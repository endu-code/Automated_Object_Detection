��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS?  �DMM�A@�  @ $��AbEREG_OFl�B�BME�HAS�C�1�A !�ARE�-   � �0�B{F S{T� �M�DTRS$ST1D6XlQCWFA� 7X �QCW�"YV�"eS/ �A~7   $�@�TINd@�0SkUL� �R_@�  $}@ S�W@�RO�RR�%	 �P�T� Ɔ@JU� �SqFS;4D6
 �2P�0�_@cFOL[d!$FIL� jjEʄP�C�S�aDI~G4RC_SCA���cINTTH�RS_BIdA�dS�MAL�bCOL��bG�`� �� ��_IVTIM��$!0B"�$S?0xCCBDSDN��-qI2wT2w�DEBUdA\!SCHN�"TOfa0�!  � Q0mr<0V� ��;!�rAUTTUuN� TRQaʤuE40N �qFS'3AXG  � 1heb}t�rI�v5�q�G_gr7 l ��!�3@WEIGYH�q�2 uS_5Q5F(�T2�WA� 	p�EsNTERVA �; - Q�� S!�t��AS0S�$J-_7STA�p JQg����1(���2��3��W���� hqx��"_COG_X�Y��Z�ҁCM�p?��p�܂RSLT �4��D��D��	"�_�p_�q7  ��~�b#0VROUN�DCMVPERIO�DA�1PUU3F2D�'TM1� �Ƒ�_D��GAMMxc1�TRXI��K�K�K��CLtbP�&O00ADJ�[GAu�UPDB
�@�:p%0 ,$�M"P30f��� d�:pG p"���HCD�GV�#G�VY��Z�JDO�5�,q��S��$R���E_8@{٣�.pAPHBC���$VF6�P��2L��蘨@IL[�����;���;�d@���R<G���NEW_���r��Q}���ڡ�5OB�OA@fY�sW2/�G�<�	����ȴ\�2�E�KP�NUCNPR�GOV����@`d_STW�c,�G�E^!�NV2#C�c0@�WT�S�TRL_SK=I2!$SJ�Q��NQpGW���s��7 �\ ;0FRf]b� � CMDC����T�b���TO�?��� �5گ���_��Ah 0 '��ALA�RM�_�*�TOT�6�FRZn l�,!Y  3��X!��mӥ�X ��@�`X �ʕ�U#��2���2
�X#Z���FIXD�8��F�"��IT��`IB�PN_d��CqH�%��_DFL �_�BF2N�ڶ�3 ����� ��3�"�怉���ʷ�� ����3���3
��X��DIAA����/#� ���%�����[1��g1 �[���Z��#��!���%���$0�@
p���7F��D�� HA¿pU�5����Q�_FwSIW6 �2P�N@�`R>!�PH;MP�`HCK%���@>0G�'*#e A����pNT��^H	��HUFRzs3��A2��UgvCa�$v0Q? ����@p�@p �  SI�0�  ��5�IRTU�_��� %SV 2���   �P6>0]@]	Q<�EF@ �o|P�  @p� � �//'/9/�K/U%@pd@p
m h K�/w/�/�/�(��$ ��/� �/�/?.8e" �/?J?\?r?8?�?|? �?�?�?�?�?�?>O4O bOO�OTO�O�OjO|O �O�O�O_�O(__\_ f_�_B_�_�_�_�_ o �_$o�_Ho>oo^b�/��o{�%�/�o�o�k�	MC: 56�78  Afs�dt1 78901234q#5w/  	q 6xzc.Ops�'���j l�o�o��� ������,�5�~DMM �)5�A ��x���𨏺�=���OR 2]	Q� ��m���_� tuB?�)DN�S�4D 
Q�!tY�d�!Ls|�q`rlƈ̀?�l�B����$ ONFIG� �(o� �� �����i!��� 2�,�
Hand g�uide��?�3����  �X���с��ь�g#?�=���A��ύ �������p�ݯ� (��L�7�p�[����m*������ʿ ܿ� ��$�6�H�Z� lɌ��ό��ϰ����Ϡ���
�C�E�I �2Q�(�0�� -�zՀ�Fտ���_`πB����d�C��  ��uq=#׽
_aNnk(��K�����̥@��=e��=D����_a�;����8I�y�_aIt$ �}$F�>���k"����Q�Fۀ3]儢ѯǯ���!�/�``+�����.������_a$�=���(4$����޷�>�E��B<�~w%�_a8E�y�5�;�jA��Ҝ{�Q�>��]�_a?��m��箑����<~u1�?�33����0�:�o����0�@����LSB�� ~uq�ӻ��m��S]���8��� ���t�	eF|���]���
�����n�O�;�.����3��'	�����B���4* 2/�V��%D�DH  *%v�+��^-���
�/��/u/~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?;)�7�?�?�o�?�8Jhq�?�?�zyjG�_FSIW Q��9��O�O �Ou�