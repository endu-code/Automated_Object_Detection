��   m�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING,��<$1_8k  �FMS*�t *v M_LIF��u,(8*x��M(DSTB0+_0>*_���*#�z&+CL_TIM>�PCCOMi��FBk M� �MAL_�EC�S��P!Q%XO �$PS� �TI����%�"r $D�TY?R. l*1E�ND14�$1�ACST1#4V22\93\9�4\95\96\6_O3VR\6� GA[7�2 h7�2u7�2�7�2�7�2ޜ8FRMZ\6DE��DX\6CURL� HSZ27Fh1DG u1DG�1DG�1DG�1DC�NA!1?( �sPL� + ���STA23TRQ_�M��/@K"�FSUX�JY�JZ�II�JuI�JI�D �$U1�SS  ����6Q�� ?P+PVE�RSI� 4W�  �5GQIRTUAL3_EQ'� 1 TX + ��(P���_��_�_�Vm���څ �!� ���~��������R?����?��J�By�4���=�t��7�Q��]�����V��u��������� ��_�Pe�ygwe�YAQ�o�^A���O ��b� I ����� �o�o�_�l/V�Set�$�w�g �B�w�un�Q�� Su���g�`� ��`���	 j�����& ~����j��b%���d�o#�5�G���=L3��R�y�?�z���@�����я���� �+�=�O�a�s���� rU������ޟ:T  2��!�3�E��W�i�{���������< ��ۯ����#�5�G��Y�k�}��������$n$ 1�\�a�Pj�J�4��J�ݖT_�b�P��N����mD�EJ���:Ha�@�J�`BB��@G(��mAɆ|1φ�|�mB�@kB�����`��C+����Pk��.dP�o�Ϙ�ϸ�+��=ϟ���M�x����2ߡ�V�A�z���s @P�� �֨�՞՞� ���{�Ђ�K�}gL��3L�X�������L�c��MZQ�MZR�<MZS�MZZU��3�8��H�L�VM]_+NN\�q�td� ���t�������6Q�Q� ������8NS_$T�i��i�����/U ��� ��� x
�� x����_����NQ��Q��sQ�WQ�BM�C��T�C���C���������E����������������Ə����%���^���p��C����C�F�C��4�C���C�������� �6g��� �7 4��7 m�t ��ZN �X� ��W �Ts ��1�5��&�N� �s�W �/4 ��4� �59�m�9������{���M��Q�� ��r�Na��,a�$a� 2���ړ����� ���vc_+�{��M��M��M��M��M�I����ѡ�š����}� t�� 0�q� 1� 1��L 1ح����u��EA����@��s���������_�������z���N����M�Ƞ�7��9��O�K��� w�3��n�	 1	 i	 � ��Ġ��1g����F Av��Wq�����#��U+��&��8��'��>�HdUc

eAPIHJ��`K���k}+����1sP�H��xtesP�EY�Q���`hsP��td��8f������� �2  ��?S	P-��sewasP!?P�O�sP������9�������}l>�����hiX�A�s�sP쩀�>����� ������{� ⩀���H楄��ssP��bsP�sP�sP�ީ�(����������sPd���ͭM��AQO���4-8���P�Ǡ_� =��WSsP��эiF.�'ce�+�/`,�/�$����??H���*���I�ڼ�D�@�^�0g��0p�D��=��.�Ħ^��맓�0��0�?������&J���L��.c��/�m�@�z�0���06�0G�0P�0Yޙ?�s��0�?��t_?�.k�����?-��?�-��?-��?�-�x?���@���?���?�)�?�~�?���?�q`!@_�?�r")@�)@����z�w9@���z�������b?��>����I.��\����v�u�l���ſ��]��2���!��{.��zۮ��z�;y@�y@�9@��@?���@���BA�=�˯@K��@5�@D��@N=%��>y��">�w�޿��@Gh�@կ@?�E�@ߍ@��@ʍ@�5Bh�b�hΪ�@��"��V��>�����,���m���;B���f���/?���?��׫�M?��:E�i�_�h�ճ�h�9�h��W�hѻ)Pm���B��B���9Q�ݫ�?��K��Jvh�J�u�MP}MP8?�����i��C�͆?+���u�9P!5P
5P�5P 5P9P�� ,�($not a program|?����_�_�_�_�_PLACE�_%o�_Io0hZERXmoTofo�o��o�o�o�o�o4dFRAM�o,7oP7I�($A�q_PO�SPIC���xA ��_q���� #�`�G���k�}������ޏ��PLCLų��� �D1�ѐ?�  ��>���?C��q�T�m�x�c��� ������������� >�P�