��   ���A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCFR_�LTST_T � l$TP�_PROG �%$DATEJ �$TIMR2SU�F_NUM  w$TlSCHm��CHSoER�Rm  $APPL_TYPR �� INI_POS�  �FRC�FIN�MAX��	�DF�FS�_��Pq V_LENORI� I  �INS'DUM_UR�GL� Q�FORCE_OK~�MOMENTe�END_AVE_�F_��OSC_�GDW�� _OFoST �  /�COM9  �$TOTAL �� 5 2  ��AL�  l ASew� ������ +=Oas���A!: ��//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?��D9 8 $~� 2 �1��@ (�A4ID�X��1�H���$$�CLASS  O���"Q��'���'PVERSIO�NX  ��53QIRTU�� _2P��@X'��� %  ����_�_�_�_��9 �S�� �_o o/oAonoeowo�o�o�o���o�o�o. @�oEW���_��_ ����_s�2�)� ;�T�_�q�����	 ����׏�.�@���E� W���������ϟ� k���!�N�E�W�p� {�����̯���� &�8���\�O���㟤� ߟ��ǿ���u��4� +�=�j�a�sόϗ��� ��������0�B߹� G�dߋ���׿�߿ߧ� ��m���#�P�G�Y� ��}��������� ��(�:���^�Q���� ���߷������w�	 6-?lcu�� ����� 2� Iz������� ���oe/%/R/I/ [/�//�/�/�/�/ ?�/*?<?�/`?S?� �?��?�?�?�g?�? OO/OAOnOeOwO�O �O�O?�O�O�O"_4_ �OD_K_|_�?�_�?�_ �_�_�?q_oo'o9o Ko]o�o�o�o�o�o_ �o�o�o,>�obU �_��_����_i ���8�C�U�g�y� ����ʏ� �ߏ$� 6���Z�M�~����� ��ş��s��2�)� ;�T�_�q�����¯	� ����ׯ�.�@���E��W����$CCFR�_D ������'� ����ܟο�� ��r� �M�D�V�h�z� �Ϟϰ��������� �I�[����r߈��� �������φ�3�*� <�i�`�r������ ��.�����A�S��� w�j����߿������� ��"OFX� |����&�� �9K]�bt�� �������5/ ,/>/k/b/t/�/�/�/ �/�/0??�/C?U? �/y?l?� /�?��? �?	O/�?$OQOHOZO �O~O�O�O�O�O(?_ _�O;_M___�Od_�_ �?�_�?�_�_oO�_ 7o.o@omodovo�o�o �o�o�o2_! E W�o{n�_��_� ��oo�&�S�J� \������������* ����=�O�Ə8�f� ������̟ޟ�� ����0�B�o�f�x��� ����ۯ�4��#�� G�Y�Я}�p������ �ֿ����1�(�:� L�^ϋςϔ��ϸ��� ,�	����?�Q���u� hߙ߬���������� ώ� �M�D�V�h�z� ��������6���� �I�[����r��ߵ� ����������3* <i`r���� �.��AS� wj��������� /�"/O/F/X/�/ |/�/�/�/�/&�/? �/9?K?]?�/b?t?� �?��?�?�?/�?5O ,O>OkObOtO�O�O�O �O�O0?__�OC_U_ �Oy_l_�? O�_�?�_ �_	oO�_$oQoHoZo �o~o�o�o�o�o(_ �o;M_�od� �_��_���o� 7�.�@�m�d�v����� ��ُ�2�!� �E� W�Ώ{�n������� ԟ�����&�S�J� \������������*� ����=�O�Ư8�f� ��������̿޿�� ����0�B�o�f�xϥ� �Ϯ�����4��#�� G�Y���}�pߢ���� �����τ�1�(�:� L�^��������� ,�	����?�Q���u� h����߽������� �� MDVhz �����6�� I[�r��� ������3/*/ </i/`/r/�/�/�/�/ �/.??�/A?S?�/w?j?�?(��?� �?�?	O/�?$OQOHO ZOlO~O�O�O�O�O�O 6?_�O_M___�O�_ v_��_�?�_�_�_O �_7o.o@omodovo�o �o�o�o�o2_!  EW�o{n�_o� �_���o�&�S� J�\������������ *܏���=�O�a�؏ f�x�����̟ޟ�� ���9�0�B�o�f�x� ���������4��#� �G�Y�Я}�p���� ſ �ֿ�� ���(� U�L�^ϋςϔ��ϸ� ��,�	����?�Q�c� ��hߙ߬��������� �ώ�;�2�D�q�h� z��������6�� %��I�[����r��� ���߲������"�� *WN`���� ��.��AS �<j������� �/��4/F/s/ j/|/�/�/�/�/�/8 ?'??K?]?�/�?t? ��?���?�?/�? 5O,O>OPObO�O�O�O �O�O�O0?__�OC_ U_�Oy_l_�_�?�_�? �_�_	oO�_$oQoHo Zolo~o�o�o�o�o�o :_�oM_�o� v�_��_���o �7�.�@�m�d�v��� ��Ǐ���2�!� � E�W�Ώ{�n���ß �ԟ�����&�S� J�\������������ *�ܯ���=�O�a�د f�x�������̿޿�� ���9�0�B�o�f�x� �ϜϮ�����4��#� �G�Y���}�pߢ�� �� ������ ϖ�(� U�L�^������� ��,�	����?�Q�c� ��h����߽������� ��;2Dqh z�����6� %I[�r�� ������"� */W/N/`/�/�/�/�/ �/�/.??�/A?S? �/<?j?�?��?��? �?O/�?�?4OFOsO jO|O�O�O�O�O�O8? _'__K_]_�O�_t_ �?�_�?�?�_�_O�_ 5o,o>oPobo�o�o�o �o�o�o0_�oC U�oyl��_��_ ��	�o�$�Q�H� Z�l�~��������� :����M�_�֏�� v�����ʟܟ�� ��7�.�@�m�d�v��� ��ǯ���2��!� � E�W�ί{�n����ÿ ��Կ�����&�S� J�\ωπϒϤ϶��� *������=�O�a��� f�xߪ��������ߴ� ό�9�0�B�o�f�x� ��������4��#� �G�Y���}�p���� �� ����� ��( UL^����� �,�	�?Qc �h�������� /�;/2/D/q/h/ z/�/�/�/�/�/6? %??I?[?�/?r?� �?��?�?�?/"/�? *OWONO`O�O�O�O�O �O�O.?__�OA_S_ �O<_j_�_�?�_�?�_ �_oO�_�_4oFoso jo|o�o�o�o�o�o8_ 'K]�o�t �_��_�_��o� 5�,�>�P�b������� ŏ���0����C� U�̏y�l������� ҟ�	����$�Q�H� Z�l�~��������� :�����M�_�֯�� v�������ʿܿ�� ��7�.�@�m�d�vψ� ���Ͼ���2��!� � E�W���{�nߠ���� �������ϔ�&�S� J�\�������� *������=�O�a��� f�x��߻��������� ��90Bofx �����4�# GY�}p�� � ��/ �(/ U/L/^/�/�/�/�/�/ �/,	??�/??Q?c? �/h?�?��?��?�? O/�?;O2ODOqOhO zO�O�O�O�O�O6?_ %__I_[_�O_r_�? �_�?�_�_�_O"O�_ *oWoNo`o�o�o�o�o �o�o._�oAS �o<j��_��_� ��o��4�F�s� j�|�������ߏ�8 �'��K�]�ԏ��t� �����ڟ���� 5�,�>�P�b������� ů���0�����C� U�̯y�l��������� ҿ�	����$�Q�H� Z�l�~ϫϢϴ����� :�����M�_��σ� vߨ������������ ��7�.�@�m�d�v�� �������2��!� � E�W���{�n������ ��������&S J\������ *���=Oa� fx�������� �9/0/B/o/f/x/ �/�/�/�/�/4?#? ?G?Y?�/}?p?�?�2