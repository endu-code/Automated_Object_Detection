��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV����RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DIS�� S�MB�	"�BC�J@"CI2AI<P6EXPS�!�gPARQ$�RCL�/
 <(C�0��SPTM�E� PWaR��X�V�SMo l5��!�"Y%�7�ICC�%� �kfR�0leP� _'DLV��YNoE3 <oNbX_�P~~#Z_INDE
C��`OFF� ~UR��iD��c�  � t �!�`M�ON�%sD�&rHOU�#EWA,vSq;v<SqJvLOCA� Y�$N�0H_HE����@I"/ >3 $ARPz&�1F�W_\ �I!F�`;FA�Dk01#�HO_� INF�O�sEL	% P� K  !k0WO�` $ACC�E� LVZk�2�H#ICE�L� � �$�s# ��)�k���
��
`�K`�SQi��Pk�5|�I�0ALh��z�'0 ��
���F�����P�܅�]$� 2ċT" �w������� č���!r�Z���4����Ċ!147.�87.224.2i0h�S���96��P��܁܁3�_{p_�  ċ� bfh.ch̟�1� C�U�g�y����������ӯ^�� _FLTRs  ��π ��������n�nx�č2n��rSH�PD� 1ĉ  �P!
robst�ation֯՚!k�.�Q�ſ�� ������޿?��c� &χ�JϫϽπ��Ϥ� ���)���M��"߃� Fߧ�j��ߎ��߲��� %���I��m�0��T� ��x��������3� ��W��{���P���t� ������������S w:�^��� ���= a$�Zׯ$ _L�A1}��x!1.��ğP�1�Q2�55.%�S���2��E �//*/<&3F/�� l/~/�/�/<&4�/�50 �/�/??<&56?�@�0\?n?�?�?<&6�? �%@�?�?�?
O1�?P���MY� M?Y��c��� Q� �VN<�O�O_�O+_=_ O_"_s_�_NPd_�_ �_�_�_�_o!o3o�_Woio{oVNLoM� �o�l�oAo
.@�U}iRCon�nect: ir�c\t//alertsE����Pu ����1�C�U�уP_R8�d�� H�~�������Ə؏ꏀ��� �2�D�V�S$���8�(p����o͟�ߟ��QA8��d�A�B4��j�h9�rQ+��@DM_�A�+��SMB 	X�8%ğVO��߯����_CLNT �2
X� 4C� ɯ0��l�c�B�T��� x���Ͽ������)π;��_�q�Pϕ��M�TP_CTRL ��%���ϙdc� ��ߋ��?�*�c߳l2��N���@{�V����Ƥ��������ѓC��USTOM' {���}�@� }�DTCPIPu�{��h�E��TEL�{��A���H!Ta�t�ç�roblol�r�  ���!KCL���F��!CRT���������!CON�S&����n+���