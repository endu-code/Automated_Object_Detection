��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER�mq�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS9?  �DMM�A@�  @ $��AbEREG_OFl�B�BME�HAS�C�1�A �DRE�-   � �0�B{F S{T� �M�DTRS$ST1D6XlQCWFA� 7X �QCW�"YV�"eS/ �A~7   $�@�TINd@�0SkUL� �R_@�  $}@ S�W@�RO�RR�%	 �P�T� Ɔ@JU� �SqFS;4D6
 �2P�0�_@cFOL[d!$FIL� jjEʄP�C�S�aDI~G4RC_SCA���cINTTH�RS_BIdA�dS�MAL�bCOL��bG�`� �� ��_IVTIM��$!0B"�$S?0xCCBDSDN��-qI2wT2w�DEBUdA\!SCHN�"TOfa0�!  � Q0mr<0V� ��;!�rAUTTUuN� TRQaʤuE40N �qFS'3AXG  � 1�eb}t�rI�v#G_|gr7 l �!|�3@WEIGH�qV�2 uS_5QF(�MT2�WA� 	pEs?NTERVA�; @- Q�� S!�t�AS0�S�$J-_ST�A�p JQg���1�(���2��3��W����� hqx��"COWG_X�Y�Z�6ҁCM�p?�p<�܂RSLT�4� �D��D���@�!�@�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDB Q:p%_0 ,$M"P380f��� d�:ppG p"��HCD��GV�#GVY��Z��JDO5�,q��Sn��$R��E_8@�{٣�pAPH�BC��$VF�6�P��2L��蘨@IL[����;���;��d@���RG���NE#W_���r�Q}����ڡ�5OBOA@fY(�sW2/�G<�	����ȴ\�2�E�KP�NUCNPRGOV��8��@`d_TW�c,�5G�E^!NV2#C��c0@�WTS�TR�L_SKI2!$�SJ�Q��NQpGW�P���7 \ m;0FR]b� � CMDC���T�b���TO?��� �5گ���_�Ah 0 '�>�ALARM�_��*�TOT6�FRZn l�,!Y 3��X!�� mӥ�X �Œ`X �ʕ�U#��2��2
�X#Z�N��FIX�8��F�"d��IT�`IB�PN_d��CH�%���_DFL _�BF2N�ڶ�3����� ��3�"�����ʷ�(� ����3��3
��X��DIA����/#� ���%��� ��[1��g1�[���Z���#��!���%����$0�@
p��7F��D,�� HA�pU�5����v�FSIW6K �2PN@�`R>!��PHMP�`HCK%���>0G�'*#eb A����pNT��p^H	��HUFRzs�3��A��UgvCa��$v0Q ��i��@p@p � � SI0��  �5�I�RTU_��� %S�V 2���  A  P4>0]@]�	Q�EF@ �oP�  	@p� � �//�'/9/K/U%@pd@p
m hK�/w/�/�/�( ��$��/� �/�/? .8e"�/?J?\?r?8? �?|?�?�?�?�?�?�? >O4ObOO�OTO�O�O jO|O�O�O�O_�O(_ _\_f_�_B_�_�_�_ �_ o�_$o�_Ho>oo ^b�/�ot��%�/�o�o��k	MC: �5678  A�fsdt1 78?901234q$#5w ��	q 6xzc.Ops�'���j l�o�o��� ������,�5�~DMM �)5�A ��x���𨏺�=���OR 2]	Q� ��m���_� tuB?�)DN�S�4D 
Q�!tY�d�!Ls|�q`rlƈ̀?�l�B����$ ONFIG� �(o� �� �����i!��� 2�,�
Hand g�uide��?�3����  �X���с��ь�g#?�=���A��ύ �������p�ݯ� (��L�7�p�[����m*������ʿ ܿ� ��$�6�H�Z� lɌ��ό��ϰ����Ϡ���
�C�E�I �2Q�(�0�� -�zՀ�Fտ���_`πB����d�C��  ��uq=#׽
_aNnk(��K�����̥@��=e��=D����_a�;����8I�y�_aIt$ �}$F�>���k"����Q�Fۀ3]儢ѯǯ���!�/�``+�����.������_a$�=���(4$����޷�>�E��B<�~w%�_a8E�y�5�;�jA��Ҝ{�Q�>��]�_a?��m��箑����<~u1�?�33����0�:�o����0�@����LSB�� ~uq�ӻ��m��S]���8��� ���t�	eF|���]���
�����n�O�;�.����3��'	�����B���4* 2/�V��%D�DH  *%v�+��^-���
�/��/u/~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?;)�7�?�?�o�?�8Jhq�?�?�zyjG�_FSIW Q��9��O�O �Ou�