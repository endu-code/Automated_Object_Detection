��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SF�TVER����_�GRP6� �2$FS_FOR�C� ��P�S_GMEA2'%� 1G�F#2G0 �GTS_K_CHKY%O �RIc"]!APP��$PS_AA�ML��$�"�	]$/!_MI2�$AS�!!�#'#�#�!��3  2 RO�M_RU2$Jn� EST2!$� ��N_NU�$�u �  
$SBn*BSCNCTO�INS29FS� _�NG$GAG�Ex� � CUToFREQY#LR*�REAL%� �2M�OMEN�T�V�C�F�C��2N�C�K1DT��1D�EVIDS�7 {	�3PATH�0]A�3FNA� 6!�	AEX� �5O �8BUF�7TDP�Y�FLGEJ5�� � � N IU�
@!(UF*����4OSs� ��DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� !�ARE-  ? � �0�BB{F S{T� M�D|TRS$STD6XlQCWFA� 7X�QCW��"YV�"eS/ �A7 �  $�@TI�Nd@�0SULگ �R_@ g $}@ SW�@�RO�RR%	� �P�T� �@J�U� �SqFS4DN6
 �2P�0_@�cFOL[d!$�FIL� jjE�P��C�S�aDIG4R_C_SCA��c�INTTHRS�_BIdA�dSMA9L�bCOL�b9G�`� �� ��_IVTIM��$!0B"$S�?0xCCBDDN���-qI2wT2wDE�BUdA\!SCHN�"TOfa0�! �  Q0mr<0V� �;!�r~AUTTUN�� TRQa�uE�40N �qFS3A	XG  � 1eb}tj�rI�v	"G_gr>7 l �!�3>@WEIGH�q�2� uS_5QF(�T�2�WA� 	pEsNTERVA�; -  Q�� S!�t�AS0S��$J-_STAF�p JQg���1(�U��2��3��W����� hqx��"COG+_X�Y�Z�ҁCM�p?�p�܂RSLT�4��D��D��	"_�p_�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDB#	"I%�0 ,$M"Pp30f��� d��:pG p"��HCDv�GV�#GVY��Z�JDO5�,q���S��$R��E_�8@{٣�pAP�HBC��$VF6�P��2L��蘨@IL[����;����;�d@���RG���NGEW_���r�Q}�8��ڡ�5OBOA@fQY�sW2/�G<�	����ȴ\�2�E�KP��NUCNPRGOVp����@`d_TW�cj,�G�E^!NV2#�C�c0@�WTS�T�RL_SKI2!�$SJ�Q��NQpG�W���	"��7 �\ ;0FR]b� � CMDC���T0�b���TO?�� � �5گ���_�Ah �0 '��ALARM��_�*�TOT6�F#RZn l�,!Y 3�� X!��mӥ�X �Œ`X P�ʕ�U#��2��2
�8X#Z���FIX�8�ґF�"��IT�`IeB�PN_d��CH��%��_DFL _�B#F2N�ڶ�3����� ��3�"�����ʷ�� ����3��3p
��X��DIA����/#� ���%�����[1��g1�[� ��Z��#��!���%���$0�@
p��7F���D�� HA�pU��5����v�FSIW.6 �2PN@�`uR>!�PHMP�`HCK%���>0G�'�*#e A����pN�T��^H	��HUFARzs3��A��Ugv�Ca�$v0Q �����@p@p ��  SI0��  �5�IRTU_��� �%SV 2���   �6>0�]@]	Q�EF�@ �oP�O  @p� �  �//'/9/K/U%@pd@p
m hK�/w/ �/�/�(��$��/�  �/�/?.8e"�/?J? \?r?8?�?|?�?�?�? �?�?�?>O4ObOO�O TO�O�OjO|O�O�O�O _�O(__\_f_�_B_ �_�_�_�_ o�_$o�_ Ho>oo^b�/�ot��%�/�o�o�k	M�C: 5678 � Afsdt1� 7890123�4q#5w  e	q 6xz.Op�s�'��j l�o�o����������,�5�DM�M �)5�A ��x�������=����OR 2	Q�� ��m��_�� tuB?�)DN�S4D 
Q�!tY�d��!Ls|�q`rƈ̀?-�l�B𴐠�$ �ONFIG ��(m� � ������i!�� �2�,
H�and guid�e��?�3���  �X��с���ь�g#�=���A��ύ����� ��p�ݯ�(��L��7�p�[����m*������ʿܿ� � �$�6�H�Z�lɌ��� ���ϰ��������
�tC�E�I 2Q�5(�0� -�z�4��Fտ��_`π�B����d�C�  ���uq=#�
_aN�nk(��K�����̥@��e��=�D����_a;��=��8I��_a�It$ �$F��>���k"��=�Q�Fۀ3]儢�ѯǯ���!�/�``+������.������_a$敕��(�4$�����>�{E��B<~w%��_a8E�y5�;�sjA��Ҝ�Q�O>��]�_a?���m��箑����~u1�?��33����0�:�o����0�����LSB��~uq�Ӡ���m�S]����8��� ����t�	eF|�@��]��߯�����n��;��.����3�'	������B��� 4* 2/V��%D�DH  *%v�+���^-��
�/��/u/~u�J/l/�)�AI��/�/�?/ #A��n5��p��4 vO?;)�7�?�?�o�?�8Jhq�?�?zyjG��_FSIW  Q��9��O�O�Ou�