��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SF�TVER����_�GRP6� �2$FS_FOR�C� ��P�S_GMEA2'%� 1G�F#2G0 �GTS_K_CHKY%O �RIc"]!APP��$PS_AA�ML��$�"�	]$/!_MI2�$AS�!!�#'#�#�!��3  2 RO�M_RU2$Jn� EST2!$� ��N_NU�$�u �  
$SBn*BSCNCTO�INS29FS� _�NG$GAG�Ex� � CUToFREQY#LR*�REAL%� �2M�OMEN�T�V�C�F�C��2N�C�K1DT��1D�EVIDS�7 {	�3PATH�0]A�3FNA� 6!�	AEX� �5O �8BUF�7TDP�Y�FLGEJ5�� � � N IU�
@!(UF*����4OS	 D�MM�A@  �@ $�AbERE�G_OF�B�BME��HAS�C1�A �!�ARE-  � � �0�B{F S{T� M�DTRS$STD6XlQCWFA� 7X�QCW�"YV�"eS/ �A7  w $�@TINd@��0SUL� ��R_@  $}@ SW@�R�O�RR%	 h�P�T� �@JU� ��SqFS4D6
� �2P�0_@cF�OL[d!$FI�L� jjE�P�C��S�aDIG4RC_�SCA��cIN�TTHRS_ByIdA�dSMALN�bCOL�bG�`α �� ��_InVTIM�$!:0B"$S?0x?CCBDDN��-q�I2wT2wDEBU�dA\!SCHN�"TOfa0�! � Q0mr�<0V� �;!�rA_UTTUN� �TRQa�uE40N| �qFS3AXG � � 1eb}t�rI��v	"G_gr7 �l �!�3@W�EIGH�q�2 �uS_5QF(�T2�W�A� 	pEsNTERVA�; - Q�� �S!�t�AS0S�$�J-_STA�p QJQg���1(���2��3��W���� �hqx��"COG_X��Y�Z�ҁCM��p?�p�܂RSLT�4��D��(D��	"_�p_�q7 � �~�b#0VR�OUNDCMVPE�RIODA�1PUnU3F2D�'TM1�� �Ƒ_D��G�AMMc1�TR�XI�K�K�K���CLbP�&O00A�DJ�GAu�UP�DB	"I%0/ ,$M"P30f��� d�:pG �p"��HCD�G]V�#GVY��Z�GJDO5�,q��S��7$R��E_8@{t٣�pAPHBCy��$VF6��P��2L��蘨@IL [����;���;�d@���RG���NEW_���r�Q}���ڡN�5OBOA@fY�sW2/�G<�	����ȴ�\�2�E�KP�NUC?NPRGOV��Ŝ�@`d_TW�c,�G�E^!NV2#C�c0�@�WTS�TRL�_SKI2!$SiJ�Q��NQpGW���	"��7 \ m;0FR]b� � CMDC���T�b���TO?��� �5گ���_�Ah 0 '�>�ALARM�_��*�TOT6�FRZn l�,!Y 3��X!�� mӥ�X �Œ`X �ʕ�U#��2��2
�X#Z�N��FIX�8��F�"d��IT�`IB�PN_d��CH�%���_DFL _�BF2N�ڶ�3����� ��3�"�����ʷ�(� ����3��3
��X��DIA����/#� ���%��� ��[1��g1�[���Z���#��!���%����$0�@
p��7F��D,�� HA�pU�5����v�FSIW6K �2PN@�`R>!��PHMP�`HCK%���>0G�'*#eb A����pNT��p^H	��HUFRzs�3��A��UgvCa��$v0Q ��i��@p@p � � SI0��  �5�I�RTU_��� %S�V 2���  A �@4>0]@]�	Q�EF@ �oP�  	@p� � �//�'/9/K/U%@pd@p
m hK�/w/�/�/�( ��$��/� �/�/? .8e"�/?J?\?r?8? �?|?�?�?�?�?�?�? >O4ObOO�OTO�O�O jO|O�O�O�O_�O(_ _\_f_�_B_�_�_�_ �_ o�_$o�_Ho>oo ^b�/�ot��%�/�o�o��k	MC: �5678  A�fsdt1 78?901234q�#5w  	q �6xz.Ops�'��j l�o�o����������,�5�DMM 1�)5�A ���x�������=���ORw 2	Q� ���m��_� tu�B?)DN~�S4D 
Q�#!tY�d�!Ls|��q`rƈ̀?�l�B�𴐠�$ ONF�IG ��(� -� �����i!s�� 2��,
Hand� guide��?��3���  ��X��с��ь��g#�=���A ��ύ�������p� ݯ�(��L�7�p�[�<���m*���� ��ʿܿ� ��$�6� H�Z�lɌ��ό��ϰπ�������
�C�E�I� 2Q�(�0�� -�zՀ�Fտ&��_`πB���Ԟd�C�  ��uq=�#�
_aNnk(���K����̥@���e��=D�����_a;����8�I��_aIt$� �$F�>����k"���Q�Fۀ3]儢ѯǯ�����!�/�``+��̞��.�����_a$�敕��(4$�x����>�E���B<~w%�_a8E{�y5�;�jA���Ҝ�Q�>�	�]�_a?��m��箑�����~u1�?�33x����0�:�o�� ��0�����LSB��~uq�ӻ��m��S]���8��� ���t�	eF|���(]��߯����<n��;�.����=3�'	�����B���4* �2/V��%D�DH#  *%v�+��^-��
�/��/u/~u#�J/l/�)AI��/p�/�?/ A��n5��p��4vO?;)@�7�?�?�o�?�8Jhq�?�?zyjG�_FSIW Q��9�� O�O�Ou�