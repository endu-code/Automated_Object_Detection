��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1d�DDd!OE4LA!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTc@�D5�F6�F7�F8�F9�G0�G�GJA��E�GbA�E�G1�G1��G �F�G2�B!S�BN_CF>"
 }8F CNV_J� �; �"�!_CMNT��$FLAGS<]�CHEC�8 �� ELLSETU�P � $H�O30IO�0� %��SMACRO�RR'EPR�X� D+�0��R{�T UTO�BACKU��0 �)DEV�IC�CTI*0��� �0�#�`B�S$�INTERVAL�O#ISP_UNI�O`_DO>f7ui�FR_F�0AIN��1���1c�C_�WAkda�jOFFu_O0N�DEL�h�L� ?aA�a1b?19a�`C?��P�1bE��#sATB�d���MO� �cE D [M�c���^qREV�BIL�rw!XI� QrR o � OD�P~�q$NO^PAM�Wp�t�r/"��w� �u�q�r�0D~`S p E �RD_E�pCq$�FSSBn&$CH�KBD_SE^eA�G G�"$SL�OT_��2=�� V��d�%��3 a_�EDIm   �� �"��PS<�`(4%$EP�1�1O$OP�0�2�an�p_OK�UST1P_C� ��d��U ^�PLACI4!�Q��4�( raCOMM� ,0$D����0��`��EOWBn�IGA�LLOW� (�K�"(2�0VAR�a��@�2ao�L�0OUy� ,Kvay�r�PS�`�0M_O]�����CCFS'_UT~p0 "�1 �3�#�ؗ`X"�}R�0  4F IMC	M�`O#S�`��up�i �_�p�BA�!���M/ h��pIMPEE_F �N��N���@O��Fr�D_�~�n�Dy�9F� dCC_�r0  T� '��'��DI�n0"��p:�P�$I��t����F�t X� �GRP0��M=qN�FLI�7��0UI�RE��$g"� SW�ITCH5�AX_�N�PSs"CF_L�IM� � �0EED��!��PqP�t�`PJ_dVЦMODEh�.Z`�P|Ӻ�ELBOF�  ������p� ���3���� FB/��0t�>�G� �� �WARNM�`/�p�qP��n�NST� �COR-0bFL{TRh�TRAT�P�T1�� $ACC�1a��N ��r$OcRI�o"V�RT�Ps_S� CHG�0I��rT2��1�I��T�I1��� x i#�Q�.�HDRBJ; C�Q�2L�3L�4L�5�L�6L�7L� N�9�{5CO`S <�F +�=�O��#92��L�LECy�"MULTI�b�"N��1�!t���0T�� �STY�"�R`�=l��)2`����*�`T  |� �&$��۱m�a�P�̱�UTO��:�E��EXT����pÁB���"2� (䈴![0������p<�b+�� "D" ���ŽQ��<煰kc��*�9�#���1��ÂqM�ԽP��" '��3�$ L� E���P<��`A�$JO�Bn�T���l�TRIG3�% dK����� ��<���\��+�Y�p��_M��& tf�pFLܐBNG AgTBA� ���M� �
�!��p� �q��0��P[`��O�'[���0tna*���"MJ��_R���CDQJ��IdJk�D�%�C�`�Z���0��Pq_�P��@ ( @F �RO.��&�t�IT�c�NOM�
�����S6�CP`T)"w@���Z�P�d���RA�0��2b"�����
$T����MD%3�T��`U31��ʩp(5!HGb�T1�*E�7�c�KAb�pWAb�cA4#YNT��>�PDBGD�� *(��PUt@X���W���AX��a��ewTAI^cBUF���0!+ � l7n�PIW�*5 P�7M�8M�9
0�6}F�7SIMQS@�>KEE�3PAT�n�^�a" 2`#�"�L�64FIX!, !���!d��D�2Bus�=CCI�:FPCH�P:BAD�aHCEhAOGhA]HW�_�0>�0_h@�f�Ak���F�q@\'M`#�"�DE3�- l�p3G��@FSOES]FgHBSU�I�BS9WC��. ` =��MARG쀳β�FACLp�SLEWxQe�ӿ�6�MC�/�\pSM_JBM����Q�YC	g�e��w0 ā�CHN-�;MP�$G� Jg��_� #��1_FP$�!TCuf!õ#@�����d�#a��V&�0�r�a;�fJR���r�SEGFR�PIO�� STRT��N��cPV5���!41�r��
r>İ�b�B��O�2` + �[���,qE`&�,q`�y�Ԣ}t��yaSI!Z%���t�vT�s� ��z�y,qRSINF }Oбc���k��`���`�`L�ĸ T`7�C3RCf�ԣCC/�9���`a�uah�ub'�MI�N��uaDs�#�G�D
�YC��C�����e�0q0��� �EV�q�UF�_�eF��N3��s�ah��Xa+p,�5!�#1�!VSCIA?� A��s1�"!3 ��`F/k��_ �U��g��]��C�� a��s��R�4� �����N����5a�R��HANC��$L�G��P�f1$+@NYDP�t�AR5@N^�`�a�q���c��ME�108���}0��RAө�CAZ 𨵰�%O��FCTK��s`"��S�PFADIJ�O J�ʠ�ʠ���<����Ր��GI�p�B�MP�d�p�Dba��AcES�@	�K�W_���BAS�� �G�5 � M�I�T�C�SX[@@�!62�	-$X���T9�{s�C��N�`�a~P_H�EIGHs1;�WI�D�0�aVT ACϰ�1A�Pl�<����EXPg���|��C}U�0MMENU���7�TIT,AE�%)�a2��a��g8 P� a�ED�E� ��PDT��R�EM.��AUTH?_KEY  ������ �b�O	�!}1�ERRLH� �9 1\� �q-�OR�DB��_ID�@l �PUN�_O��Y�$SY�S0��4g�-�I��E�EV�#��(�PX�WO�� �: $�SK7!f2�DBT�d�TRL��; ��'AC�`��ĠINMD9DJ.D��_��bf1��f���PL�A��RWAj���SD��A��!+r|��U�MMY9d�F�10�d�&���J�<��}1P�R� 
3�PO9S��J�= ��$V$�q�PLB~�>���SܠK�?�����CJ�@����EN5E�@T��A���S�_�RECOR��B�H 5 O�@7=$LA�>$~�r2��R��`�q�b`�_DLu��0RO�@�aT[� Q��b������! }О��PAUS���dE�TURN��MR�U�  CRp�E�WM�b�AGNAL:s2$LA�!�?$PX�@$P�y A �Ax�1C0 #ܠDO�`X��k�W�v�q�GO_A7WAY��MO�ae����]�CSS_C�CSCB C �8'N��CERI����J`u�QA0�}���@�GAG� R �0�`��{`��{`OF�q�5��#kMA��X��&���LL�D� �$���sU�D)E%!�`���OVR10�W�,�OR|�'�$�ESC_$`�eDSGBIOQ��l �\�B�VIB&� �c�,�����f�=pSS�W���f!VL��P�L���ARMLO�
��`����d7%SC �bALspH�MPCh �Ch �#h �#h 5�UU���C �'�C�'�#�$'�d�#AC\4�$�pH��Ou�0�!Y��!�SB�� �`k$4�C�P3Wұ~46$VOLT37#$$`�*�^1�0�$`O1*�$o��0�RQY��2b4�0DH_THE����0xSЯ4�7ALPH�4�`���7�@ �0�qb7�rR�5�88� �×���"��Fn�MӁVHBPFUBAFLQ"D�s�`�THR��i2dB�����G(��PVP�����(������1�J2�B�E�C�E�CPSu�Y@� �Fb3���H�(V�H:U �G�
X0��FkQw�[��Na�'B���C IN{HBcFILT�� �$��W�2�T1�[� ��$���H Y6АAF�sDO��Y �Rp� fg�Q�+�c�5h�Q�iSh�QPL��Wqi�QTMOU �#c�i�Q\��X�gmb���vi�h�bAi�fI��aHIG��ca	xO���ܰ��W�"vAN�-u!��	#AV�H!Pa8$P�ד#p��R_:�A�a��B��N0�X�MCN`���f1[1�qVE�p��Z2;&f�I�QO�uh�rx�wGldDN{G|d��aF>!�9�r�aM:�U�FWA�:�Ml���X�Lu��$ !����!l�ZO�����0%O�lF�s�13�D	I�W�@��Q����_��!CURV�A԰0rCR41ͰZ �C<�r�H�v���<�`0��<�(�f�CH�QR 3�S���t���Xp�VCS_�`�ד�F���ژ���?N�STCY_ E L����1�t�1�T�U��24�2B�NI �O7������DEV�I|� F��$�5�RBTxSPI2B�P���BYX�����T��HNDG>��G H tn���L��Q�C���t5��Lo0 H���閻�FBP�{tF�E{�5�t��T��I��DO���uPMC�S�v>�f>�t�"HOTSW�`s�%҈wELE��J T��@�e�2��25�� O� ��HA7�E��344�0q?��A�K �� �MDL� 2J~PE��	A��s��t��È�s�JÆG!��r�D"�ó�����\�TO���W�	��/��SL{AV�L  \0INPڐ���`%ن�_CFd�M� $��ENU��O�G��b�ϑ]զP�0�`ҕ�]�IDMA0�Sa��\�WR�#���"]�VE�$a�SK�I�STs��sk$��2u���J�������	��Q���_SVh�E�XCLUMqJ2M!ONL��D�Y��|�P�E ղI_V�A�PPLYZP��HI�D-@Y�r�_M�2��VRFY�0��r�<1�cIOC_f��"� 1������O��u��LS���R$DU/MMY3�!���S=� L_TP/Bv��"���AӞ�ّ Ns ���RT_uN�� P@�G&r�[�O D��P_B�A�`�3x�!IF ��_5���H������� �� P� $�KwARGI���� q�2O[�_wSGNZ�Q �~P/�/PIGNs�l��$�^ sQANNUN�@�T<�U/�ߴ�LAzp]	Zh�d~,�EFwP}I�@ R @��F?IT�	$TOTA%��d���j�!�M�NIY�CS+���E�A[��
DAYS\�AD�x�@��	� �E�FF_AXI?�T�I��0zCOJA ��ADJ_RTRQ��Up��<P�1D �r5̀Ll��T�p? ]P�"p��M��Atpd��V 0@w�G���������SK�SU� ��C�TRL_CA�� �W�TRANS��6PIDLE_PAW���!��A�V���V_�l�V ��DIAGS���X� /$2�_SE�#TAC���t!�!00z*@��RR��vP�A���p ; SW��!�!�  ��ol�U���oOH��PP̱ ��IR�r��BR1K'#��"A_Ak��� x 2x�9ϐZs2���%l�W�pt*�x%R7QDW�%MSx�t5�AX�'�"��LIF�ECAL���10��N�1{"�5Z�3{"�dp5�ZU`}�MOT�N°Y$@FLA��cZOVC@p�5H�E	��SUPPOQ�ݑAq� Lj (C��1_X6�IEYRJZRJWRJ�0TH�!UC��>6�XZ_AR�p�Y2�HCOQ��S�f6AN��w$
�U C�TE�Y `��CACHE�C9��M�PLAN��UFFIQ@�Ф0<Ѩ1	��6
���M�SW�EZ 8�K�EYIM�p��TM~�SwQq�wQ#���>��OCVIE� �w[ A�BGL��/�}�?��@�?��D�\p�ذST��!�R� �T� �T� �T<	��PEMAIf�ҁ���_FAUL��]�Rц�1�U��� �TRE�?^< $Rc�u�S�% IT��BU!FW}�W��N_� 'SUB~d��C|��8Sb�q�bSAV�e�b�u �B��� �gX�^P �d�u+p�$�_~`�e�p%yOTT����s�P��M��OtT�LwAX � ��X~`9#�c�_G�3
�YN_1�_�D��1 �U2M���T��F��H@ g�`� 0p��Gb-s7C_R�AIK���r�t�RoQ�u7h�q'DSPq��rP��A�IM�c6�\����s2��U�@�A�sM*`I�P���s�!DҐ6�T!H�@n�)�OT�!6��HSDI3�ABSC���@ Vy���� �_D�CONVI�G���@3�~`	F�!�pd��psq�SCZ"���sMER�k��qFB��k��pEiT���aeRFU:@�DUr`����x�CAD,���@p;cHR�	A!��bp�ՔՔV+PSԕC���	C��p�ғSp�_cH *�LX� :cd�Rqa�| ����W� �U��U��U�	�U�TOQU�7R�8R�9R���0T�^�1k�1x�1���1��1��1��1*��1ƪ2Ԫ2^�k�U2x�2��2��2��U2��2��2ƪ3Ԫ%3^�3k�x�3���To���3��3��3ƪ54Ԣ&%�XTk!0�d <� 7h�p�6�p�O��p����NaFDR^Z$eT^`V��Gr����䂴2REMr� Fj��BOVM�z�A�TROVٳDT�`-�MX<�I�N��0,�W!IND�KЗ
w�׀�p$DG~q36��P�5�!9D�6�RIV���2��BGEAR�IO�%K�¾DN�p��J��82�PB@�CZ_MCCM�@�1��@U���1�f ,②a?� ���PI�!?I�E��Q�$��a�m���g� _0Pfq�g RI9ej�k!UP?2_ h � �cTD�p���! a�纱���BAC�riC T�P�b�`�) OG��%���p��IFI�!�pm�>���	�PT�"i�MR2>��j ��Ɛ +"����\��������P$�B`x%��_ԡ��"�_���� M���߾��DGCLF�%D7GDY%LDa��A5�6�ߺ4@��UkM`��� T�FS#p�Tl P���e�|qP�p$EX_����1M2��2� 3��5��G ���m� ��Ѝ�SW�eO>e6DEBUG����%GR���pU�#B�KU_�O1'� �@PO�I5�l5MS��OOfswSM��E�b�Q�0��0_E n ��0 Ɛ�TERM�o��UPORI�+�p�P�SM�_���b�q�!� �TA�r�2�O �UP�Rs� -�1�2n$|�' o$SEG,*�> ELTO��$wUSE�pNFIA�U"4�e1���#$p$UFR���0ؐO!��0����OT�'�TqAƀU�#NST��PAT��P�"PTHJ����E�P rF�V"ART�``%B`�a�bU!REL:�aS�HFT��V!�!�(_�SH+@M$���� ���@N8r����OV9Rq��rSHI%0���UN� �aAYLO����qIl����!�@��@ERV]��1� ?:�¦'�2��%��5��%�RCq��EAScYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba��
5aPo��0�p6OR��MY� `GR��t 2b5n� � ��UPaN�Uu Ԭ")���TOCO!S�1POP ��`�pC�����e��Oѥ`REP�R3��aO�P�b�"ePR�%WU.X1���e$PWR��IM�IU�2R_	S�$VI�S��#(AUD�����Cv" v��$�H���P_ADDR
��H�G�"�Q�Q�Q�БR~pDp1�w H� SZ�a��e�ex�e��SE��r���HS��MNvx ���%Ŕ��OL���p<P��-��ACROlP_!QND_C��ג�1�T� �ROUPT��B_$�VpQ�A1Q�v� �c_��i���i��hx�`�i���i��v�ACk�IOU��D�gfsu<^d�y $|�P�_D��VB`bPR�M_�b�ATT�P_אHaz (��OBJEr��P��[$��LE�#�s>`{ � ��u��AB_x�T~�S|�@�DBGLV���KRL�YHITC�OU�BGY LO: a�TEM��e�0>�+P'�,PSS|�P��JQUERY_F;LA�b�HW��\!�a|`u@�PU�b�PIO��"�]�ӂ�/dԁ=dԁ�� �IWOLN��}����CXa$SLZ�$INPUT_g�$IP#�P��'���SLvpa~��!�\��W�C-�B%�IO^�pF_ASv��$L ��w �F1G�U�B0m!��F�0HY��ڑ����wUOPs� `�� ����[�ʔ[�і"�[PP�SIP�<�іI�2��?�IP_MEMBܿ�i`� X��IP�P�b{�_N�`�����R�����bS�P��p$FOCUgSBG�a~�UJ�Ə� �  � o7JsOG�'�DIS[�J7�cx�J8�7�� Im!�)�7_L�AB�!�@�A��A7PHIb�Q�]�D� J7J\���� �_KEYt� {�KՀLMONa=���$XR��ɀ~��WATCH_����3���EL��}Sy�~���s� �Ю!V8�g� �CTR3�쓥��LG�D� ��R��I�
LG_SIZ���J�q IƖ�I�FDT�IH�_�j V�GȴI�F�%SO��� q �Ɩ���v��ƴ�ǂK�S����w�k�N����E��\���'�*�U�s5��@�L>�4�DAUZ�E�A�pՀ�Dp�f�GH��B�ᢐBOO���� C���PITp���� ��REC��OSCRN����D_p<�aMARGf�`���:���T�L���S��s��W�Ԣ�Iԭ�J{GMO�MNCH�c���FN��R�Kx�PRGv�UF��p0��FWD��HL��STP��V��+������RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28��2��Gh�0PO���������M8�Ģ��EX.��TUIv�I��(�4�@�t�x�J0J�~�P��J0��N�a�#ANA��O"�0�VAIA��dCLE�AR�6DCS_H�I"�/c�O�O&�SI��S��IGN_�vpq�uᛀ�T�d� DEV-�L1LA �°BUW`Ո�x0T<$U�EM��Ł�����A�R��x0�σ\�a�@OS1�2��3�7a�`� �ࠜh�AN%-���-��IDX�DP�2MRO���Գ!�ST��R�q�Y{b! �$E&C+��p.&pA&d���a� L���ȟ%Pݘ��T\Q�UE�`�Ua��_ � �@(��`�����# �MB_PN@ �R`r��R�w�TRIqN��P��BASS\�a	6IRQ6,Ϡ{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?��?RIAt,1ID`�D�� d1��RQQp�rpDSTB
`� 1�F�HAXD2��|�G�LEXCES?R��EMhPa��D�BD4َE�q`�`�F_A�J�C[�Ot�H� K��� \��d�bTf$� ��LI�q��SREQUIRE��#MO�\�a�XDESBU��,1L� M�� �p���P�c��AA,1N��
Q�q�0/�&���-cDC��B�sIN�a?�RSM��Gh� N#B��N�iP�ST9� � 4n��LOC�RI��v�EX�fANG���A,1ODAQ䵗ƞ@$��9�ZMF �����f��"��%u\#ЖVSUP�%Ϡ�FX�@IGGo�� �rq�"��1��#B��$���p%#by���rx���vbPDAT	AK�pE;����R���M��*� t�`MD�qI��)�v� �tĀA�wH�`��tDIyAE��sANSW�P�th���uD��)�b�ԣ(@$`� PC�U_�V6�ʠ�d�PL�Or�$`�R���BD���B�p�����
,1�RR2�E� � ��V�A/A d�$CALI�@��G�~�2��!V��<;$R�SW0^D"��ABC�hD_J�2SE�Q�@�q_Ju3M�
G�1SP�$,��@PG�n�3m�u�3p�@��JkC���2�'AO)IMk@{BCSKP^:ܔ9�wܔ	Jy�{BQܜ�����`_AZ.B��?��EL��YAOCMaP�c|A)��RTьj���1�ﰈ��@1ќ������Z��SMaG��pԕ� ER!���ˀINҠACk�p����b�
n _�������D4�/R��DIU��C�DH�@
�#a�qc$V�Fc�$x�$���`@���b���̂�E�H ��$BELP����!A/CCEL���kA>°IRC_R�p P��T!�$P9S�@B2L  �����W3�ط9� ٶPACTH��.�γ.�3���p�A_��_�e�-Br�`C���_MG�$DD��ٰ��$FW�@�p����γ칲��DE��PPA�BN�ROTSPEEu��O0���DEF>Q����$OUSE_��JPQP�C��JY����-A 6qYN�@A�L�̐��L�MOU�NG̭�|�OL�y�INCU��a�¢ĻB��ӑ�AENCS���q�B������D�IN�I`�����pzC�VE��<���23_U ��b^�LOWL���:�O0��0�Di�B�P�Ҡ� ��PRC����M3OS� gTMOpp�@�-GPERCH  M�OVӤ ����� !3�yD!e�]�6�<�$� ʓA����LIʓ�dWɗ��:p3�.�I�T3RKӥ�AY���� ?Q^���m�b��`p�CQ�� MOM�B?R �0u��D���y�0�̂��DUҐZ�S_�BCKLSH_C ����o�n��TӀ����
c��CLAL�J��A��/PKCH�KO0�Su�RTY�� �q��M�1�q_�
#c�_UMCP�	C����SCL���LMTj�_L�0X����E�� �� � ��m�h���6��PC����H� �P��2�CN@�"XT����CN_��N^C�kCSF����V6�����ϡj���nCAT�SHs�����ָ1����֙���������P�A���_P���_ P0� e���O1u�$x�JG� P{#�OG|���TORQU(� p�a�~����Ry������"_W��^�����4Pt�
5z�
5I;I ;Iz�F�`�!��_8�1��VC��0�D�B�2�1�>	P�?�B�5JR�K�<�2�6i�DBL�_SM�Q&BMD`_sDLt�&BGRV4`
Dt�
Dz��1H_��8�31�8JCOSEKr�EHLN�0hK�5oDt� jI��jI<1�J�LZ1�51Zc@y��1MYqA�H�QBTHWMYTHE{T09�NK23z��/Rn�r@CB4VCBn�CqPASfaYR<40gQt�gQ4VSBt��RN?UGTS���Cq���a��P#���Z�C$DUu ��R䂥э2��Vӑ��Q�r�f$N	E�+pIs@�|� �	$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b��F�c�j�FR�VrhV�ghd��lV�jV�kV��kV�kV�kV�kV�iHrh�f�r�m!�x��kH�kH�kH�kH��kH�iOclOrhOT��nO�jO�kO�kUO�kO�kO�kO�F�F.bTQ���E��egS�PBALANCEl��RLE�PH_'USP衅F��F��FPFULC�3���3��E��1�l�UT�O_p �%T1T2t���2NW������ǡ��5�`�擳�T��OU���� INSsEG��R�REV���R���DIFH��1ٟ��F�1���OB��;C��2� �b~�4LCHWAR���i�ABW!��$MECH]Q�@k�q��AXk�P��IgU�i�� 
���!����7ROB��CR��ͥ�7*�C��_s"T� � x $�WEIGHh�9��$cc�� Ih�.�I9F ќ�LAGK�8qSK��K�BIL?�cOD��U��STŰ�P�; �����
�����
�Ы�L���  2�`�"�DEKBU.�L&�n��POMMY9��NA#�δ9�$D&���q$��� Q ��DO_�A��� �<	���~��L�B$X�P�N��+�_7�L��t�OH  ��� %��T���ѼTx�����TICK/�C�T1��%������!N��c�Ã�R L��S���S�����PRO�MPh�E� $IR� X�~ ���!�MAI�0��j���_9����t�l��R�0COD��FU`�+�ID_" =������G_SUFF�<0 3�O����DO��ِ��R��� �ن�S����!{�����u�	�H)�_FI���9��ORDX� ����36��X�����GR9�S��ZDTD�"�v��ߧ4 *�L_�NA4���K��DEF_I[�K���g�� _���i��Ɠ�š���IS`i �萚���"��e����4�0Bi�Dg����D� �O��LOCKE A!uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ� {����}��v�Ա� ��g������^��� K�Փ����!w�N��P'���^���,`�W�\�[R�7�TE�FĨ �OU�LOMB_u�0��VISPITY��A�!OY�A_FcRId��(�SI�ᄺ�R������3���W�W��0�r�0_,�EAS%���!�& "���4�p�G;� h ���7ƵCOEFF�_Om���m�/�Gd!%�S.�߲CA5�����u�GR` ?� � $R� �X]�TME�$R��s�Z�/,)�ER�T�;�:䗰�  ]�L�L��S�_SVL�($~���0܀��� "SE;TU��MEA��Z��x0�u������ �� � �� ȰI�D�"���!*��&P�H��*�F�'����)3��#���"�5;t`*��REC��:�!7�SK_���� P	�1_USER��,��4���D�0��VEL,2�0��ȯ2�5S�I�|��M�TN�CFG}1� � ���Oy�N�ORE��3��2�0S�I���� ��\�UaX-�ܑPDE�A� $KEY_�����$JOG<EנSVIA�WC�� 1DSWy���
��CoMULT�GI�@�@C��2� 4 ��#t�+�z�XYZ���|�����z� �@_7ERR��� ��S L�-���@��s0BB_$BUF-@X1�7ࡐMOR�� H	�CU�A3�z�1Q��
��3���	$��FV��2��A�bG�� � �$SI�@ G�0VOx B`נOBJE&��!FADJU�#EEGLAY' ���SD�W�OU�мE1PY���=0QT i�0�W�DIR$ba�pےʠDYN�He	T�@��R�^�X����OPWORK}1��,�SYSB9U@p 1SOP�aR$�!�jU�k�PR��2�ePA�0�!�cu� 1+OP��UJ��a'�zD�QIMAG�A1	��`i�IMACr�IN,�bsRGO�VRD=a�b�0�aP �`sʠ� �^uz��LP�B�@��!PMGC_E,�Q��N@�M�rǱ��1Ų7�=q�SL&�~0���$OVSL\G*E��"*E2y�Ȑ�_=p�w ��>p�s���s	�����y�ׯt�#}1� @h�@;���OE�RI#A���
N��X�s�f��{��PL}1�,RT�v�m�ATUSRBT�RC_T(qR��B  �����$ �Ʊ��,�~0� D��`-CSALl`�SA���]1gqXE���%���C�1�J�
���UP(4�����PX��؆�q��3��w� �PG�5�� $SUBࠁ����t�JMP�WAITO��s��L�OyCFt�!D=�CV!F	ь�y���R`�0~��CC_CTR�Q��	�IGNR_P�Lt�DBTBm�P���z�BW)����0UL@���IG�a��Iy�OTNLN��Z�R]a�K� N��`B�0�PE��s���r��f�SPD.}1� L	�A�`g����S��UN�{���r]�R!�`BDLY��2���7�PH_�PK�E��2RET�RIEt��2�b����FI�B� �x���8� 2��0�DBGLV�LO�GSIZ$C�KT�ؑUy#u�D7�_�_YT1@�EM�@C\1�aA����R��D�FC�HECKK�R�P��0����@&�(bLYEc�" PA9�T����P�C߰PN�����ARh�0���Ӯ��PO�BORMATTnaF�f1h���2�S��UXy`	����PLB��4�  �rEITCH���7�9PL)�AL_ � $��XP)B�q� C,2D�!���+2�J3D��� =T�pPDCKyp��|oC� _ALPH�Æ�BEWQo���� ���I�wp � ��b@PAYLOA,��m�_1t�2t���J3AR��؀դּ��laTIA4��5:��6,2MOMCP�Ӡ���������0BϐA�D��������PUBk`R��;���;������z4�` I$PI\Ds�oӓ1yՕ��w�2�w�Z��I��I��I���p����n���y�e`�9S)bT�_SPEED� G�� (�Е��/���Е�`�/�e�>��M��ЕSAMP�6V��/���FЕMO�@ 2@�A ��QP���C��n����� ������LRf`kb�ІE9h�EIN09�� 7S.В9
yPy^�GAMM%S��>�D$GET)bPҺcD]��2
�IBt�q�I�G$HI(0";A��LREXP1A8)LWV M8z)��g���C5�CHKKp]�0�I_��h`eT�� n�q��eT,����� �$�� �1�iPI� RCH_D�313\��30LE�1�1\�o(Y�7 }�t�MSWFL �]M��SCRc�7�@`�&��%n�f�SV���PB``�'�!�B>�sS_SAV&0ct,5B3NO]�C\�C2 ^�0�mߗ�uٍa�� u���u:e;��1���8��D�P������� ��)��b9��e�G@E�3��V�����Ml��� � �YL(��QNQSRlb fqXG�P�RR#dCQ�p� �S:AW70�B �B[�CgR:AMxP�K�CL�H���W�r�(1�n�g�M�!o�� �8F�P@}t$WP�u �P r��P5�R<�R C�R��%�6�`��� (��qsr X��OD�q�Z�Ug�ڐ>D� ��OM#w�J?\? n?�?�?��9�b"۱e�:]�_��� |��X 0��bf��qf��q`���gzf��Eڐ���FbJ�"�ܰ��FdPB���PM�QU�� �� 8L�QCO�U!5�QTHI�H�OQBpHYSY�ES��qUE�`�"�]O���  �P�@L\�UN���Cf�9O�� P��Vu���!����OGRA�ƁcB2�O�tVuI�Te �q:pINFOB�����{�qcB�e�OI�r� (�@SLEQS��q��p�v�gqS���� 4�L�ENABDRZ�PTIONt�����Q�\��)�GCF��G��$J�q^r�B� R���U�g��r�S_ED����� I�F��PK���E'NU߇وAUyT$1܅COPY��P���n�00MN����PRUT8R ��Nx�OU��$�G[rf��e�RGAkDJ���*�X_:@�բ$�����P��W��P��} ��)�}�[EX�YCDR|��NS.��F@r�LG�O�#�NYQ_FREQR�W� �#�h�TsLAe#������ �CRE� s��IF��sNA���%a�_Ge#STA�TUI`e#MAIL�����q t��������ELEM��� �/0<�FEASI?�B��n�ڢ�vA�]� � I�p��`Y!q]�t#A�ABM����E�p<�VΡY�BCASR�Z��S�UZ��0$q���RMS_TR;�qb  ���SY�	�ǡ��$����>C�Q`	� 2� _�TM�� ����̲�@ �A��)ǜ��i$DOU�s]$NLj���PR+@3���r�GRID�qM�BA�RS �TY@�|�O�TO�p��� Hp_"}�!����d�O�P/��� � �p�`P�OR�s��}���SReV��)����DI&0T����� #�	�#�U4!�5!�6!�7!�I8�e�F�2��Ep?$VALUt��%���=b��/��� !;�1�q�����(F_�AN�#�ғ�Rɀ|(���TOTAL��,S��PW�Il��REGEN�1�c�X��ks(��a���`T1R��R��_S� ��1ଃV�����⹂Z�E��p�q��Vr���7V_H��DA�S�����S_Y,1�R4�S�� AR�P2� >^�IG_SE	s��d��å_Zp��C_��~��ENHANC�a�� T ;�8������INT�.���@FPsİ_OVRsP�`p�`��Lv�҂o��7�}��Z�@�SSLG�AA�~�2 5�	��D��S�BĤ�DE�U�����T�E�P���� !�Y��
�J��$2�IL_MC�x r#_��`TQ�`��q���'�B5V�C�P_� 0ڽM�	V1�
V1��2�2�3�3
�4�4�
�!���`� � m�A�2IN~VIBP���1�U2�2�3�3�4�4�A@-�C2�p� MC_YFp+0�0L	1(1d���M50Id�%"FE� S`�R/�@�KEEP_HNA�DD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0�#i�.�#REM�"�$�P�½%�!�(U}�e�$�HPWD  �`#SBMSK|)G��qU2:�P	�COLLAB� �!K5��B�� ��g��pI�TI1{9p#>D� �,�@FLAP��$�SYN �<M�`C�6���UP_DL�YAA�ErDELAh�0ᐢY�`AD�Q���QSKIPN=E� ���XpOfPcNTv�A�0P_Xp �rG�p�RU@,G��:I +�:IB1:IG�9JT�9J@a�9Jn�9J{�9J9<���RA=s� X����4�%1�QB� N�FLIC�s�@J�Ux�H�LwNO_H�0X�"?��RITu��@�_PA�pG�Q�S ��^�U��W���LV�d�NGRLT �0_q��O�  " ��OS���T_JvA V	�A�PPR_WEIG=H�sJ4CH?pvT�OR��vT��LOO��]�+�tVJ�е�ғaA�Q�U�S�XOB'��'���J2P���
7�X�T�<a43DP�=`Ԡ\"<a�q\!��RsDC��L� �рER��R�`� �RV�p�jr�b�RGE��8*��cN�FLG�a�Z����SPC�s�U�M_<`^2TH2�NH��P.a 1�� m`EF11��� lQ �!#� <�p3AT� g�S�� Vr�p�tMq�Lr���HOMEwr�t2'r�-?Qcu��w3'r���P����w4'r�'�@9�K�]�o����w5'r뤏��ȏڏ����w6'r�!�3�E�W�i�{��w7'r힟��Pԟ����w8'r��@-�?�Q�c�u��uS$0
�q�p�� sF��`ala�!`P����a�`/���-�IO[�M�I֠��qPOW=E�� ��0rZa*��� �5ވ�$DSB GN�AL���0Cp���laS2323�� Ɍ~`��� / ICEQP��PEp��5PsIT����OPBx0ޣ�FLOW�@TR`vP��!U���CU�M��UXT�A��w�ERFAC�� U���ȳCH��� tQ  _��>�Q3$����OM���A�`T�P#UPD�7 A�ct�T��UE�X@�ȟ�U EFA8: X"�1RSPT��ѧ��T ��PPA��0o񩩕`EXP�IAOS���)ԭ�_�0��%��C�WR�A���ѩD�ag֕`ԦFR�IENDsaC2UFx7P����TOOL���MYH C2LENGTH_VTE���I��Ӆ$SE�����UFINV_t���RGI�N{QITI5B��Xvl��-�G2-�G17� w�SG�X��_��UQQD=#���AS��d�~C�`��q�� ��$$C/�S�`������ Ȱ����V�ERSI� ��]Ȱ�5��I���������AAVM_�Y�2 �� 0  �#5��C�O�@�r� )�r�	 ������ ���������� ������
?QYf�BS���1��� <- ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O��O�O�OiCC�@XgLMT��C�7  ��DIN�O�A\�Dq�EXE�HPV_��ATQz
���LARMRECOV �RgLMDG *��5�OLM_IF' *��`d�O�_ �_�_�_j�_'o9oKo<]onm, 
��o db��o�o�o�o^���$� z, A  � 2D{�PPIN�FO u[ @�Vw������� �`�������*� �&�`�J���n�����DQ����
��.� @�R�d�v����������a
PPLICATf��?�P��`�Handl�ingTool �
� 
V8.3�0P/40Cpɔ_LI
883���ɕ$ME
F�0G�4�-

�398�ɘ�%�z��
7DC3x�ɜ
�Noneɘ�Vr���ɞ@�6d� Vq_A�CTIVU��C죴�MODP���C��I��HGAPONp���OUP�;1*�� i�m�����Қ_����1�*�  �@���� ����Q���Կ濸@�
����� g���5�Hʵ�l�K�HTTHKY_��/�M�SϹ��� ������%�7ߑ�[� m�ߝߣߵ������� ���!�3��W�i�{� ������������� �/���S�e�w����� ����������+ �Oas���� ���'�K ]o������ ��/#/}/G/Y/k/ �/�/�/�/�/�/�/�/ ??y?C?U?g?�?�? �?�?�?�?�?�?	OO uO?OQOcO�O�O�O�O �O�O�O�O__q_;_ M___}_�_�_�_�_�_�_kŭ�TOp��
��DO_CLEAN�9��pcNM  !{衮o�o�o�o�o���DSPDRY�Rwo��HI��m@ �or����������&�8�J���MAXݐWdak�H�h��XWd�d���PL�UGGW�Xgd��P�RC)pB�`�k�aS�Oǂ2DtSEGF0�K� �+� �o�or����������%�LAPOb�x��  �2�D�V�h�z�����య¯ԯ�+�TOT�AL����+�USE+NUO�\� e�A��k­�RGDISPWMMC.���C6�&z�@@Dr\�OMpo��:�X�_STRI�NG 1	(�
��M!�S��
��_ITEM1Ƕ  n����� �+�=�O�a�sυϗ� �ϻ���������'��9�I/O S�IGNAL���Tryout M�odeȵInp�y�Simulat{eḏOut��OVERRLp� = 100˲In cycl��̱Prog A�bor��̱u�S�tatusʳ	H�eartbeat�ƷMH Fauyl	��Aler� L�:�L�^�p����8������ Scû Saտ��-�?�Q�c�u� ���������������);M_q��WOR.�û���� ��+=Oa s�������8//'.PO���� M �6/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?H"DEVP.�0d/�?O *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�J_\_n_PALT 	��Q�o_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o�_GRIm�û9q�_ as������ ���'�9�K�]�o� ������'�R	�݁ Q����)�;�M�_� q���������˟ݟ����%�7�I�ˏPREG�^����[����� ͯ߯���'�9�K� ]�o���������ɿۿ��O��$ARG_�� D ?	����0�� � 	$O�	+[D�]D��O�e��#�SBN_CON?FIG 
0˃����}�CII_SAVE  O������#�TCEL�LSETUP �0�%  OME�_IOO�O�%M�OV_H������R�EP��J��UTOoBACK�����FRA:\�o� Q�o���'�`��o���� �� f�o������*�!�3�`�Ԉ��f���������� o�{��&�8�J�\�n� ��������������� ��"4FXj| �������ׁ  ��_i�_\�ATBCKCTL�.TMP 6.V�D GIF .TP D_q���N.E#��f�IN�I�P�Օ�c�MESSAG�����|8��ODE_D�����z��O�0�c�P�AUSM!!�0� ((O3�U/g+ Q/�/u/�/�/�/�/�/ �/�/)??M?;?q?7�0$: TSK  �@-��T�f�UPDT���d�0
&XW?ZD_ENB����6STA�0��5"��XIS��UNT �20Ž� � �	 �/� 0/� 3���;:: �n�o� U@�?��o�}O�O�O�O��O�O�O"_�?7AME�T߀2CMPTA>��oH=	��=�R�^�?�I��>Ë�_�_4_A�XSCRDCFG� 1�6�Ь�Ź��_�_o@o(o:oLo��o�Q�� �_�o�o�o�o�o�o]o �o>Pbt��0�o9�i�GR<@MX/�s/NA�/�s	i��v_ED��1�Y� 
 ��%-5EDT-��'�GETDA3TAU�o�9��?�(j�H�o�f�\�ּA��  ���2 �&�ȏE�D���~� ŏ׏m����3��&� �J�\�ߟJ�����9�ǟ�4���ϯ�\�����]�o�����5 N������\�w��)�;�ѿ_��6ϊ�g� ��\�CϮ���ϝ�+��7��V�3�z�\��@z�����i����8������]���F� �ߟ�5����9~������]����Y�k�����CR�!ߖ� ��W�q���#�5���Y���p$�NO_DEL���rGE_UNU�SE��tIGAL�LOW 1���(*SYS�TEM*S	$SERV_GR��V� : REG�q$�\� NUM�
<��PMUB U�LAYNP\PMPAL�>CYC10#6� $\ULSU`�8:!�Lr~�BOXORI��CUR_��PoMCNV��10L�T4DL!I�0��	����B N/`/r/�/�/�/�/�/����pLAL_OU�T �;���qW?D_ABOR=f��q;0ITR_RT�N�7�o	;0NON�S�0�6 
HCC�FS_UTIL s#<�5CC_@�6A 2#; h� ?�?�?O#O�]CE�_OPTIOc8�qF@RIA_IIc f5Y@�2�0�F�Q�=2q&}ނA_LIM�2�.� ��P��]B���KX�P
�P�,2O�Q��B�r�qF�PQ5T1)TR�H�_:JF_PA�RAMGP 1�<g^&S�_�_�_��_�VC�  C��d�`�o!o`��`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?���2HE ONFI�� E?�aG_P�1#; ���o 1CUgy�a�KPAUS�1�yC ,���� �����	�C�-� g�Q�w���������я4���rO�A�O�H~�LLECT_�B1�IPV6�EN. QF܍3�NDE>� ��G�71234567890���sB�TR����%
 	H�/%)����� ��W���0�B���f�x� ��㯮���ү+���� �s�>�P�b������� ���ο��K��(Ϡ:ϓ�^�|��B!F�� �I|�IO #��<U%e6�'��9�K���TR�P2$���(9X�t�Y޼`�%�̓ڥH��_MO-R�3&�=��i� �A�$��H�6�l�Z���~S��'�=�r_A? �a�a`��@K��RʭdP��)F�haÃ-�_�'�9�%
@�k��G� ��%Z�^%��`�@c.��PDB��+���cpmidbg���	3 :�  %' QU��p��N�' ��@���)����]�`@�s<�^��@�bsg�$�.s�fl�q��u�d1:��:J��D�EF *ۈ��)��c�buf.�txt����_�L64FIX ,������l/[Y/�/ }/�/�/�/�/
?�/.? @??d?v?U?�?�?�?��?�?�?,/>#_E -���<2ODOVO�hOzO�O6&IM��.zo�YU>���d�l
�IMC��2/��b��dU�C��20�M�QT:Uw�Cz  �B�i�Aep�?����?2]8�+;�CG�A�n&`w�XQ�á�@/
?�f�9��SD�%�A�Mes]C �"A:�R@�q�u=7m�E\C g��kJ��22o�D|���.U ���C�C-����
�xObi�D4cdv`D��`/��`v`s]E�D D��` E4�F�*� Ec��F�C��u[F���E���fE��fF�ކ3FY�F��P3�Z��@�3�3 ;��>L̩��Aw�n,a@��@e�5Y���a���`�A��w�=�`<#����
��?�ozJRS�MOFST (X�,bIT1��D @3��
д����a���;��bw?����<�M�NT�EST�1O�CR�@�4��>VC5`A�w�Ia+a�aORI`mCTPB�U�C�`�4���r��:d�T���qI?�5��q�T_�PROG 	��
�%$/ˏ�t���NUSER  �k�������KEY_?TBL  �����#a��	
��� !"#$%&'�()*+,-./���:;<=>?@�ABC�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~��������������������������������������������������������������������������������͓���������������������������������耇���������������������9�����LCK�
�<���STAT/��s�_AUTO_DO� �	�c�IND�T_EN�PR���R�pqn�`�T2����ScTOr`���XC��� 26���8
�SONY XC-�56�"b����@���F( А=�HR50w����>�P�7b�t�Af!f����ֿ� Ŀ� ���C�U�0�yϋ�f� ���Ϝ��������-���TRL��LET�Eͦ ��T_S�CREEN >��kcs����U�MMENU {17�� <� ����w�������� �K�"�4��X�j�� �����������5�� �k�B�T�z������� ��������.g >P�t���� ��Q(:� ^p����/� �;//$/J/�/Z/l/ �/�/�/�/�/�/�/7? ? ?m?D?V?�?z?�? �?�?�?�?!O�?
OWO .O@OfO�OvO�O�O(y~��REG 8�y�����`�M�ߎ�_?MANUAL�k��DBCO��RIG�Y�9�DBG_ER�RL��9�ۉq���_�_�_ ^QNOUMLI�pϡ�p�d
�
^QPXWO_RK 1:���_�5oGoYoko}oӍDBwTB_N� ;������AD�B_AWAYfS^�qGCP 
�=�p�f_AL�pR��bbR�Y�[�
�WX_�P +1<{y�n�,�%o`c�P��h_M���ISO��k@L��sOoNTIMX��
����vy
��2sM?OTNEND�1t�RECORD 1�B�� ���sG�O�]�K��{�b�� ������V�Ǐ�]�� ��6�H�Z������� ��#�؟������2� ��V�şz�������� ԯC���g��.�@�R� ��v�寚�	���п� ��c�χ�#ϫ�`�r� �ϖ�Ϻ�)ϳ�M�� �&�8ߧ�\�G�Uߒ� ߶�����I������4�� �p7�n���� ����������"� ��F�1���|������ ��[�����i���B�Tf���bTOL�ERENC�dB��'r�`L��^PCS�S_CCSCB �3C>y�`IP�t }�~�<�_` r�K�����/�{��5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O��O�O�O�O_�~�L5L� D��&qET|�c�a C[�C��PZP^r_ A�� p� �sp�x�QGPt[	 A�p�Q�_�[? �_�[oU�p�P�pSB�V�c�(a�PWoPio{h+�o�X�o�oY��[	r�h�LUwN2E*��5��:�N7�2ܘ��c��aD@VB���|�G���+��K� �otGhXGr�So�����eB   =���Ͷa>�tYB��� �pC�p�q�aA"�H�S�Q-��q����ud�v�����AfP w` 0���D^P���p@�a
�QAXTHQ�z�a a"W>� �a9P��b�e :�L�^�h�Hc�́PQ�RFQ�PU�z�֟ �o\^��-�?��c��u����zCz��ů�b2�Щ�RD�;Rl��p����� �S̡0��]�0�.��@���EQ�p��F�X� ѿUҁп�VSȺ�NSTCY 1E��]�ڿ��K� ]�oρϓϥϷ����� �����#�5�G�Y�k��}ߏߒ��DEVI�CE 1F5� MZ�۶a��	� ��?�6�c���	{䰟�����_HNDGD �G5�VP���R�LS 2H�ݠ��/��A�S�e�w����� ZPARAM I��FgHe�RBT [2K��8р<�߬WPpC�C��,`¢�P�Z�����%>{�C*  �2�j�MTLU,`"nPB , s���M� }�gT�g��
B��!�bcy�[2Dch z����/���/gT#I%D��CǓ` b!�R��A���A,��Bd���A��P��_C14kP�!2�C��$Ɓ��]�ffA�À���B�� �| �0��/�/�T (��5 4a5�}%/7/d?/ M?_?q?�?�?�?�?�? O�?OO%O7OIO�O mOO�O�O�O�O�O�O �OJ_!_3_�_�_3�_ �_�_�_�_o�_(oo Lo^oЁ=?k_IoS_�o �o�o�o�o�o�o #5G�k}�� �����H��1� ~�U�g�y�ƏAo�Տ ���2�D�/�h�S��� go����ԟ����ϟ� ��R�)�;���_�q� ���������ݯ�<� �%�7�I�[�m����� ����}�&��J�5� n�YϒϤϏ��ϣ�ѿ ������F��/�A� ��e�w��ߛ߭����� ����B��+�x�O�a� �����������,� ��%�b�M���q����� ����������L #5�Yk}�� � ��61 CUg����� ���	//h/���/ w/�/�/�/�/�/
?�/ .?@?I/[/1/_?q? �?�?�?�?�?�?�?O O%OrOIO[O�OO�O �O�O�O�O&_�O_\_ 3_E_W_�_?�_�_�_ �_�_"ooFo1ojoE? s_�_�om_�o�o�o�o �o0f=Oa �������� ��b�9�K���o��� Ώ��[o��(��L��7�I���m������$�DCSS_SLA�VE L��}�ё���_4D  љ�~�CFG Mѕ���������FRA:\ĐL�-�%04d.CS�V��  }�� ����A i�CHq�z�������|�����  �����Ρޯ̩<ˡҐ-��*�����_CRC_OUT N������_FSI ?њ ����k� }�������ſ׿ ��� ��H�C�U�gϐϋ� �ϯ��������� �� -�?�h�c�u߇߰߫� ����������@�;� M�_��������� ������%�7�`�[� m�������������� ��83EW�{ ������ /XSew�� �����/0/+/ =/O/x/s/�/�/�/�/ �/�/???'?P?K? ]?o?�?�?�?�?�?�? �?�?(O#O5OGOpOkO }O�O�O�O�O�O _�O __H_C_U_g_�_�_ �_�_�_�_�_�_ oo -o?ohocouo�o�o�o �o�o�o�o@; M_������ ����%�7�`�[� m��������Ǐ��� ���8�3�E�W���{� ����ȟß՟��� �/�X�S�e�w����� ���������0�+� =�O�x�s��������� Ϳ߿���'�P�K� ]�oϘϓϥϷ����� ����(�#�5�G�p�k� }ߏ߸߳����� ��� ��H�C�U�g��� ����������� �� -�?�h�c�u������� ��������@; M_������ ��%7`[ m������ �/8/3/E/W/�/{/ �/�/�/�/�/�/?? ?/?X?S?e?w?�?�? �?�?�?�?�?O0O+O =OOOxOsO�O�O�O�O��C�$DCS_C�_FSO ?�����A P �O�O_ ?_:_L_^_�_�_�_�_ �_�_�_�_oo$o6o _oZolo~o�o�o�o�o �o�o�o72DV z������ �
��.�W�R�d�v� ������������ /�*�<�N�w�r����� ����̟ޟ���&� O�J�\�n��������� ߯گ���'�"�4�F� o�j�|�������Ŀֿ ������G�B�T��O_C_RPI�N_ jϳ����ς��O���ϰ1�Z�U��NSL��@ &�h߱���������"� �/�A�j�e�w��� �����������B� =�O�a����������� ������'9b ]o������ ��:5GY� }������/ //1/Z/U/g/y/�/ �/�/�/�/�/�/	?2? -???Q?z?u?��ߤ� �?�?�?�?OO@O;O MO_O�O�O�O�O�O�O �O�O__%_7_`_[_ m__�_�_�_�_�_�_ �_o8o3oEoWo�o{o �o�o�o�o�o�o /XSew�� ������0�+� =�O�x�s��������� ͏ߏ���'�P�K��]�o����� �PRE_CHK P����A ��,8��2��� 	c 8�9�K���+� q���a�������ݯ� ͯ�%��I�[�9�� ��o���ǿ��׿��� )�3�E��i�{�Yϟ� �Ϗ����������� -�S�1�c߉�g�y߿� �߯����!�+�=��� a�s�Q������� ��������K�]�;� ����q����������� ��#5�Ak{ ����� �CU3y�i� �����/-/G /c/u/S/�/�/�/�/ �/�/??�/;?M?+? q?�?a?�?�?�?�?�? �?�?%O?/Q/[OmOO �O�O�O�O�O�O�O_ �O3_E_#_U_{_Y_�_ �_�_�_�_�_�_o/o oSoeoGO�o�o=o�o �o�o�o�o= -s�c���� ���'��K�]�wo i���5���ɏ������ ��5�G�%�k�}�[� ������ן�ǟ�� ��C�U�o�A�����{� ��ӯ����	��-�?� �c�u�S�������Ͽ ῿�����'�M�+� =σϕ�w�����m��� ���%�7��[�m�K� }ߣ߁߳��߷���� !���E�W�5�{��� ����e�������	�/� �?�e�C�U������� ��������=O -s����]� ���'9]o M������� /�5/G/%/k/}/[/ �/�/��/�/�/�/? 1??U?g?E?�?�?{? �?�?�?�?	O�?O?O OOOuOSOeO�O�O�/ �O�O�O_)__M___ =_�_�_s_�_�_�_�_ o�_�_7oIo'omoo ]o�o�o�O�o�o�o !�o1W5g�k }������/� A��e�w�U������� я��o����	�O� a�?�����u���͟�� ���'�9��]�o� M���������ۯ��ǯ �#�ůG�Y�7�}��� m���ſ�����ٿ� 1��A�g�E�wϝ�{� ��������	�߽�?� Q�/�u߇�e߽߫ߛ� �������)���_� q�O��������� ����7�I���Y�� ]��������������� !3WiG�� }����%� A�1w�g�� ����/+/	/O/ a/?/�/�/u/�/�/�/ �/?�/9?K?�/o? �?_?�?�?�?�?�?�? O#OOGOYO7OiO�O mO�O�O�O�O�O_�O 1_C_%?g_y__�_�_ �_�_�_�_�_o�_+o Qo/oAo�o�owo�o�o �o�o�o);U__ q������ ��%��I�[�9�� ��o���Ǐ�����ۏ !�3�M?�i��Y��� ����՟�ş���� A�S�1�w���g�����������ӯ�+�=���$DCS_SGN� QK�c��7�m� 17-�JAN-19 13:15   O��l�4p�08:38�}����� N.DѤ����������h�x,rWf*�σ�^M��  �O�VERSION� [�V3�.5.13�EF�LOGIC 1R�K��  	���P�?�P��N�!�PROG_E_NB  ��6����o�ULSE  �TŇ�!�_AC�CLIM�����Ö��WRSTgJNT��c��K�EMOx̘��� ���INIT S.��G�Z���OPT_S�L ?	,��
 	R575��VY�74^�6_�7_�+50��1��2_�@�����<�TO  �Hݷ���V�DE�X��dc����P�ATH A[�A�\�g�y��HC�P_CLNTID� ?��6� �@ȸ����IAG_�GRP 2XK�� , `���� �9�$�]�H������1234?567890����S�� |�������8!�� ��H؀��;�dC�S��� 6�����. �Rv�f�� H��//�</N/ �"/p/�/t/�/�/V/ h/�/?&??J?\?�/ l?B?�?�?�?�?�?v? O�?4OFO$OjO|OO E��Oy��O�O_�O 2_��_T_y_d_�_,
�B^ 4�_�_~_ `Oo�O&oLo^oI��T jo�o.o�o�o�o�o  �O'�_K6H�l �������#� �G�2�k�V���B]��?�  ��3:/3\E�������޾���aƁD|�Ο@㈙D�"���Ƈ����(���L�B\ډC4  ��E2���c >���:�����ߟʟܟ����CT_CON�FIG Y��|Ӛ�egU����STBF_TTS��
��b����Û�:u�O�MAU��|�~�MSW_CF6��Z��  �OCoVIEW��[ɭ������-�?�Q� c�u�G�	�����¿Կ ������.�@�R�d� v�ϚϬϾ������� ߕ�*�<�N�`�r߄� ߨߺ��������� &�8�J�\�n���!� �������������4��F�X�j�|����RC£\�e��!*�B^�� ����C2g{��SBL_FAUL�T ]��ި�G�PMSKk��*�TDIAG ^:��աI��UD�1: 6789012345�G�BSP�-?Qcu �������/@/)/;/M/tJ��
�@q��/$�TRECP��

��/ ?"?4?F?X?j?|? �?�?�?�?�?�?�?O�O0OBOi/{/xO�/U�MP_OPTIO1Nk���ATR¢l�:�	�EPMEj��O�Y_TEMP  È�3B�J��P�AP�DUNI�m�Q��YN_B�RK _ɩ�E�MGDI_STA�"U�aQSUNC_S1`ɫ �FO�_�_
�^
�^dpOoo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{�E���� �y�Q��� �2�D� V�h�z�������ԏ ���
��.�@�R�d� �z�������˟�� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i������� ��ÿݟ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�{�iߗߩ߻�տ�� ����'�9�K�]�o� ������������� �#�5�G�Y�s߅ߏ� ����i������� 1CUgy��� ����	-? Qk�}������� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?u? �?�?�?��?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_m?w_�_�_�_�? �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9Ke_W ����_�_��� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�]oy������� �ӟ���	��-�?� Q�c�u���������ϯ ����)�;���g� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�_�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�W� E�s������ߧ����� ��'9K]o �������� #5O�a�k}� E������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-?G Yc?u?�?�?��?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_Q?[_m__ �_�?�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ I_Sew��_�� �����+�=�O� a�s���������͏ߏ ���'�A3�]�o� ������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 9�K�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� �����ߑ�C�M�_� q߃ߝ��߹������� ��%�7�I�[�m�� ������������� !�;�E�W�i�{��ߟ� ����������/ ASew���� ���3�!O as������� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?+=G?Y?k?!?� �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	_#?5??_ Q_c_u_�?�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o -_7I[m�_ �������� !�3�E�W�i�{����� ��ÏՏ����%/� A�S�e�q������� џ�����+�=�O� a�s���������ͯ߯ ����9�K�]�w� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������'� 1�C�U�g߁��ߝ߯� ��������	��-�?� Q�c�u������� ����m��)�;�M�_� y߃������������� %7I[m �������� !3EWq�{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/�/+?=?O? i_?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O?� �$ENETM�ODE 1aj5��  
0054_F[P�RROR_PRO/G %#Z%6�_��YdUTABLE  #[t?�_�_�_�gdRSEV_NU�M 2R  ��-Q)`dQ_AU�TO_ENB  qPU+SaT_NO>a� b#[EQ(b�  *��`��`��`��`4`+�`�o�o�oZdHIS%c1+P�Sk_ALM 1c.#[ �4�l0+�o;M_q���o_b``  �#[aFR�zPTC�P_VER !�#Z!�_�$EXTLOG_REQ�fs�Qi,�SIZ5��'�STKR�oe��)�TOL  �1Dz�b�A '�_BWD�p��Hfܻ�D�_DI�� dj5SdDT1KRņSTEPя�P>��OP_DOt�Q�FACTORY_�TUN�gd<�DR_GRP 1e#YNad 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ� ԟ���1��U�@�y� d�v�����ӯ����LW
 I�4y�,��tۯ�j�U���~y�B�  B୰}���$  A@��s�@UUUӾ����|���E�� E�`�F@ F�5U�/�,��L���M���Jk�L�zp�JP��F�g�f�?�  �s��9�Y9}��9��8j�
�6��6��;��m����y �_� �� Q�(������[FEATU�RE fj5���JQHand�lingTool� � "
P�English� Diction�ary�def.4D St��ard�  
!� hAnal�og I/OI� � !
IX�gle ShiftI��d�X�uto S�oftware �Update  �rt sѓ�mat�ic Backu�p�3\st���ground �Edit��fd�
Came�ra`�Fd�e��CnrRndIm����3�Commo�n calib �UI�� Ethe��n��"�Moni�tor�LOAD�8�tr�Reli�aby�O�ENS�D�ata Acqu�is>��m.fd~p�iagnos���]�i�Docume�nt Viewe�J��870p�u�al Check Safety*�� cy� �hanc�ed Us��Fr�����C �xt.� DIO :�fi�� m8���end.��ErrI�L��S�������s  t KPa�r[�� ����J944F�CTN Menur��ve�M� J9l��TP InT�fa}c{�  744���G��p Mask� Exc��g�� �R85�T��Pr�oxy Sv�� � 15 J�ig�h-Spe��Sk}i
� R738�����mmunic��ons�S R�7��urr�T�d�0�22��aю�con�nect 2� {J5��Incr���stru,Қ�2 �RKAREL Cmd. L��{ua��R860h�Run-Ti��E[nvL�oa��KU�el +��s��S�/Wѹ�7�Lic�ense���ro�du� ogBoo�k(System�)�AD pMACROs,��/Offs��2�N�Ds�MH�� ����MMRC�?���ORDE� ech/Stop��t? �7 84fMi$�|� 13dx��]еи׏���Modz�w/itchI�VP��t?��. sv��2Optm�8�2��fil��I ��2�g 4 !+ulti-T������;�PCM f3unY�Po|���x4$�b&Regi� �r �Pri��F�K+7���g Numo SelW  �F�#�� Adju���60.��%|�� fe���&tat�u�!$6���%�� � 9 J6R�DM Robot�)�scove2� w561��RemUz�n@� 8 (S�>F3Servo��ҩ�)SNP�X b�I�\dcys�0}�Libr1Ӟ�H� �5� �f�0��58��Soz� tr�ssag4%^G 91�p ��d&0���p/I���  (ig TMI�LIB(MӋ�Fi3rm����gd7���Ns�Acc����0��XATX�Heln���*LR"1��Swpac�ArquzПimulaH��� �Q���Tou�Pa���I��T��c��&���ev. f.s�vUSB pYo��"�iP�a���  r"1Unexcept��`0i$/�����H59� VC"&�r��[6���Px{��RcJPRIN�V��; d T@�TS?P CSUI�� �r�[XC��#We�b Pl6�%d -c�1R�@4d��8���I�R66?0FVx�L�!FVGridK1?play C�lh�@����5RiR�R.�@���R-35iA����Asciip���"��� 51f��cUpl� � (�T����S��@ri�tyAvoidM� �`��CE��rk��Col%�@�GEuF� 5P��j}P�����
 B�L�t� 1+20C C� o�І!�J��P��y��� o�=q�b @DCS b ./��c��O��q���`�; ���qc�kpaboE4�DH�@�OTШ�main� N��1.�H��a�n.��A> aB!F#RLM���!i ��пMI Dev�  9(�1� h8j��spiJP��� �@��A"e1/�r���!hP� M-2� i��߂�^0i�p6�PC���  iA/'�Passwo�qT��ROS 4����qe�da�SN��Cli ����G6x Ar��G 47�!���5s��DER��Tsup�>Rt�I�7 (M��a�T2DV�
�3?D Tri-���H&��_8;�
�A�@�Def?����B�a: deRe p 4t0��e�+�V��st64MB DwRAM�h86�΢FRO֫0�Arc� visI�ԙ�yn��7| ), �b�Heal�wJ�\=h��Cell`��p� �sh[��� tKqw�c� - ��v���p	VCv�ty�y�s�"Ѐ6�ut��v�m���xs ���TD_0��J�,m�` 2��a[�>R� tsi�MAILYk�/F2�h���>�� 90 H��F0�2]�q�P5'���Ta1C��5����FC���U�F9�GigE�H�S�t�0/A� i�f�!2��boF�d�ri=c �O�LF�S����" H=5k�OPT ���49f8���cr�o6��@��l�Ap�A�Syn.(RS�S) 1L�\1y�rH�L� (2x5�5�d��pCVx9����es�t�$SР��> \p�ϐSSF�e$�tex�D o���A�	�� BP���a�(R00�Qirt��:���2)�D��1�e�VK�b@l Bui, n��WAPLf��0b��Va�kT�XCGM�ċD��L����[CR1G&a�YBU��Y�KfL��pf��k�\sm�ZTAf�@��
��Bf2�и��V#��s���� r���CB����
f���WEB��!��
���T�p���DT�&4 Y�V�`��EH����
F�61Z��
�R=2L�
�E (Np��F�V@�PK�B���#��Gf$1`?G���H�р�?I�e ����LDh�L��N��7\s@����`���M��d�ela<,��2�M.�� "L[P��`�?��_�%�����S���-F�TSO�W�J57��VGF܋|�VP2֥ 5\b�`0&�cV:����T;T� �<�ce�,?VPD��$�
T;F��DI):�<I�a\so<��a-�6Jc6s6�4L��M�V9R�h���Tr@i�� ���5�` �f�@ �������P
� ���|�`��Img PH��[l��I/A � VP�S��U�O�w��!%S�Skastd�pn)ǲt�� SW_IMEST�BFe�300��-Q� �_�P8B�_�Rued�_�T��!�_�S ��_bH'573o2c2��-o�NbJ5N�Iojb)�Cdo�cxE��o�_�lp� �o�TdP�o�c�B�or �2.rٱ(Jsp�EfrSEo�f1�}�r�3 RGoeELS��sL����s������B	��S\ $�F�r�yz�ftl�o~�g �o���������?�����P  �n�&�"�l ��T�@<�^��Y���e�u8Z���alib��Γ��ɟ3����埿�\v ��e\c��6�Z�f�T�v�R� VW���8S��UJ�91����i�ů[c9�1+o�w8���847�:��A4�j���Q��t6�m���vrc�.����HR���oqt�0ݿ��  ��28ޯ�460�>e3S0L�97���U�ЄϦ�60.� g�Ѐ��+��'�ܠ�Ϻ�8Lco��DM߱U"������ߕpi�߲T! L��na;�� �� �u%��ⅰI���loR�d��1a590gϱŭ���95�ϔ�	R����1��?��o�@#��1A�/���vt{UWeǟ���ￇ7�3[���7�ρ�C �W��62K�=fR���8��������d����2�ڔ����@��@" "http�����t7 ��� v R7��78����4�� ��TTPT�#	��eGPCV4/v߀�j�&Q�Fa7��$N�0�/2�rIO�)/;/M/6'.sv3�64i�oS�>l? torah?*�8|`�?��AM/�?
?�?.?0�k/��1 J`O��� ,O�tro��`�[P��OB4c.K?��g'�)�24g?�� c(B�Od�\iO�A5sb�?U_�?vi �/i��/�/Wn��`�o%�Fo�4l�$of8��oXF I)xo�cgmp\7��mp���duC��lh����o�(A�_Bt� �o]6P���m�I?�w�@���nIaO��4*O0wip�%P�?"�bsg?� ]7�YEM���8woV�J�/ե11?o��D�Ms�BC��7�J�\���(�52�XFa# AP�ڟ<�v�`/�şaqs����/�Of��1�9�VRK���ph�ք3H5+�=�IN/¤�SkiW�/�IF`��_�%��fs�$I�O�l����"<�0�$�`����\jԿz5�bO�vrouς�3(�ΤH (DϮ��? sG��|��F�Ou����@���D)O��*�3P $�FӅ�k��ϻ���럊�� �PL��ʿ��pgbox�ߦebo�&��Sh �>�R.�0w1T{����fx6�� P��D��3��#_I�\m;YEe�OԆMp�hxW�=Ete,����dct\���O$k R������Xm*��փro3��D�l�j�9��V'�  �FC���|@�ք <f?6KARE0�_��~ (Kh��.c1f���WpoO�_K�up��a���H/�j#- Eqd/�84���$qu�o��/  o2o?Vo<�7C�)��s�NJԆ�|?�3l\sy�?�40�?Τ�wio�u]?�w58�?,F�$OJ�
?Ԇ�"io�!�V��u&A���PR�ߩ5, �s��v1\  ?H552B�Q�21p0R7�8P510.R0�  nel �J614Ҡ/W?ATUP��d�8P545*�H8R6���9VCAM:�q97PCRImP\1�tPUIF�C8Q28  ingsQy0��,4P P63P @P P�SCH��DO�CVڀD �PCSUȾ��08Q0=PqpVEIOCr��� P�54Pupd�PR�69aP���PSET�pt\hPQ`Qt�8P�7`Q�!MAS�K��(PPRX�Y���R7B#POCO  \pppb36���PR�Q��b1P�d60Q$cJ539�.eHsb��vL�CH-`(�OP[LGq\bPQ0]`:��P(`HCR���4`S�aund�PM�CSIP`e0aPle5r=Ps�p(`DSW�  �  qPb0`�aPa��(`PRQ`Tq�RE`(Poas601P<cPCM�P�HcR0@q\j23�b�V�`E`�S`UPvisP`E` c�`UP�cPRS	a�bJ699E`sFRDmPs�RMCN:eH93<1PHcSNBARa�r7HLB�USM�qc�Pg52�fHTC<IP0cTMIL�e"P4�`eJ �PA�PdSoTPTX6p967PTEL�p��P�`�`4
Q8P8$Q48>a"PPX�8P95�P`[�s95qqbUEC-`wF
PUFRmP�fahQCmP90ZQV�CO�`@PVIP�%�537sQSUI�zVSX�P�SWEB�IP�SHTTIPth�rQ62aP�!tPGL���cIG؁�`c�wPGS�eIRC%�N�cH76�P�e Q��Q|�Ror��R51`P s:P�P,t53=PR8u8=Py�C�Q6]``�b�PI��q52]`sJ56E`s���P�DsCL�qPt5�\�rd�q75UP cR�8���u5P sR55]`,s� P8s��P��`CP�PP�SJ77.P0\o�6��cXRPP�cR6�ap�`��QtaT�79P`�6�4�Pd87]`�d90P0c��=P,���5�Y9ta�T91P� ���1P(S���Qpaiv�P06=P- C�PF�T	���!aLP PsTS�pL�CAB%�)I БIQ` ;�H��UPPaintPMS��Pa��D�IP|�ST�Y%�t\patPT�O�b�P�PLSR7�6�`�5�Q��WaN�N�Paic�qNN�E`�ORS�`�cR�681Pint'�FCB�P(�6x�-W`iM�r��!(`OBQ`�plug�`L�ao;t �`OPI-���rPSPZ�PPG�Q�7�`73ΒPRQ�ad�RL��(+Sp�PS��n�@��E`�� �PTS�-�� W��P�`a�pw�`��P`cFV9R�PlcV3D%�l��PBVI�SAPL��Pcyc+PAPVv1�pa_�CCGIP� - U��L�Pr;og+PCCR�`�JԁB�P �PԁK=�C"L�P��p��(h��<�P��h�̱�@g�Bـ
TX�%���7CTC�ptp��2��P927"0ҝPs�2�Qb��TC-�rm�t;�	`#1ΒTC�9`HcCTE�Per�j�EIPp.p/�Ep�P�c��I�use��-Fـvrv�F%��ăTG�P� CP��%�d� -h�H-�Tra��PCTI�p��TL� TRS���p�@Pנ��IP�PTh�M%��lexsQTMQ`vGer, �p�SC:�8��F��Pv\e�PF�IPSV"+�H�$cj�vـtr�aCTW-����CPVGF-��SV{P2mPv\fx����pc�b��e��bVP4�fx_m��-��S�VPD-��SVPF.�P_mo�`V� c�V��t\��LmPo�ve4��-�sVP�R�\|�tPV�Qe5.W`V6�*u"��P�}�o`���`��CVKd��N�IIP��CV����IPN9�Gene���D��D�R�D������  ��f谔�p�os.��inal"��n��DeR���`2��d�P��omB���on,���R�D�R��\��TXf��D$b��womp�� "N��dP��m���! ���=C-f����=F�XU�����g Fx��(��Dt II��hr�D��u�� "�<���Cx_ui X������f2��h	�Crl2��D,r9u�i�Ԣ� it2�c�0co��e"�����ا(.)�� ���� ���� IQnQ� �I[ ��{_= wo��,�bD� ��|�GG� ��݅��4 �{e� vʷ� &� 2���Z uz����{�� ��TW&wq~q 5�׷&��o? ;0��  �2� �w�y� ���W&���� ?�3�� A��e��/> �\�3&T���� 77߸� ���� ����� ֵ��&���8 �l1���S�) ����d *J� F�'s ~���� 6:0� ��,���s�- Q�{v� ��� �,�T �ZB�Lx6���6 ���6���ParD ��s>�E��j�6wdsq��F  ��p�����ЁDhel������ti-S`�� �Ob��Dbcf��O�����t OFT��P<A�_�V�Z I��D��V\�qWS��= dtle�Ea�n�(bzd��tiStv�Z�z�Ez :XWO H6�6����5 H�6H69�1�E4܀Tofkst�F� Y682�4܌`�f804�E91�g�`30oBkmon�_�E��eݱ�� q�lm��0 J�fh���B�_  ZDTrfL0�f(P7�EcklKV� �6|��D�85��ّ�m\b�����xo�k�ktq��g2.g���yL�bkLVts��IF��bk������IdG I/f��GR� �han�L��V0y��%��%ere���v��io�� ac�- A�n�h����cuACl�_�^i!r��)�g��	.�@�&� G��R630 ���p v�p�&H�f�f�un��R57v�OJavG�`Y��wowc��-ASF���O��7���SM`�����
af���rafLa�v(l�\F c�w a����?VXpoV �30��NwT "L�FFM���=����yh	a�G-�w:�� �m2.�,�xt��̹�6ԯ6��sd_�MC'V��➟D���fslm��isc.  H5522���21&dc.p�R78����0��708J6�14Vip �ATUu�@�OL�5�45ҴINTL�6��t8 (VC�A���sse�CRI��ȑ��UI����rt\rL�28�g��NRE��.f�,�63!��,�SC�H�d Ek�DOCV���p��C,�<�L��0Q�isp��EI1O��xE,�54��z��9��2\sl,��SET���lр�l�t2�J7�Ռ�MASK��̀�PRXY҇��7����OCO��J6�l�3�l�� (SVl�A�H�L�@Օ��7539Rsv���;#1��LCH����OPLGf�out�l�0��D��HCR.
svg��S@�hƌ�CSa�!�{�50���D�l�5!�lQ��DSW��S����̀���OP����7��PR����L�ұ�(Sg9d���PCM���[R0 \s��5PՄ����0���n�q� EAJ�1��N�q�2��gPRSa���69��� (AuFR�D�Խ��RMCN̪��93A�ɐC_SNBA�F9� 'HLB��� M��h4���h�2A�95z��HTCaԈ�TMI�L6�j95,��8�57.,PA1�i{to��TPTXҴ; JK�TEL��pIiL�� XpL�80ՃI)��.�!��P;�J{95��s "N�ܱ�H�UEC��7\cs�FR��<Q���C��57\{VC�Oa�,���IP1j�H��SUI�	CS�X1�AWEB�a��HTTa�8�RK62��m`��GP%v�IG %tutK�IPGSj�| RC�1_me�H76t��7P�ws_+��?x�R51�\iaw�N���H�53!���wL�8!�h�R66��H���Ԡ����@;J56��1���(N0��9�j��L��ӣR5`%�A|�5q�r��`,�8 5��{165�!��@�"5��H84�!�29��0��PJ����n B[�J77!Ԩ�R6�5h3n�d��y36P��3R6��-`;о Ԩ@��e;xeKJ87��#wJ90!�stu+��~@!䬵�k90�kop�B����@"!�p�@|BA�g*�n@!��Q��06!�@[�F�FaP�6��́,лTS� NC[�CKAB$iͰl1I���R7��@q�y�C�MS1�rog+QM��� �� TY$x�C;TOa�nv\+���1�(�,�6�con��~0��15��JN�N�%e:��P��9O�RS%x���8A�8�15[�FCBaUn�ZQ�P!��p{��CM�OB��"G��OL܀�x�OPI�$\lEr[�SŠ�T	D7�U޹�CPRQR9RL���S�V�~`���K�ETS�$1��0����3�Ԩ�FVR:1�LZQV3D$ ���BVa�SAPLn1�CLN[�PV���	rCCGaԙ��C�L�3CCRA�n� "W!B�H�CSKQn\0�p��,)�0CTPn�ЌQpe��p!$bCt�aqT0U�pCTC�tyЋRC1�1 (�s���trl,�r��
�TX��TCaerr9m�r�MC"�s���#CTE��nrr�REa�XPj�^��Grmc�^�a"�PQF!$���$p e"�rG1�tTG$�c8��QH�$SCT�I�! s��CTLqdACK�Rp)���rLa�R82��M`��YPk�.���OF��.���e�{�CN���^�1�"M�^�a�С@�Q`US��!$��M�QuW�$m�VGF�$oR MH��P2�� H5� ΐq��ΐn�$(MH[�VP�uAoY����$)��D���hg��VPF��"�MHG̑`e!�+�V/vpcm�N��ՙ�8N��$�VPRqd)�&�CV�x�V� "�X�,�1�($TIa�t�\mh��K��et!pK�A%Y�VP%ɠ�!PN���Gen=eB�rip���x�8��extt���Y�m�"�(� �HB���)��x�������Ȣ�r�es.�yA�ɠn@����*���p�@xM�_�NĀ6L�p��Ș�yAvL�0Xr�Ȉ2��"R;�Ƚ�\ra��	P�� h86��Gu+ʸ�φ��SeLɨm�9�69�P�Ȩr�Ȩ2�ɹ1&��n2�h� �0L�,XR}�RI{�e� L�x���c�Ș���N��vx�L��"��2\r@�]�N�82�d����b�ɉa��y1��/�kp�@���A��ruk��� L�sop��H�}�Cts{�����s�ʼ9��j965��S�c��h��5 J9��{�
�PL�J	e;en��t I[
x��com��Fh�L�4c J��fo��DIF+�6�Q���ڏrati|��p��1L�0�
R8l߾�M�����P��8� �j�mK�X�HZ�����N�oڠ��3̹q��vi���80�~�l Sl�yQ�F�tpk�xb�j� .�@�R�d������,/n(�8�8�0���
�:�O8�<�Q}�COt���PT��O (��.�Xp|�~H���?�ov �wv���8�22�pm���722��j7�^�@�̙���cf�=Yvr���vcu���O��O�O�O_#_5_7�3�Y_��wv4{_�_yw�ʈ�ust_�_�cus�_�Z��o�o,o>oPo�io��n�ge��(pLy747��jWelʨHM47ZKEq {���[�m�MFH�?�(ws K�8J�n���oΝ�fhl;��wm�f���? :�}(4�	<g J{��II�)̏މw��X�7714kﭏ/7ntˏ݊�e+���se�/�a!w��8�ɐ��EX \��!+: �p��~�002��nh�,:Mo+�xO���1 "K�O��\a��#0��.8���{�h�L?�j+�mond�:��t�/�st�?-�w�:���)�;��p(=h�;
d Pۻ��{:  ���� �J0��re�����STD�!t�reLANG����81�\tqd��������rch�.������ht�wv�WWָ� wR79��"Lo�51 (�I�W�h�8Ո�4�aww�� �vy �623�c�h a?�cti �֘!�X�iؠ�	t ��n,�։�����j��"AJ1P@�3p�vr{�H��6��!��- Se�T� E3�) G�J9�34��LoW�4 (S������ <����91 ��8!4�j9 �所+���y�
��	�btN�ite{�R  ��I@Ո�����P� ������	 ����Z�vol��X ��9�<�I�p���ld*���F�864{��?��K�	�k扐�֘1�/wmsk��M�q�Xa�e����rp��0RBT�1�ks.OPT�N�qf�U$ RTCamT��y��U ��y��U��UlU6L�T�1Tx����"SFq�Ue�6T���USP W�b DT�qT2h�T�!�/&+��TX�U\j6&�U U�UsfdO&�&ȁT����662DPN�bi��%�Q�%62V��$���%�� ��#(�(6To6e #St�%��#5y�$\�)5(To�%tT0�%5�W6T���%�#�#orc��#I���#���%cct�6ؑ?��4\W6965"8p6}"�#\j536�p��4�"�?kruO O,Im?Np�C �?�t�0<O�;�e ��%���?
;gcJ7 �"AV�?�;avs�f�O__&_8Wtp�D_V_0GT�F|_:Uc�K6�_�_r�O�3e\�s�O2^y`O:�miugxGvgW! m�%��!�%T�$E A`{6�po6��#37N��)5R5_2E���$0\���$Ada�Vd�Ѐ�V�?;Tz7�_�e7DCDTF9���#8�`��%��4y�te�d Z@�A}�@�}�0�4N�}�}���}�d�c& }����u 6��v��v1�u1\b��u$2}���}� R8�3�u�"}��"}�vaClg���Nrh�&�8�J�Y�o�ue���� j70�v=1��M{IG�uerfa��{q���E�N�ء���EYE�ce A ���񁏯pV�e�A!�� �2Յ�Q�%��u1�e�i�@��H�e����J0�� '��b��T��E In�B�  W�|��537g�����(MI�t�Ԇr��ݟ�am���n�ҵv!g�U -�v J�߆8⹖F���P�y�a�c���2���Rɏ j�o��2�� djdx�8r}� og\k��0��g��wmf��Fro/� Eqx'�4"}�3 J8��oni[��ᅩ}Ĵ�� o� ��ʛ���m@�R�e��{n�Д�V�o�������  �������"POS\����ͯ menϖ�⑥OMo�43��� �w(Coc� An[�0t���"e�a\�vp�z��.��cflx$�le��8�hr�trᅻNT� CF+�x E/�t	qi�M�ӓcxc��p�f�lx��,��Z�cx��
0 h�6��h8��mo��=�c H���)� (�vSER,���g�0߆0\r�vX�= ���I � - �tiغ�H��VC�82�8�5��L"�RC���n G/���w�P��y�\v�vm " o�lϚ�x`��=e�ߠ-�R-3?�����x�vM [�AX/2�\)�S�rxl�v#�0氆h8߷=� RA�X�A�����9�H��E/Rצ����hN߶"RXk��F�v˦85��2L/�xNB885_�q�Ro��0iA��5\r�O�9�K��v����88���.�n "�v��88��8s�i ?�9  ��/�$�y O��MS"���&�9R� H74&�`�74�5�	p��p��yc�r0C�c�hP0� �j�-�a%?o��6D95�0R7trl��c;tlO�APC����j�ui"�L���  ]����^棆!�A���qH��&-^7�w��� ���616C�q�794h���� M�ƔI���99��(���$FEAT_A�DD ?	����Q%P  	�H._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����������& 8J\n���������TDE�MO fY   WM_ �������� //%/R/I/[/�// �/�/�/�/�/�/�/? !?N?E?W?�?{?�?�? �?�?�?�?�?OOJO AOSO�OwO�O�O�O�O �O�O�O__F_=_O_ |_s_�_�_�_�_�_�_ �_ooBo9oKoxooo �o�o�o�o�o�o�o >5Gtk}� �������:� 1�C�p�g�y������� ܏ӏ���	�6�-�?� l�c�u�������؟ϟ ����2�)�;�h�_� q�������ԯ˯ݯ�� �.�%�7�d�[�m��� ����пǿٿ���*� !�3�`�W�iϖύϟ� ����������&��/� \�S�eߒ߉ߛ��߿� ������"��+�X�O� a����������� ����'�T�K�]��� �������������� #PGY�}� ����� LCU�y��� ���/	//H/?/ Q/~/u/�/�/�/�/�/ �/???D?;?M?z? q?�?�?�?�?�?�?
O OO@O7OIOvOmOO �O�O�O�O�O_�O_ <_3_E_r_i_{_�_�_ �_�_�_o�_o8o/o Aonoeowo�o�o�o�o �o�o�o4+=j as������ ��0�'�9�f�]�o� ��������ɏ����� ,�#�5�b�Y�k����� ����ş����(�� 1�^�U�g��������� ������$��-�Z� Q�c������������ �� ��)�V�M�_� �σϕϯϹ������� ��%�R�I�[߈�� �߫ߵ��������� !�N�E�W��{��� �����������J� A�S���w��������� ����F=O |s������ B9Kxo ������/� />/5/G/t/k/}/�/ �/�/�/�/?�/?:? 1?C?p?g?y?�?�?�? �?�? O�?	O6O-O?O lOcOuO�O�O�O�O�O �O�O_2_)_;_h___ q_�_�_�_�_�_�_�_ o.o%o7odo[omo�o �o�o�o�o�o�o�o* !3`Wi��� �����&��/� \�S�e���������� ����"��+�X�O� a�{����������ߟ ���'�T�K�]�w� ���������ۯ�� �#�P�G�Y�s�}��� �����׿���� L�C�U�o�yϦϝϯ� �������	��H�?� Q�k�uߢߙ߫����� �����D�;�M�g� q����������
� ��@�7�I�c�m��� ������������ <3E_i��� ����8/ A[e����� ���/4/+/=/W/ a/�/�/�/�/�/�/�/ �/?0?'?9?S?]?�? �?�?�?�?�?�?�?�? ,O#O5OOOYO�O}O�O �O�O�O�O�O�O(__ 1_K_U_�_y_�_�_�_ �_�_�_�_$oo-oGo Qo~ouo�o�o�o�o�o �o�o )CMz q������� ��%�?�I�v�m�� �������ُ���>;�  2�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s��������'9  :>Ugy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������/=C6Yk }������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ������/�A��$FEA�T_DEMOIN�  E��q���>�Y�INDEX�f�u��Y�ILE�COMP gw�����t��T���SETUP2� h������  N ܑ��_�AP2BCK 1�i��  �)�B���%�C�>� ��1�n�E����)��� M�˯�������<�N� ݯr������7�̿[� �ϑ�&ϵ�J�ٿW� ��Ϥ�3�����i��� ��"�4���X���|ߎ� ߲�A���e����� 0��T�f��ߊ��� ��O���s�����>� ��b���o���'���K� ��������:L�� p����5�Y� }�$�H�l~ �1��g��  /2/�V/�z/	/�/ �/?/�/c/�/
?�/.? �/R?d?�/�??�?�? M?�?q?O�?O<O����P� 2��*.VRCO�O�0*�O�O�3�O�O�5w@�PC�O_�0FR6:�O=^�Oa_�KT���_�_&U�_�\h�xR_�_�6*.FzODo�1	(SoEl�_<io�[STM �b�oН^+P�o�m�0i�Pendant �Panel�o�[H �o �g�oYor�ZGIF|��e�O8a��ZJPG �*���e���z��JJS������0@���X�%�
JavaScrgiptُ�CSʏ�1��f�ۏ %C�ascading� Style S�heets]��0
�ARGNAME.SDT���<�`\���^���Д៍�АDISP*ן���`$��d��V�e��CLLB.ZI��=�/`K:\��\�����Collabo����	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V���zό�!ߘ�TPEINS.XML(��@�:\<����Cu�stom Too�lbar}��PA?SSWORD���>?FRS:\���� %Passw�ord Config��?J���C�� "O��3�����i���� "�4���X���|��� ��A���e�����0 ��Tf����� O�s��>� b�[�'�K� ��/�:/L/�p/ ��/#/5/�/Y/�/}/ �/$?�/H?�/l?~?? �?1?�?�?g?�?�? O �?�?VO�?zO	OsO�O ?O�OcO�O
_�O._�O R_d_�O�__�_;_M_ �_q_o�_�_<o�_`o �_�o�o%o�oIo�o�o o�o8�o�on�o �!��W�{� "��F��j�|���� /�ďS�e�������� �T��x������=� ҟa������,���P� ߟ񟆯���9���� o����(�:�ɯ^�� ����#���G�ܿk�}� ϡ�6�ſ/�l����� ϴ���U���y�� � ��D���h���	ߞ�-߀��Q߻��߇��,���$FILE_DG�BCK 1i������� ( �)
S�UMMARY.DyG,���MD:`������Diag� Summary����
CONSLOG��y����$����Console� log%���	T�PACCN��%�g�����TP A�ccountin�F���FR6:I�PKDMP.ZI	P����
��)�����Exceptio�n-����MEMCHECK������8�Memory� Data��L�N�)�RIP�E���0�%�� Packe�t LE���$S<n�STAT*|#� %L?Status�i	FTP�/�/��:�mment� TBD=/� >�)ETHERNE�/o�/�/��EthernU~<�figuraL���'!DCSVRF�1//)/B?�0 �verify a�llE?�M(5DIFF:? ?2?x�?F\8diff�?�}7o0CHGD1p�?�?�?LO �?,sO~3&�
I2BO)O;O�O bO�O�O�GD3�O�O�OT_� �O{_
VUP?DATES.�P�_~��FRS:\�_��]��Updates List�_���PSRBWLD'.CMo���Ro��_9�PS_ROB�OWEL^/�/:G�IG��o>_�o��GigE ��no�sticW�N��>�)�aHAD�OW�o�o�ob��Shadow C�hange���8+"rNOTI�?=O��Notific�"���O�A�PMIO�o��h��f/��on�^U�*�UI3�0E�W��{�UI������B���f��_��� ����O��������� >�P�ߟt������9� ί]�򯁯�(���L� ۯp������5�ʿܿ k� Ϗ�$�6�ſZ�� ~��wϴ�C���g��� ߝ�2���V�h��ό� ߰���Q���u�
�� �@���d��߈��)� ��M���������<� N���r����%����� [����&��J�� n��3��i ��"�X�| ��A�e�/ �0/�T/f/��//�/=/�/�/�$�$FoILE_�PPR�P���� �����(MDO?NLY 1i5� ? 
 �z/Q? �/u?�/�?�?t/�?^? �?O�?)O�?MO_O�? �OO�O�OHO�OlO_ �O_7_�O[_�O_�_  _�_D_�_�_z_o�_ 3oEo�_io�_�oo�o �oRo�ovo�oA �oew�*�� `����&�O��*?VISBCK,81>;3*.VDV�����FR:\o�I�ON\DATA\�/��Vis�ion VD filȅ��&�<� J�4�n������3�ȟ W������"���F�՟ �|������m�֯e� �����0���T��x� �����=�ҿa�s�� ��,�>���b���� �ϼ�K���o��ߥπ:���^����ϔ��*M�R2_GRP 1�j;�C4 w B�}�	 71�������E�� E��  F@ F��5U������L����M��J�k�Lzp�JP��Fg�f�?�  S����9��Y9}�9���8j
�6��6�;���A�  ���BH���B���B���$�������������@UUU#����� Y�D�}�h����������������
C��_�CFG k;T M���]��NO :
�F0� � \�RM�_CHKTYP  0�}�000���OM_MI9N	x���50�X� SSBdl.5:0��b�x�Y���%TP_?DEF_OW0x��9�IRCOM���$GENO�VRD_DO*�62�THR* dz%d�_ENB�{ �RAVC��9mK�� ��՚�/3�/��/�/�� �M!OUW s��}��ؾ��8�g�;?�/7?�Y?[?  C��0�a���(7�?�<B�?B����2��*9�N SMTT#t[)��X��4�$HOSTC�d1ux��֮? 	zHzKdzOx��O�Ie�O �O	__-_;Z�O^_p_��_�_�O�_KP	anonymous�_ �_�_oo1o yO�O �Ozo�_�OM_�o�o�o �o?_.@Rd�o �_�_�����;o Mo_oqos`��o���� ����̏����&� 8�[����������� ȟ�!�3��G�4�{� X�j�|���Տ��į֯ �����e�B�T�f� x���џ����	�� =��,�>�P�bϩ��� �Ϫϼ����'�9�� (�:�L�^ߥ���ɿw� ������� ��$�6� ��Z�l�~��ߴ��� ������� �g�yߋ� ��z����߰������� ��?�.@Rd�� ��������;� M�_�q�s`���� ����//&/ I7/�n/�/�/�/�/�#O\AENT 1v�
; P!J/?  ��/3?"?W? ?{?>?�?b?�?�?�? �?�?O�?AOOeO(O �OLO^O�O�O�O�O_ �O+_�O _a_$_�_H_ �_l_�_�_�_o�_'o �_Koooo2o{oVo�o �o�o�o�o�o5�o Y.�R�v���zQUICC0 ���3��t14��"����t2��`�r�ӏ�!ROUTER�ԏ��#�!PC�JOG$���!�192.168.�0.10��sCA�MPRTt�P�!bd�1m�����RT�🟱���$NAME� !�*!RO�BO���S_CF�G 1u�) ��Auto�-started^FTP&�� =?/֯s����0� B��f�x��������� S������,���� �����ϼ�ޯ������ ���ʿ'�9�K�]�o� ��ߥ߷��������� (:~�k�Ϗ� ������������ 1�C�f���y������� �����,�>�R�? ��cu��`��� ��(�$M_ q������  /H%/7/I/[/m/4 �/�/�/�/�/�~/? !?3?E?W?i?��� �?�/�?/�?OO/O �/�?eOwO�O�O�?�O RO�O�O__+_r?�? �?�?�O|_�?�_�_�_ �_o�O'o9oKo]ooo �_o�o�o�o�o�o�o F_X_j_~ok�_� �����o��� 1�TU��y����������U�)�_ERR �w3�я�PDU�SIZ  g�^ڀp���>�WR�D ?r�Cq� � guestb�Q�c�u��������"�SCDMNG�RP 2xr����Cqg�\��b�K� 	P0�1.00 8(q _  �5p�5p�z�5pB  ��{ ���H����L��L��>L�����O8������l�����a4� �x��Ȥ�x��8��U�\���)�`蠍;�������d��.�@�R�ɛ_GR�OUېy���⽒	ӑ���QUPOD  ?u����VİTYg�����TTP_AUTH� 1z�� <!�iPendan䷗-�l���!KAREL:*-�6�H�KC]�m���U�VISION SET���ϴ�g� G�U������R�0�� H�Bߏ�f�x��ߜ߮����CTRL {�����g�
S�?FFF9E3��At�FRS:DEF�AULT;�F�ANUC Web Server;� )����9�K��ܭ����������߄WR_�CONFIG �|ߛ ;��I�DL_CPU_P5CZ�g�B�Dpy�w BH_�MINj��)�}�GNR_IO���g���a�NPT?_SIM_D_������STAL_S�CRN�� ���T�PMODNTOL8������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMAST�E��ɾeSLAV�E ~��c�O�_CFGٱBU�O�O@CYCL�En>T�_ASG� 1ߗ+�
  ����//+/=/ O/a/s/�/�/�/�/���NUM��
�@IPCH�^R?TRY_CNZ��@�@��������1 @kI�+E��z?E�a�P_MEMBERS 2�ߙ�� $���2����ݰ7�?�9a�SDT�_ISOLC  �����$J23�_DSM+�3J?OBPROCN���JOG��1�+��d8�?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSRE�QO��KANJI_����a[�MONG ����b�yN_ goyo�o�o�o�Y�`3	�<� ��e�_ִ���_L���"?`EY�LOGGINL�E�������$L�ANGUAGE Y��<T� {q��LGa2�	�b����g�xP��  *��g�'��b����>�MC:�\RSCH\00�\<�XpN_DISP �+G�J��O��O߃LOCp�D�z���AsOGB?OOK ����`��󑧱����X� ����Ϗ����a�*��	p������!�m��!���=p_B�UFF 1�p��2F幟���՟�D� Collaborativǖ ���F�=�O�a�s��� ����֯ͯ߯����B�9�K���DCS ��z� =��� '�f��?ɿۿ���H@�{�IO 1��# ~?9ü��9�I� [�mρϑϣϵ����� �����!�3�E�Y�i� {ߍߡ߱��������-E��TMNd�_B� T�f�x�������� ������,�>�P�b��t�������L��SE�VD0��TYPN1�$6���Q�RS"0&��<2FLg 1�"�J0��� �����G�TP:pOF�NGNAM1D�mr�t7UPS�GI"5�a�O5�_LOAD�N@G %�%�TG1#$$MA?XUALRM�'��8�(��_PR"4F0�d��1�B_PN�P� V 2�C�	MDR077���BL"806=3%�@ �_#?�hߒ|/�C��z��6��/���/Po@P �2��+ �ɖ	��	t  ��/�%W?B?{?� k?�?g?�?�?�?O�? *OONO`OCO�OoO�O �O�O�O�O_�O&_8_ _\_G_�_�_u_�_�_ �_�_�_o�_4ooXo joMo�oyo�o�o�o�o �o�o0B%fQ �u������ ��>�)�b�M����� {��������Տ�� :�%�^�p�S��������D_LDXDI�SApB�MEM�O_APjE ?=C
 �,� (�:�L�^�p�������ISC 1�C ����4�����૟4��X���C_M?STR ���w��SCD 1��� L�ƿH��տ���2� �/�h�Sό�wϰϛ� �Ͽ���
���.��R� =�v�aߚ߅ߗ��߻� ������<�'�L�r� ]���������� ����8�#�\�G���k� ��������������" F1jUg�� �����B -fQ�u����h�MKCFG 񓆽�/�#LTAR�M_��7"�0�0N/V$� MEgTPUᐒ3�����ND� ADCOLxp%� {.CMNT�/s �%� �����.E#>!�/4�%PO�SCF�'�.PR�PM�/9ST� 1���� 4@��<#�
1�5�?�7 {?�?�?�?�?�?�?)O OO_OAOSO�OwO�O��O�O�O_�A�!SI�NG_CHK  ��/$MODAQ�,#����.;UDE�V 	��	M�C:o\HSIZE�ᝢ��;UTASK� %��%$12�3456789 ��_�U9WTRIG +1���l3%%��9o���"ocoFo5#�VYP�QNe��:SEM_�INF 1�3'� `)�AT&FV0E0�po�m)�aE0V�1&A3&B1&�D2&S0&C1�S0=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o '��K������ ��я:�L�3�p�#� 5���Y�k�}������ $�[�H���~�9��� ��Ưد��������ӟ �V�	�z�������c� Կ����
��.��� d��)�;��Ͼ�q��� ����˿<���`�G� �ߖ�IϺ�m�ϑϣ� ���8�J��n�!ߒ��M�������h_NIwTOR� G ?�[�   	EX�EC1�/�25�3�5�45�55��P7�7*5�85�9�0�� ��4��@��L��X� ��d��p��|�������2��2��2���2��2��2��2���2��223ʡ�3��3@�;QR_�GRP_SV 1ݚ�k (�5W�r>���������MO�Q_�D��^�PL_N�AME !3%�,�!Defa�ult Pers�onality �(from FD�) �RR2� �1�L6(L�?�,0	l d �������� //(/:/L/^/p/�/��/�/�/�/�/�/ZX2 u?0?B?T?f?x?�?�?�?�?\R<?�?�? O O2ODOVOhOzO�O��O�OZZ`\RD�?�N
�O_\TP�O :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo _)_~o�o�o�o�o�o �o�o 2DVh z�[omo���� 
��.�@�R�d�v����������Џ� �Ef  Fb� gF7�����!��d�?�Q�6� t���������ʜ8����� ݘ� ���"�@�F�d���� �"𩯹�� A� � ϩU[�$n��B�E ��� � @D��  �?�� �?x�@��A@�;f�|�FH� ;�	l,��	 |��j��s�d�>��� ���� K(��Kd�$2K ��J7�w�KYJ���ϜJ�	�ܿ��� @I���_f��@�z��f��γ�N�������	Xl�������S�Ľ�Ô��X������5���  �����A?oi#��;���� � �l� �Ϫ�-���ܛ�G�G����@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=������@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj�a�Be�Ci��@#��Bи�M L� 2���~��bbdʷBР��P����̠�����ADz՟�n�3� �C�i�@�R�R�Yщ���  �@� ����  ��?��ff������n�  ɠ#�y9G
(�$��I�(�@uP~�����t�t���>����;��Cd;��.<�߈<�g�<F+<L��������,�d�,�̠?f7ff?��?&&���@��@x���@�N�@���@T�H�ِ�! -�ȹ�|��
`� ������//</�'/`/r/]/�/��eF���/�/�/�/m?Б�/J?�(E��G=�#�� FY�T? �?P?�?�?�?�?�?O �?/OO?OeO�ħO �IQOG�?�O1?�OmO _0_B_T_������A_�_	_�_�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�o�o����W�����oC�E� q�H�d���؜a@q��e�F�B�µWB]�NB�2�(A��@�u\?�D��������b�0�|��uR����
�x~�ؽ���Bu*C��$��)`�$ ����GC#������rAU����1�eG�D��I�mH�� �I:�I�6[�F���C�I���J�:\I�T�H
~QF�y��p�*�J�/ I8Y��I��KFjʻCe�o��s�����Џ ���ߏ�*��N�9� r�]������������ ۟���8�#�\�G��� ��}�����گů��� "���X�C�|�g��� ��Ŀ�������	� B�-�f�Qϊ�uχ��� ���������,��P� b�M߆�qߪߕ��߹� ������(��L�7�p� [���������s=(la��3:��s��$�le3���d8�,�4��@�R�wa����l�~�wa����e����wa4 �{������(PL:ueP�P~�A�O�����<�	���� G2W}h��� ���/���O�O7/m/[(d=�s/U/�/ �/�/�/�/?�/1??�U?C?y?�=  2 wEf9gFb��7�7�9fB)aa)`C%9A`�&`w`@-o�?�9de�O-OOQOpn��?�?�O�O�O�O9c?��0�A7hldw`�w`!w`xn
 �O9_K_]_o_�_�_ �_�_�_�_�_�_o#o�zzQ ��h��G����$MR_CABLE 2�h� �a�T� @@�0�Ae��a,�a�a��`��0�`�C�`�aO8�tB��n��ECG+���F�o�f�#���0��0�DO���By`,�0/��EAA�V���o�h�8  ��a�07�d4
v3���v�O�"4�Ƞ`y`
qC�p�bHE��
v�y�mҠ`�p�0�q�p�b0��`�����#�5C�0��y��c-��� H� �2���V������� ����'�"���D������o��\����������������*,�** \cOM� �ii������cr�%% 2�34567890	1i�{� f�����������1�����
��`�not? sent 5����;�TES�TFECSALG�R  eg`��1d�.�š
:�� ��DCbS�Q�c�u��� �9UD1:\m�aintenances.xml���ֿ  Z�DEFAULT-��i4\bGRP 2��M�  =��7�E � �%Forc�e�sor ch�eck  �����Bz��p����h5-���ϻ��������%!�1st clea�ning of cont. v�ilation��}�Rߗ+��[�ߔ��߸���mec�h�cal`�������0��h5 k�@�R�d�v����(�rolle_Ƶ����/���(�:��L��Basic� quarterCly�������,������������MH��:(�"GpP(�X_h5�������#C���M"��{Pbt����Suppq�grease���?/&/8/J/\/���C+ ge��. batn�y`/��/h5	/�/�/�/? ?X_�ѷen'�v��/�/��/��?�?�?�?�?�G=?O(��Dp"CrB1O��0 �/`OrO�O�O�O�t$,��Lf��C-(��A�O:�OO$_6_H_Z_�l_�t*cabl,�O(���S<(��Q�_:�
_�_�_oo�0oo)(Ӂ/�_�_����_�o�o�o�o�o��O@hau1�l�2r x(�<qC:��op������_ReplaW�fU��2�:�._4�F�X�j�|�(�$%���ߟ ����#���
��.�@� ��d���ŏ׏����П ����U�*�y����� r���������	�q�� ?�߯c�8�J�\�n��� ϯ�����ڿ)���� "�4�Fϕ�jϹ�˿�� ����������[�0� ϑ�fߵϊߜ߮��� ��!���E�W�,�{�P� b�t����߼��� ��A��(�:�L�^��� ������������  $s�H������q �����9] o�Vhz��� U�#�G/./@/ R/d/��/�/��// �/�/??*?y/N?�/ �/�?�/�?�?�?�?�? ??Oc?u?JO�?nO�O��O�O�O+Jkb	 H �O�O__6M2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o�*<ND@ ̾bA?�  @!Q _���Fwp�� �H* �** @A>F�pRT��f�x�:�������ҏ��eO^C7�Տ#�5� G�	�k�}���ُ��� c�����W��C�U� g���ß)�����ӯ� ��	��-�w�����9� ������m�Ͽ��=��O�E!Q�$MR�_HIST 2��>EN�� 
 \�
B$ 2345678901^�f�#�
�]�9O���φ� ��O�)�;����q� �ߕ�L�^߬����ߦ� ���7�I� �m�$�� ��Z���~������!� ��E�W��{�2������h�����:�SKCF�MAP  >EKQ��r5�!P�����ONREL7  .�3����EXCFENB�8
��QFNC�XJJOGOVL�IM8dNá ��K�EY8��_�PAN7����R�UN����SFSPDTYPx<C��SIGN8J�T1MOT�G���_CE_GRP7 1�>EV� �@�����/Ⱥ ��/�/U//y/ 0/n/�/f/�/�/�/	? �/???�/c??\?�? P?�?�?�?�?�?O)O�OMO,���QZ_E�DIT5 )TC�OM_CFG 1����[�O�O�O }
�ASI �yB3�
__+[_�O_��>O�_bHT__ARC_U.���	T_MN_MO�DE5�	UA�P_CPL�_gN�OCHECK ?��� ��  o.o@oRodovo�o�o �o�o�o�o�o*�!NO_WAITc_L4~GiNT�A����EUwT_E�RRs2���3��@ƱJ�����>_�)��|MO�s��}x�:I8@�oA�M�˞´4�8�?����� �~��rPARAM�r�.����r_�p:H5�5�G� = �� d�v�~�X�������������֟�0��:G��b�t�����SUM_RSPACE������Aѯۤ�$OD�RDSP�S7cO�FFSET_CAqRt@�_�DIS���PEN_FIL�E:�7�AF�PT?ION_IO���q�M_PRG %��%$*����M�WORK �y=f ��춍�@�� �E����	 ���Í��It��RG_DSBL  ���C�{u��RIE�NTTO7 �C�~�A �UT__SIM_Dy����V�LCT ���}{B �٭��_�PEX�P=��RA-T�W dc���UP ���`����e�w�]ߛߩ���$�2r�L6�(L?���	l d������&� 8�J�\�n����� ���������"�4�F�X���2�߈��������������*�< w�Tfx��������J` �DT��Tz��Pg������ /"/4/F/X/j/|/�/ �/�/���/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?�/�/,O>O PObOtO�O�O�O�O�O �O�O__(_:_��O�Z��y_�]2ӆ� �_�^�_�_�W^]^]��/ooSog��Hgro hozo�o�o�o�o�oF`��#|`�A� � 9y����OK�1��k������<�E�A�nq @D�C  �q����nq?���C��s�q1� ;��	l��	 �|�Q�s�r�q>���u �sF`H<�zH~�H3�k7GL�zH?pG�99l7�0k_B�T�F`C4��k��H���t��-�Z�����k�����~s���  �ሏ�����EeBVT����dZ�����ڏ ���q�-�Fk�y�{FbU����n@6�  ���z�Fo���[�	'� � ���I� � � �:p܋=��q�ڟ웆�@�@��B�,���B����g�
�N����  '�|���g��B��
p�BӀC׏����@?  #�Bu�&����� �_bbd�B:p 2���>�m�6p�Z���Dz?o}�܏�������׿������Ǒ��� ~f�  � �M�z��*�?�ff�_8�J�ܿ 3pϑ�ñ8= �ϵʖq.·�	(= ��P���'��s��tL�>��/�;�C�d;��.<���<�g�<F+<L ��^oiΚr�d@��r6p?fff�?�?&���@���@x��@��N�@���@T싶�Z���ћtމ �u�߈w	�x��ti�>� )�b�M��q����� ��������:�%�^��������W���S�E��  G�=F�� Fk��������� 1U@yd�� ����q��	�� {�A��h����D�a��ird��A{�/w/J/5/n/vA�A���":t�/ C�^/�/Z/ ލ?����/�/1??���Wҵ���g��pE�! ~1�?04�0
1ή1@IӀ��B���WB]�NB2��(A��@��u\?��������������b�0�|�uR����
�>��ؽ��B�u*C��$��)`�? ����GC#����rAU�����1�eG���I��mH�� I�:�I�6[Fߍ��C4OI���J�:\IT��H
~QF��y�Ol@�*J��/ I8Y�I���KFjʻC ��-?�O�O__>_)_ b_M_�_�_�_�_�_�_ �_o�_(oo%o^oIo �omo�o�o�o�o�o  �o$H3lW� {������� 2��V�h�S���w��� ��ԏ�������.�� R�=�v�a�������П ����ߟ��<�'�`� K�]���������ޯɯ���&�8�#�\��3(�J���3:a���9���J�3��c4�����������������ڿ�n�����e��n�4 �{2�2�r�`ϖτ�(�Ϩ��%PR�P���!�h�!�K�6�o�Z�����u�|ߵ� �����������3�� W�B�{�f�4���������d�A����!�� 1�3�E�{�i��������������  2 �Ef�7Fb�7���6B�!�!� C9� �� n�@�/`r@������#x�@�+=�3?, TV�8v�n�n���n��.
  D�����// %/7/I/[/m//�/�:� ��ֻ�G����$PARAM�_MENU ?�2�� � DEFP�ULSE�+	W�AITTMOUT��+RCV? �SHELL_W�RK.$CUR_oSTYL� 4<�OPTJJ?PTB�_?Y2C/?R_DECSN 0�Ű<�?�? �?�?�?OO?O:OLO�^O�O�O�O�O�O�!S�SREL_ID � .����EUS�E_PROG �%�*%�O0_�CCC�R0�B��#CW_H�OST !�*!HT�_=ZT��O_�S�h_zQ�S�_<[_TGIME
2�FXU� ?GDEBUG�@�+��CGINP_FLgMSKo5iTRDo�5gPGAb` %l��tkCHCo4hTY+PE�,� �O�O �o#0Bkfx �������� �C�>�P�b������� ��ӏΏ�����(��:�c�^�p�����7eW�ORD ?	�+
? 	RSc`n�/PNS��C4�sJOv1��TE�P�COL�է�2�Z�gLP 3��n���OjTRACEC�TL 1�2���! �� �Қ�q�DT� Q�2�Ǡ���D � ���:�� ܠ�)ԯ�����}��`�,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �Щ*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6Fl~� ������� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�x�N�߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`?�r?�?�?�?�?�9�$�PGTRACEL�EN  �1  ���0���6_UP �/���A@�1�@�1_CFG7 �E�3�1
@�<D�3UOaH�SO�0$BDEFSP/D �/L�1�0���0H_CON?FIG �E�3W �0�0d�DM��2 �1�APpD�sA�A�0��0IN~'@TRL �/M�OA8pEQPE�E��G�A<D�A�ILID(C�/M	~bTGRP 1ýI� l�1B�  �����1A��33FC� F�8� E�� @eN	�A�AsA�Y�Y�A~�@� 	 vO8�Fg�_ ´8cokB;`baBo,o>oxo�bo�o�1>о�?�B/�o�o~�o �=%<�� 
C@yd���"������  Dz@�I�@A0�q�  �������ˏ���ڏ ���7�"�4�m�X����|���Ú)ґ
V�7.10beta�1HF @��=��Aq��Q�  �?� �B�ܠP�p �C���&�B�EQA� ��Q�P�Q�� ß[�m����<CA��0�b �A��̯ޯ��1!CeQ�KNOW_M  �lE7FbTSV ĽJ�BoC_�b� t�������������1��]aSM�SŽK ���	NB�0����ĿK���-�bb��A�R� �P����0�Ŗ��bQ+MR�S��T�iN�`��d���V]ST�Q�1 1�K
 4MU�i��c�kFK�]� oߠߓߥ߷������� 2��#�h�G�Y��}� �������
�������,�27�I��1�<t�H��P3^�p�����,�4��������,�A5(:,�6Wi{�,�7����,�8�!3,�7MAD�6 F,�OVLD  K�D�xO.�PARNUM  �/�_T_SCH� E�
9'!G)�3Y%UP�D/%�E�/P�_C�MP_��0@�0'�7E�$ER_CH�K�%5H�&�/�+RqS���bQ_MO��+?=5_'?O�_RES_G6��:�I�o �?�?�?�?O�?O7O *O[ONOOrO�O�O�{4]��<�?�Oz5�� �O__|3 #_B_G_ |3V b_�_�_|3� �_ �_�_|3� �_�_o|3�Oo>oCo|2V 1��:�k1!�@c?��=2THR_IN�Rc0i!}�o5d�fM�ASS�o Z�gM�N�o�cMON_QUEUE �:ը"�j0��t4N� U�1Nv�+DpEND8Fqd?`yEXEo`uƅ BEnpPAsOP�TIOMwm;DpPR�OGRAM %�$z%Cp}o(/BrT�ASK_I��~O?CFG �$/��K�DATA��&T���j12,ź� ̏ޏ�����&�8�J� \�n��������ȟ{��INFO�͘�� 3t��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����
�Θ� 4�FJ�a K_N��T��˶�ENBg ڽw1��2���GN�2�ڻ� P(O�=�{��]ϸ�@���v� �u�uɡd�Ʒ_EDIT ��T�����G�WER�FL�x�c)�RGA�DJ Ҷ�A�  $�?j00��a��Dqձӆ5'�?��ʨ�<u�j0�%e������FӨ��2�R��	H;plR�G�b_�>�pAodw�t$�*�=/� **:�j0�$�@�5Y�T���^��q�߈b~�L�� \�n��������� ������4�F�t�j� |�������������b LBT�x� ���:��$ ,�Pb���/ ����/~/(/:/ h/^/p/�/�/�/�/�/ �/V? ??@?6?H?�? l?~?�?�?�?.O�?�? OO O�ODOVO�OzO �O_�O�O�O�O�Or_ _._\_R_d_�_�_�_�_�_�_�f	g�io�p Wo�o{d�o�~o�o�zoB�PREF� �Rږp�p
~�IORITY�w�[���MPDSP�q��pwUT6�����ODUCT3������OG��_�TG��8��ʯrTO�ENT 1׶�� (!AF_I�NE�p,�7�!�tcp7�_�!�udN���!iccmv��ޯrXYK��ض���q)� 0,�����p��&� 	��R�9�v�]�o��� ��П������*��$N�`�*�sK��9}�߸����Ư ,�/�6쒯�����خ�A~t�,  �Hp ��P�b�t����u�w��HANCE �R��:�wd��连��2s�9Ks��PO�RT_NUM�s�p���_CARTREP{p�Ω��SKSTA�w nd�LGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_�a_seiban �o\��olߒ�}߶ߡ� ��������"���X� C�|�g�������� �����	�B�-�f�Q� ��u����������� ��,<bM�q �������(�L�VERSI�yp�w} disabledWSAVE ߾z�	2600H7K68S?�!ؿ0����/ 	5(�r$)og+^/y�e{/�/�/�/�/�*�,/?� �p���_�p 1��Ћ� �����Wh?z?�W*p/URGE��B�p}vlgu,�WF�0DO�v�Ʋ�vW%��4(�C�W�RUP_DELA�Y �\κ5R_?HOT %Nf�q�׿GO�5R_NORMAL&H�r6O�OZGSEMIjO�O�O(q_QSKIPF3��W3x=_98_J_\_ ]�_�_{_�_�_�_�_ �_�_	o/oAoSoowo eo�o�o�o�o�o�o�o +=aOq� �������'� �7�]�K�������)Eo�$RA{���K�/�zĀÁ_PAR�AM�A3��K �@.�@`�61�2�C<��y��C��6$�BÀBTI�F�4`�RCVTMkOUu�c��À�DCRF3��I ��+QB
$��D�ZD2Y��1>��78�I]�÷<ޅ���x.�p�]��"-W_��k_ �;�Cd;��.�<߈<�g��<F+<L�� �Ѱ��d�u�L��� ����ϯ����)��;�M�_���RDIO�_TYPE  �M=U�k�EFPOS�1 1�\�
 x4/�����+�$/ <��$υ�pϩ�D��� h��ό��'������ o�
ߓ�.ߤ�Rߌ��� ����5���Y���i� ��*�<�v���r���� �����U�@�y���� 8���\������������?��c����2 1�KԿX�Tx�x��3 1�����nY�S4 1�'9K��/�'/�S5 1���/�/�/�/>:/S6 1�Q/c/�u/�/-??Q?�/S7 1��/�/
?D?�?��?�?d?S8 1� {?�?�?�?WOBO{O�?�SMASK 1����L��O�D�GXNO����F&�^��MOT�EZ�Ż��Q_ǁ��%]pA݂��PL_�RANG!Q]�_QO�WER �ŵ��P1VSM_DRY�PRG %ź%�"O�_�UTART ��^�ZUME_�PRO�_�_4o��_�EXEC_ENB�  J�e�GSP�D`O`WhՅjbTD�Bro�jRM�o�hI�NGVERSIOoN Ź#o��)I_AIRPU�RhP �O(�MMKT_�@T�P#_À�OBOT_ISO�LC�NTV@A'q^huNAME�l��o��JOB_ORD_�NUM ?�X�#qH768w  j1Zc@�r�
�rV�s��r�?�r�?�r�pÀPC_OTIMEu�a�xÀoS232>R1��� LTEA�CH PENDA1Nw�:GX�!O� Mainte�nance CoKnsj2����"���No Use B�׏������1�C�y�V�NPO�P@�YQ��cS�CH�_L`�%^ �	�ő��!UD1�:럒�R�@VAI�L�q@�Ӏ�J�QS�PACE1 2�ż ��YRs�i��@Ct�YRԀ'{��8�?��˯� ���"���7�2�c�u� ����G���߯ѿ򿵿 �(��u�AC�c�u� ����Ͻ�߿���ϵ� �(��=�_�qσϕ� C߹������߱��$� �9�[�m�ߑߣ�Q� �����߭��� ���	� W�i�{���M����� ��5���.S�e� w�����I������ �*?as� �E�����/ &//;/]o��� ���/2/�/?"?�/ 7?Y/k/}/�/�/O?�/ �/�?�?�?O0OOK�A��*SYPpM�*�8.3026�1 yB5/21/�2018 A ��WPfG|�H�_T�X`� !$CO�MME�$�USAp $ENABLEDԀ�$INN`QpIO�R�B�@RY�E_SOIGN_�`�AP�AsIT�C�BWRK�B=D<�_TYP�CRINDXS�@W�@�%VFRI{�_GR�PԀ$UFRAyM�rSRTOOL\V�MYHOL�A$�LENGTH_V{TEBTIRST�T�  $SEC�LP�XUFINV_�POS�@$M�ARGI�A$WgAIT�`�ZX2�\��VG2�GG1�AI �@�S�Q	g�`_WR�B�NO_USE_DyI�BuQ_REQ�B�C�C]S$CUR�_TCQP�R"a^f ��GP_STAT�US�A @ `�A3`�BLk�H$zcQ1�h�P@���@_�F�X �@E_�MLT_CT�CH�_�J�`CO�@OLt�E�CGQQ$W�@�w�b#tDEAD�LOCKuDEL?AY_CNT�a3q�Gt�a$wf 2W R1[1$X�<�2[2�{3[3 $Zwy�q%Y�y�q%V�@��c�@�b$V�`�RV��UV3oh>b�@ Ǡ �d�0arMS	KJ�LgWaZ�C`NR�K�PS_RATE�0$���S
`�Q�T;AC��PRD���e��S*��a4�b  :�DG�A 0�P�f�lp bquS2�ppI�#`
`�P 
��S\`  ؾA�R_ENBQ ��$RUNN�ER_AXI�<`A�LPL�Q�RU�THI�CQ$FLIP�7��DTFEREN|��R�IF_CHS�U�IW��%V)�G1�����$PřA�Q�Pnݖ_JF�PR_P��	�RV_DA�TA�A  =$�ETIM���_$VALU$�	��OP_   ��A  2 ��SC*�	�� �$ITP_0!�SQ]PNPOU}�o��TOTL�o�DSP>��JOGLIb��P'E_PKpc�Of�i���PX]PTAS��$KEPT_MI�R��¤"`M�b�A	Pq�aE�@�y�q��g@١c�q�PG�BCRK6�x���L�I��  ?�SJ�q�P��ADEz�ܠBSO�Cz�MOTNv�D�UMMY16Ӂ�$SV�`DE_O�P��SFSPD_�OVR
���@L�D����OR��TP8�LE��F������OV��SF��F����bF�d�ƣ&c)�fQ~c�LCHDLY��RECOV���`���W�PM��gŢ�ROȲ�����_F�?� �@v�S �NVER\�@�`OFS�PC,�CSWDٱc�ձ���B,����TRG�š�`�E_FDO��MB�_CM}���B��BALQ�¢	�Q�̄VzaF�BUP�g��G
��AM���@`KՊ�fe�_M!�d�AMf�<Q��T$CA����uDF���HBKd��v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�Dd�9�1A��9�3A�^��ATIO�0���͠��US����WaAB��R+c�`tá`Dؼ�A��_AUXw�S�UBCPUP���S �`����3Եжc����3�FLA�B�HW�_Cwp"�Ns&�]sA�a��$UNIT�S�M�F�ATTR�Iz�Z�CYCL��CNECA���F�LTR_2_FI~��TARTUPJp0����A��LP����ޖ�_SCT*cF_�F�F_P���b�FS8��+�K�CHA/Q��p*�d�RSD��`Q����Q���_TH��PROr���հEM�PJ���G�T�c �Q�DI�@~y�RAILAC/��bMX�LOf�xS���ځ���拁���P�R#�S`app�C�� 	��FUsNC���RIN``QQP� ԱRA)]R ��AƠ��AgWAR֓��BLZa�WrAkg�ngD�AQ�B�rkLD@�र&q�M�K����TI���j���$�@RIA_SWV��AF��Pñ#���%%�p9r1��MO9IQ���DF_~P(��PD"LM-�FA��PHRDY�DORG�H; _QP�s%MULSE~Pz���**�� J��Jײ���FAN_ALMsLVG��!WRN�%�HARDP��UcO��� K2$SHADOW]�kp�a02��N� STOf�+�_^�w�AU{`R��eP_SBR�z5���:�F�� �3MPIN�F?�\�4��3R3EGV/1DG�+c1Vm �C�CFL(��?�DAiP���Z`Ɨ� �����Z�	 ��P(Q$�A$�Z�Q V�@�[�
7� ��EG߀o����kAAR���㌵2p�axG��AXE��wROB��RED���W�QD�_�Mh�SY�A��AF��FS�GWRqI�P~F&�STR��(��E�˰EH�)��D�a\2kPB6P��=V���Dv�OTO�1)���ARYL�tR��v�3���FI&�ͣ$LINKb!\��Q%�_3S���E�N�QXYZ2�Z5�V'OFF���R�R�X%xPB��ds�G�cFI�03g�h������_J���'�ɲ�S&qR0LTV[6����aTBja�"�bCL���DU�F7�TUR� X��e�Qb�2XP�ЊgFL�@E���x@�`�U9Z8��^�� 1	)�K��	Mw��F9��劂����ORQj��G;W3���#�Ґd ���upz����1�tOVE�q_�M��ё?C�uEC�u KB�v'0�x-�wH��t ���& `��qڠ� B�ё�u�q�wh�ECh�L���ER��K	�!EP����AT�K�6e9e�W���AXs�'��v�/�R  ����!�� ��P ��`��`�3p�Yp�1�p�� �� � � (�� 8�� H�� X� � h�� x�� ������oDEBU�$`%3�I��·RAB�ȱ�ٱ�sV��� 
d�J、��@񘧕� ������Q���a���a ��3q��Yq+$�`%"<�.cLAB0b�u��'�GRO���b<��B_s��"Tҳ*`��0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθu�ݸ��PNT0����SERVE �Z@� $`EAV�!�PO����nP!��P@�$!Y@ w $>�TRQ�b�
=��BG�K�%"2�\��� _ � l��5�D6ERRVb(�I��V0`;���'TOQ:�7�L�@
�(R��e G�%�Q��q <�50F� ,��`�z�>�RA� �2 d!�����S�  M��px�U ����OCuG��  ��COU�NT6Q��FZN_wCFGF� 4#��6��TG4�_�=������Î�VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@HE�L�0�� }5b`B_BAS��RSR�6�CSHH����1�Ǌ�2��U3��4��5��6���7��8��}�ROO0����P�PNLEA�c�AB)ë ��ACK�u�INO�T��(B$�UR0� =�_PUX��!0��OU+�Pd��8j��� V��TPFWD_KAR��L� ��RE(ĉ P�Pܺ>QUE�:RO �p�`r0P1I� x��j�P�f��6�QSE�M��0��� A��S�TYL�SO j�D�IX�&�����S!_�TMCMANRQ܉�PENDIt$�KEYSWITCaH���kHE�`�BEATM83PE�{@LE��>]��Uү�F��SpDO/_HOM# O�@�EF�pPRaB�A#PY�C� O�!��яOV_M|b<0 I�OCM�dFQ���h�HKYA DH�Q�7��UF2��M�x��p�cFORC�3gWAR�"�OM|@  @S�#o0UU)SP�@1�2&E3&4E���T�O���L���8UNLiOv�D4K$EDU1�  �SY�HD�DNF� M�B�LOB  p�SNPX_AS�҇ 0@�0��81�$SIZ�1$V�A{���MULTI�P-��# A�? � $��� H/4`�BS��0�C����&FRIFBO�S����3� NF�ODBUP߰�%@3;9�(�����Z@ x6��SI��TEs�r.�cSGL�1T�Rp�&�Н3B��@�0ST�MTq�3Pg@VByW�p�4SHOW�5n@�SV��_G��; 3p$PCJ�PЬ����FB�PHS�P AW�EP@VD|�0WC� ���A00��PB XG �XG XG$ XG5VI6�VI7VI8VI9VIAVIBVI�XG�YF�0BXGFVH��XbI1oIU1|I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1YU1Y2UI2bI2oI2|I2�I2�I�`�XP�I2p�X�I2�I2�IU2�I2�I2Y2Y��p�hbI3oI3|I3��I3�I3�I3�I3��I3�I3�I3�I3��I3�I3Y3Y4��i4bI4oI4|I4��I4�I4�I4�I4��I4�I4�I4�I4��I4�I4Y4Y5��i5bI5oI5|I5��I5�I5�I5�I5��I5�I5�I5�I5��I5�I5Y5Y6��i6bI6oI6|I6��I6�I6�I6�I6��I6�I6�I6�I6��I6�I6Y6Y7��i7bI7oI7|I7��I7�I7�I7�I7��I7�I7�I7�I7��I7�I7Y7T�ցVP� UD��y"ՠ��
<A62��t�R��CMD� ��M5�Rv�]��Q_h�R���e�����<�YSL���  � �%\2��+4��'��W�BVA�LU��b��'���F�H�ID_L���H�I��I���LE_���㴦�$0C�S�AC�! h ��VE_BLCK���1%�D_CPU5ɧ 5ɛ ������C�� ��R " � PWj��#06��LA�1SBћ������RUN_FLG�Ś����ĳ ����������H���ХĽ��TBC2��#/ � @ B��e ��S�8=�FTD	C����V���3dՆQ�THF�����R��L�ESERVE9��F��3�2�E�|�Н�X -$��LEN9��F��f�cRA��W"G�W_5��b�1��д2�MO$-�T%S60U�Ik�0�`ܱF����[�DEk�21LACEi0�CqCS#0�� _MA� pj��z��TCV����z�T�������.B i�'A�z�'AJh�#E�M5���J��@@i�V�z���2Q �0&@�o�h��JK��VK�9��{���щ�J0l����JJ��JJ��AAL���������e4��5�ӕ N1��P����.�LD�_�1�* �CF�"%{ `�GROU��(�1�AN4�C�#m ?REQUIR���EBU�#��6�$Tk�2$���z�܏ #�& \�AP�PR� C� 0�
$�OPEN�CLO�S�St��	i�
\��&' �Mf�p����W"-_MG�7CB@�A���B�BRK@NOLD|@�0RTMO_5�H�p1J��P�� ������������6��1�@ �m1�#�(� ������'��+#PATH''@!6#@!��<#� � '��1SCaA���6IN�ңUCJ�[1� C0@UM�(Y ��#�"������*���*��� PAYwLOA~J2LؠOR_AN^�3L���91�)1AR_F�2LSHg2B4LO�4�!F7�#T7�#ACRL_�%�0�'�$r��H��.�$HA^�2FLEX��J!�) P�2�D��߽���0��* :����z�FG]D��`��z���%�F1]A �E�G4�F�X�j�|���BE���������� ��(��X�T*�A���@�XI�[�m�\At�T$g�QX<�=��2TX ���emX���������� ��������+	�J>+ �-�K]o|�٠AT�F�4�CELFPѪs�J� �*� JEmCTR��!�ATN�vzH�AND_VB.���1��$, $8`Fi2Av���SWu�	#-� $$M*0.�]W�lg��PZ����A��� 1�����:AK��]A�kAz��LN�]D*kDzPZ G��C�CST_K�lK�N}DY��� A����0 ��<7]A<7W1�'��d�@g`�P��������"
"J"�. M�2D%"��H�����ASYMj%0��� j&-��-W1�/_ �{8� �$�����/�/�/�/ 3J<�:p9�/�89�D_VI��v����V_UN!I�ӛ��cD1J���� ╴�W<��n5Ŵ�w=�4��9��?�?<�uc$�4�3��%�H����/�j��0�DIzuO�ğ�k�>�0 �`��I��A ��#���@ģ���@���IPl� 1 �[ /�ME.Qph��9�ơT}�PT� ;pG �+ Gt� ����'��T�0 �$DUMMY1���$PS_�@RMF�@  G b�'7FLA@ YP(c|���$GLB_T P�ŗ���9 P�q���2 X� z!SuT9�� SBRM �M21_V�T$_SV_ER*0O�pL����CL����AGP�O��f�GL~�EW�>�3 4H �$YrZrW@�x�A1B+�A���"	""�U&�4 8`NZ�"�w$GI�p}$&�� -� �Y�>�5 qLH {��}$F�E��NEAR(PN��CF��%PTANC��B	!JOG�@� �6.@$JOI�NTwa?pd�MSE]T>�7  x�E��HQtpS{r��up>�8�� �pU.Q?��� LOCK_F�OV06���BGLV��sGLt�TEST�_XM� 3�EMP������_�$1U&@%�w`24� Y�B��5��2�d��3���CE- ���� $K�AR�QM��TPD�RA)�����VECXn@��IU��6��{HEf�TOOL�C�2V�DRE IS�3ER6��@AC)H� 7?Ox ӦQ�29Z�H I� � @$RAIL__BOXEwa�oROBO��?��?HOWWAR�1�<_�zROLMj���:qw�jq� �@ O{_Fkp! d�tl>�9�� �R �O8B: �@��c�OU�;�Һ�3�ơ�r�q_�$PIP��N&`H�l�@���#@CORDEADd�p >f�fpO�� < D ��OB⁴sd���K�p����qSYS��ADR�qf��TC}Ht� = ,8`SENo��1Ak�_{��-$Cq,Be�VWV�A��> � � &��PREV_�RT�$EDI}Tr&VSHWRkq��֑ &R:�v�D���JA�$�a$H�EAD�6�� ��z#KE:�E�CPS�PD�&JMP�Ld~��0R*P��?�T�1%&I��S�rC�p�NE; �q�wTIC�K�C��M�13�3H=N��@ @� 1Gu�!_GPp6��0gSTY'"xLO���:�2l2?�A t 5
m G3%%$R!{�u=��S�`!$�� w`���ճ���Pˠp6�SQU��E��u�T�ERC�0��TSUtB ����hw &`gw�Q)�pO���F�@IZ��{��^уPR�kюB1XP9U���E_DO��, �XS�K~�AXI4�@���UR�pGS@�r� ^0�&��p_) �ET�BPm��o�%�0Fo��0A|���CRԍ��a  z1@R�Cl>@ P��b_�yUr��Y��yU ��yS��yS���UЇ�U ���U���U�]��Ul [��Y�bXk�]Cm�h����0ASC��� D h�DS�~0��Q�SP���eA	Tހ���A]0,2NҿADDRES<B�} SHIF{s��_W2CH�p�I�Ю=q�TVsrI��E�"���a�Ce�
��
�;�VW�A��F \��q��0l|\A@�rC�_B"R{zp�ҩq��TXSCREE��Gv��1TIN!A���t{����A�b?�H T1�ЂB �����I��A��BE�y RRO������ �B��D��UE4I ��g�!p�S��R�SM]0�GUNEX0(@~Ƴ�j�S_S�ӆ@��Á։񇣣�ACY򼯂0� 2H�pU�E;�J�����@G+MT��Lֱ�A�нO	�BBL_| W�8���K ��0s�OM��LE/r��� �TO!�s�RIGHΓ�BRD
�%qCKsGR8л�TEX�@|����WIDTH��� �B[�|�<��I�_��Hi� L 	8K���_�!=r���R:�_��Yґ��)O6q�Mg0紐�U��h�Rm��LUqMh��FpERVwD �P���`�N���&�GEUR��F4P)�)� LP��(R	E%@�a)ק�a�!���f �5�6�7�8Ǣ#B�É@���t�P�fW�S@M��USR&�O �<����U�Qs�FsOC)��PRI;Q�m� :���TRIP>�m�UN����Pv��0��f%��'8���@�0 Q���.�AG �0T� �aL>q�OS�%�RPo���8�R/�A�H�L4����U¡�S�U�g��¢5��OF�F���T�}�O�� 1R����ĝS�GUN��>6�B_SUB?���N,�SRTN�`TUg2���mCOR| D�R�AUrPE�TZ�#'��VCC��	3V �AC36MFB1�f$c�PG �W �(#��ASTEM�0����0PE��T3�G�X �\ ��M�OVEz�<���AN��� ���M���LIM_X��2��2�� 7�,�����ı�
��VF�`E���~��04Y��IB�7���5S��_Rp� 2���/ WİGp+@���}СP��3�Zx# ���3����A�ݠCZ�DRID����Vy08�90�� De�MY_UBYd���6��@��!q��X��P_S���3��L�KBM,��$+0DEY(#EX�`�����UM_MUb� X����ȀUS��� ���G0`PACI���а@��:��:0,�:����RE/�3qDL�+��:[��/TARG��P�rr��R<�\ d`�H�A��$�	��AR��#SW2 ��-��@�Oz�%qA7p�yRE�U�U�01�,�HK�2]g0�qP�� N� �EAM0GW�OR���MRC]V3�^ ���O�0M�C�s	���|�REF_���x (�+T� ������p���3_RCH 4(a�P�І�hrj�NA8�5��0�_ ��2�����L@��n�@@OU ~7w6���Z��a2[��RE�p�@;0�\�c�a'2K�@S+UL��]��C��0�3^��� NT��L� 3��(6I�(6q�(3� L��Q5��Q5I�]7q��}�Tg`4D`�0|.`0�AP_HUCv�5SA��CMPz��F�6�5�5�0_�aR ��a�1I\!X�9�@��VGFS��ad ��M��0p�UF_x��B� �ʼ,�RO��Q��'����U�R�3GR�`.�3I Dp���)�D�;�X�A��~�IN��H{D���V@AJ���S͓UWmi=�����LTYLO*�5���|�bt +�c�PA� �cCACH�vR�UvQ��Y���p�#CF�I0sF�R�XT���Vn+$H	O����P!A3󯂀XBf�(1 ���$�`V�Py� ^b_SZ3d13he6K3he12J�`eh chG�chWA�UsMP�j��IMG9�uPAD�iiIM�RE�$�b_SIZ©$P����0 ��AS�YNBUF��VR�TD)u5tqΓOLE_2DJ�Qu5R��%C��U��vPQu�ECCUlVEM�V �U�r�WVIRC�aIuVTPG���r`v1s��5qMPLAq�a��v�V0�cm�� CKLAS�	8�Q�"��d  �ѧ%$ӑӠ@}¾�$�Q���Ue |�0!�rSr�T�#0! �r�iaI��m�vK�BG��3VE�Z�PK= �v8�Q�&�_HO�0��f � >֦3�@<Sp�SLOW>�{RO��ACCE���!� 9�VR�#���p�:���AD�����PQAV�j�� D�����M_B"���^�JM�PG ��g:�#E$SSC��F�vPq���hݲvQS�`qVN���LEXc�i �T`�sӂ��Q�F�LD �DEsFI��3�02���:��V�P2�Vj� �A��V�4[`MV_PIs��t���A�L�@��FI��|�Z�� Ȥ�����A���A��~�sGAߥ1 LOO��1 JCB���Xc��<^`�#PLANE��R��1F�c�����p�r�M� [`�噴��S ����f����Af��R�A�w�״tU��pRKyE��d�VANC��A���� k����ϲϡ�R_AA� l��2� ��p�#B��m h���O K��$������kЍ0O)U&A�"A�
p�p�SK�TM@FVIEM 2l ��P=���n <<��dK�/UMMYK1P���`D��AC�U��#AU��o �$��TIT�g$PR����OP���VSHIF�r�p`J�Qs�ؙ�fOxE$� _R�`U�#����s��q ������G�"G�޵'�9T�$�SCO{D7�CNTQ i�l�>a� -�a�;�a�H�a�V����1�+�2u1��Dx����  D�ЋMO�Uq��a�J,Q�����a_�R[�ir�n�*@LIQ��AA/`�XVR��s��n�TL���ZABC�t�t�c�]
AZIP��u撖��LVbcLn"�^��MPCFx�v:��$�� ���DMY_LN�������@y�w Ђ(a�u� �MCM�@CbcCA�RT_�DPN� �$J71D ��=NGg0Sg0�B�UXW� ��UXE#UL|ByX@���	��|!Z��x 	���m��YH�Db  y �80���0EIGH��3n�?(� H����$z ���|������$B� Kd'��_X��L3�RVS�F`���OVC�2' �$|�>P&��
q����5D�TR�@ �V�c��SPHX��!{� ,� *<�$�R�B2 2 ����C!�?  �@V+�| b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/?�/�/V(7%3@/R/d/ v/�/6?�/�/�?�?�? O4OOION;4]?o? �?�?�?SO�?�?�O_@�O0_Q_8_f_N;5zO �O�O�O�Op_�O_o�8o�_MonoUo�oN;6 �_�_�_�_�_�oo%o 4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8�����Ǐ =�_�n���R���ş���ڟN;G �S џ�
���� ��W�i�{������� ï�.�������A��dW�<�N�|��� ����Ŀֿ�ޯ�� �0�B�_�R�d�꿤� �������������� *�L�^��rτ�
��� ���������&�8߸J�l�~� `ҟ @�з����ߩ��-����&�,�� �9�{�����a����� ����������A 'Y������ ���a#1��
��N;_MOD�E  ��S ���[�Y� B���
/\/*	|/�/�R4CWORK_A�D�	�A�T1R  ���� �/�� _INTVAL��+$��R_OPoTION6 ��q@V_DATA_GRP 27���D��P�/~?�/ �?�9��?�?�?�?O O;O)OKOMO_O�O�O �O�O�O�O_�O_7_ %_[_I__m_�_�_�_ �_�_�_�_!ooEo3o ioWoyo�o�o�o�o�o �o�o/eS �w������ �+��O�=�s�a��� ����͏���ߏ���9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_TI�M����ΑR ���Ƙ��5�;#U!AP"�Z���� �? E�W�i�{�����.�ï�կ�����'(�~�T"2F��Q�dDF�a��2�o+@a�@������)�u��� k0~ϴ��_ ��  T� � �2�D�~)�T D��Q� zόϞϰ��������� 
��.�@�R�d�v߈���/V凷������߽��R�;W�o �W�p���
�t��Di�z$� �0 � �T"%!������ ������������ *�<�N�`�r������� ��������&8 J\n����� ���"4FX ��࿁���� ���/`4�=/O/ a/s/�/�/�/�/�/�/�!!/ �0޲k�ݵu� 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  ok$o6oHoZolo~o �o�o�o�o1/�o�o  2DVhz�/5 ?�������� &�8�J�\�n������� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q�0c�u��� ���`� ��ϯ����)�;� M�_�q���������˿ݿ� ����3� ���&2,��	�1234567�8v�h!BW!��2�Ch���0�ϵ��������� �!�3�9ѻ�\�n߀� �ߤ߶���������� "�4�F�X�j�|�h�K� ����������
��.� @�R�d�v��������� �����*<N `r������ �&��J\n �������� /"/4/F/X/j/|/; �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�/�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_�?L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o =_�o�o�o�o�o�o  2DVhz�����h�������u�o.�@�R���C�z  B��  � ���2&� �� _�
���/  	�_�2�Տ�����_�p������ďi�{����� ��ß՟�����/� A�S�e�w��������� N������+�=�O� a�s���������Ϳ߿����'�9�K�_�������<v�_��$�SCR_GRP �1
� �� t ���� ��	 _����� �����������_���p���)�a����~&�DE� DW8����l�&�G�CR�-35iA 90�12345678�90��M-20���8��CR35 ��:�
��������������:֦� Ӧ�G���&������	��]�o����~:���H���>�����������&���ݯ:��j���`��g������B�t�!���������A�����  @�`��@�� ( ?�=��H�t�P
��F@ F�`z�y��� ��� �$H ��Gs^p��B��7��/� 0//-/f/Q/�/u/�/ �/�/8���P�� 7%?����"?W?-2?<5��]? H�14�?t�ȭ7�������?-4A, �&E$@�<�@G�B-1A 3OZOlO-:HA�H��O�O|O P�B(��B�O�O_��EL_�DEFAULT � �����`SHOTS�TR#]A7RMIP�OWERFL  �i�/UYTWFD�O$V /URRV�ENT 1�����NU L!DUM_EIP_�-8�j!AF_�INE#P�_-4!�FT�_->�_;o!���`o �*o�o!�RPC_MAI�N�ojh�vo�o�cV�IS�oii��o!7TPpPU�Y�dk!
PMON_PROXYl��VeZ�2r��]f���!RDM_'SRV��Yg�O�G!R��k��Xh>����!
�`M��\i����!RLSY3NC�-98֏3��!ROS�_-<�y4"��!
CE4p�MTCOM���Vk�n�˟!	��CON�S̟�Wl���!>��WASRC��V�m�c�!��US	Bd��XnR���Noӯ �������!��E���i�0���WRVICE_KL ?%�[� (%SVC�PRG1��-:Ƶ2�ܿ�˰3�	�˰4�,�1�˰5T�Y�˰6|ρ�˰7�ϩ�˰��$���9����ȴf� !�˱οI�˱��q�˱ ϙ�˱F���˱n��� ˱���˱��9�˱�� a�˱߉��7߱�� _��������)� ���Q����y��'� ���O����w���� ������˰�� İd�c����� �=(as^ ������/� /9/$/]/H/�/l/�/ �/�/�/�/�/�/#?? G?2?k?V?}?�?�?�? �?�?�?O�?1OCO.O gORO�OvO�O�O�O�O��O	_�O-_��_DE�V �Y��MC:5Xd�>GTGRP 2SVK ���bx 	�/ 
 ,�P5_�_ �R�_�_�_�_�_�_3o oWo>o{o�oto�o�o �o�o�o�o/A�_ e������ ��� �=�$�6�s� Z���~���͏���H �'�ޏK�2�o���h� ����ɟ۟���#� 5��Y�@�}�d�v��� 
�ׯ�Я���1�� *�g�N���r������� �̿	���?�&�c� u�̯��PϽ��϶��� ���)��M�4�q�X� jߧߎ��߲������ %�|��[���f�� ������������3� �W�i�P���t����� ����>�A( eL^����� �� =O6s Z�� ���/ �'//K/]/D/�/h/ �/�/�/�/�/�/�/#? 5??Y?�N?�?F?�? �?�?�?�?O�?1OCO *OgONO�O�O�O�O�O`�O�O�O_kT �"V		_R_=_v_a_�_�_��_�[%��_�_�S���a�Qeo)g oIo7omo[o�o�i�_ �oi�o�o�o% '9o�o��o_� �����!�w� n��G�����ŏ��� ׏�O�4�s���g��� w����������'�� K�՟?�-�c�Q�s��� �������#����� ;�)�_�M�o���ׯ�� �����ݿ��7�%� [ϝ��ϔ�K�m�Gϵ� �������3�u�Zߙ� #ߍ�{ߝߟ߱����� �M�2�q���e�S�� w������%�
�I� ��=�+�a�O���s��� �����!���9 ']K������q �m��5#Y ���I���� �/�1/sX/�!/ �/y/�/�/�/�/�/	? K/0?o/�/c?Q?�?u? �?�?�??�?O�?�? �?)O_OMO�OqO�O�? �OO�O_�O__%_ [_I__�O�_�Oo_�_ �_�_�_oo!oWo�_ ~o�_Go�o�o�o�o�o �o	_o�oV�o/� w�����7� [�O��_���s��� ��͏��3���'�� K�9�[���o����̟ ������#��G�5� W�}������m�ׯů �����C���j�|� 3�U�/���ӿ����� �]�Bρ��u�cυ� �ϙ��Ͻ���5��Y� ��M�;�q�_߁߃ߕ� �����1߻�%��I� 7�m�[�}�������	� ������!��E�3�i� �����Y���U����� ��A��h��1 ������� [@	sa�� ����3/W� K/9/o/]/�/�/�/� �/�/�/�/�/?G?5? k?Y?�?�/�?�/?�? �?�?�?OCO1OgO�? �O�?WO�O�O�O�O�O �O	_?_�Of_�O/_�_ �_�_�_�_�_�_G_m_ >o}_oqo_o�o�o�o �o�ooCo�o7�o Gm[���o� ���3�!�C�i� W�������}��Տ ���/��?�e����� ˏU������џ��� +�m�R�d��=���� ����߯ͯ�E�*�i� �]�K�m�o������� ۿ��A�˿5�#�Y� G�i�k�}ϳ������ �����1��U�C�e� ���ϲ��ϋ�����	� ��-��Q��x��A� ��=���������)� k�P������q����� ������C�(g��� [Im����  ?�3!WE {i������ ��///S/A/w/� �/�g/�/�/�/�/�/ +??O?�/v?�/??�? �?�?�?�?�?�?'Oi? NO�?O�OoO�O�O�O �O�O/OUO&_eO�OY_ G_}_k_�_�_�__�_ +_�_o�_/oUoCoyo go�o�_�oo�o�o�o 	+Q?u�o� �oe������ '�M��t��=����� ˏ���ݏ�U�:�L� �%���m�����ǟ�� �-��Q�۟E�3�U� W�i�����ï��)� ����A�/�Q�S�e� ��ݯ¿������� �=�+�Mϣ�ɿ��ٿ s��ϻ�������9� {�`ߟ�)ߓ�%ߣ��� �������S�8�w�� k�Y��}������� +��O���C�1�g�U� ��y��������'��� 	?-cQ��� ��w�s� ;)_���O� ����//7/y ^/�'/�//�/�/�/ �/�/?Q/6?u/�/i? W?�?{?�?�?�??=? OM?�?AO/OeOSO�O wO�O�?�OO�O_�O _=_+_a_O_�_�O�_ �Ou_�_�_o�_o9o 'o]o�_�o�_Mo�o�o �o�o�o�o5wo\ �o%�}���� �="�4����U� ��y�����ӏ���9� Ï-��=�?�Q���u� ���ҟ�����)� �9�;�M���ş��� s�ݯ˯��%��5� ��������[�����ٿ ǿ���!�c�Hχ�� {�ϋϱϟ������� ;� �_���S�A�w�e� �߭ߛ������7��� +��O�=�s�a��� ���������'�� K�9�o������_��� [�������#G�� n��7����� ��aF�y g������9 /]�Q/?/u/c/�/ �/�/�%/�/5/�/)? ?M?;?q?_?�?�/�? �/�?�?�?�?%OOIO 7OmO�?�O�?]O�O�O �O�O�O!__E_�Ol_ �O5_�_�_�_�_�_�_ �_o__Do�_owoeo �o�o�o�o�o%o
 �o�o�o=sa����o�!+q�$S�ERV_MAILW  +u!����OUTPUT��$�@�RV �2�v  $� �(�q�}��SAV�E7�	�TOP10� 2W� d 'ݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w����������ѿ�u��Y�P���FZN_C�FG �u�$�~����GR�P 2�D� ?,B   A[�+q�D;� B\���  B4~�R�B21��HELL���u��j�k��2�����%RSR �������
�C�.�g� Rߋ�v߈��߬������	���-�?�Q��  �_�%Q���(_���,p��⦼�ޖ�g�2,pd�����HK 1�� ��E�@�R� d��������������� ��*<e`r����OMM ������FTOV_�ENB�_���HO�W_REG_UI��	�IMIOFW�DL� �^�)WAIT���$V�1�^�NTIMn���VA�|_)_UNIT����LCTRY�B��MB_HDDN 2W� 2�:%0 �p Q/�qL/^/�/�/�/�/�/�/�/�"!ON_�ALIAS ?e�	f�he�A?S? e?w?�:/?�?�?�?�? �?OO&O8OJO�?nO �O�O�O�OaO�O�O�O _"_�OF_X_j_|_'_ �_�_�_�_�_�_oo 0oBoTo�_xo�o�o�o �oko�o�o,�o Pbt�1��� ����(�:�L�^� 	���������ʏu��  ��$�Ϗ5�Z�l�~� ��;���Ɵ؟�����  �2�D�V�h������ ��¯ԯ���
��.� ٯR�d�v�����E��� п���ϱ�*�<�N� `�r�ϖϨϺ���w� ����&�8���\�n� �ߒߤ�O��������� ��4�F�X�j�|�'� ������������ 0�B���f�x������� Y���������> Pbt���� ��(:L� p����c��  //$/�H/Z/l/~/ )/�/�/�/�/�/�/?� ?2?D?V?]3�$S�MON_DEFP�RO ����1 �*SYSTEM�*0m6RECA�LL ?}9 �( �}-cop�y frs:*.�dt virt:�\temp\=>�147.87.1�49.40:8008 �5�?OO*O�}
xyzrate 61 �?�?�?O�O�O6E?GXOj@@^OpO__%_8C8�6�orderfil�.daKFmpba�ckWO�O�_�_�_ �}/�2mdb�0*�T_f_o_ oo$o7D3x�4:\�_I`�_�Ap�_�o�o�o }4?eaGoYo�Eto) <_N_�_�_����_ U�_p��%�8o�o �ono������oG�Y� �o���!�4F�j {�������_���� ��0�B�Տf�w��� ������Q��v������:�4h:\su�pportɨI�=�>2611609�60:56058�9+�����/Ltp?disc 0߯�@�\�n����#�6Et�pconn 0 �ȿڿ�}Ϗϡ�4G=���olptest.tpLI��ǿ��� �0�B�˟���ωߛ� ����[��v���� >�ѯg��߅��Ｏ M�_��x�	��.O@G ������������O�N2552 ^�p� %��������� �6�HZl�!<����:731�� ��6J�l� /!/�F�����/ �/1�C���Mx/	?? �����/S�/�?�?�? 7�H?\�Xs?OO(O ���?�?[�?�O�O�O �/�/W?r?__'_:? �O^?�O�_�_�_�?KO ]O�?�_o#o6O�_�_ lO}o�o�o�O�OO_�O �o2_D_�oh_�o����z�$SNP�X_ASG 2�����q�� P 0 �'%R[1]�@1.1��y?��s%�!��E�(�:� {�^�������Տ��ʏ ���A�$�e�H�Z� ��~���џ����؟� +��5�a�D���h�z� ����ů�ԯ���
� K�.�U���d������� ۿ������5��*� k�N�uϡτ��ϨϺ� �����1��U�8�J� ��nߕ��ߤ������� ���%�Q�4�u�X�j� ������������� ;��E�q�T���x��� ��������% [>e�t��� ���!E(: {^������ /�/A/$/e/H/Z/ �/~/�/�/�/�/�/�/ +??5?a?D?�?h?z? �?�?�?�?�?O�?
O KO.OUO�OdO�O�O�O �O�O�O_�O5__*_ k_N_u_�_�_�_�_�_ �_�_o1ooUo8oJo��ono�o�o�d�tPA�RAM �u}�q �	��jUP�d9p�ht���pOFT_KB_CFG  �c��u�sOPIN_S_IM  �{v�n��p�pRVQSTP_DSBW~�r"t�HtSR �Zy � &� ZERO S�T���vTO�P_ON_ERR�  uCy8�PT�N Zuk��A4�RINGo_PRMB� �`�VCNT_GP �2Zuq�!px 	r��ɍ���׏���wVD��RP 1	�i p�y��K� ]�o���������ɟ۟ ����#�5�G�Y��� }�������ůׯ��� ��F�C�U�g�y��� ������ӿ��	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�qߘߕߧ߹��� ������%�7�^�[� m����������� ��$�!�3�E�W�i�{� �������������� /ASew�� �����+ =Ovs���� ���//</9/K/ ]/o/�/�/�/�/�/�/ ?�/?#?5?G?Y?k? }?�?�?�?�?�?�?�?�OO)�PRG_CgOUN�:t�k��GuKBENB��FEM�pC:t}O_UPD �1�{T  
 4Or�O�O�O__!_ 3_\_W_i_{_�_�_�_ �_�_�_�_o4o/oAo So|owo�o�o�o�o�o �o+TOa s������� �,�'�9�K�t�o��� ������ɏۏ���� #�L�G�Y�k������� ��ܟן���$��1� C�l�g�y��������� ӯ����	��D�?�Q� c���������ԿϿ� ���)�;�d�_�q��=L_INFO 1��E�@ �2@����������� ��8@�oA˛Mˋ�´*�H@Y?SDEBUGU@�@����d�If�SP_�PASSUEB?~x�LOG  �ƕ�C��Qؑ� � ��A��UD�1:\��Uߦ�_M�PC�ݵE&�8�A���V� �A�SAV !�������X����SVZ�TE�M_TIME 1u"���@ 0����X�X������$�T1SVGUNS��@VE'�E��A�SK_OPTIO�NU@�E�A�A+�_�DI��qOG�BC2_GRP 2#�I������@�  C����<Ko�CFG 3%z��� ���`��1�.> dO�s���� ���*N9r ]��������/�8/#/\/n/v$ Y,�/Z/�/�/H/�/? �/'??K?]�k?=�@0 s?�?�?�?�?�?�?O �?OO)O_OMO�OqO �O�O�O�O�O_�O%_ _I_7_m_[_}__�_ �_�X� �_�_oo/o �_SoAoco�owo�o�o �o�o�o�o=+ MOa����� ����9�'�]�K� ��o���������ɏ�� �#��_;�M�k�}��� �����ß�ן�� 1���U�C�y�g����� ����������	�?� -�c�Q�s��������� �Ͽ����)�_� Mσ�9��ϭ������� m���#�I�7�m�� ��_ߵߣ��������� ��!�W�E�{�i�� ������������� A�/�e�S�u�w����� ��������+=O ��sa����� ��9']K mo������ �#//3/Y/G/}/k/ �/�/�/�/�/�/�/? ?C?��[?m?�?�?�? -?�?�?�?	O�?-O?O QOOuOcO�O�O�O�O �O�O�O__;_)___ M_�_q_�_�_�_�_�_ o�_%oo5o7oIoo mo�oY?�o�o�o�o �o3!CiW�� ������� -�/�A�w�e������� ���я���=�+� a�O���s�������ߟ ͟��o�-�K�]�o� ퟓ�����ɯ���צ���$TBCSG_GRP 2&ץ��  ��� 
 ?�  6�H�2�l�V��� z���ƿ��������(�d�E�+�?�	 HC�=���>���G���~�C�  A�.��e�q�C��>ǳ3�3��S�/]϶�Y���=Ȑ� C\  B�ȹ��B���>�c���P���B�Y��z��L�H�0�$�����J�\�n�����@ �Ҿ���������=��Z�%�7����?3������	V3�.00.�	cr;35��	*�����
�������� �3��4�   �{�CT�v�}��J�2�)������C�FG +ץ�'� *������rI���� .<
�<bM�q �������( L7p[�� ����/�6/!/ Z/E/W/�/{/�/�/�/ �/.�H��/??�/L? 7?\?�?m?�?�?�?�? �? OO$O�?HO3OlO WO|O�O����Oӯ�O �O�O!__E_3_i_W_ �_{_�_�_�_�_�_o �_/oo?oAoSo�owo �o�o�o�o�o�o+ O=s�E��� Y�����9�'� ]�K�m�������u�Ǐ ɏۏ���5�G�Y�k� %���}�����ßşן ���1��U�C�y�g� ������ӯ������ 	�+�-�?�u�c����� �����Ͽ���/� A�S�����qϓϕϧ� �������%�7�I�[� ��mߣߑ߳����� �߷��3�!�W�E�{� i����������� ��A�/�e�S�u��� ������������ +aO�s�� e�����'K 9o]���� ���#//G/5/k/ }/�/�/[/�/�/�/�/ �/??C?1?g?U?�? y?�?�?�?�?�?	O�? -OOQO?OaO�OuO�O �O�O�O�O�O___ M_�e_w_�_3_�_�_ �_�_�_oo7o%o[o moo�oOo�o�o�o�o �o!3�o�oiW �{������ �/��S�A�w�e��� ����я������� =�+�M�s�a������� ��ߟ�_	���_ן ]�K���o�������ۯ ɯ���#���Y�G� }�k�����ſ׿���� ����U�C�y�g� �ϋ��ϯ�������� 	�?�-�c�Q�s�u߇� �߫��������)�� 9�_�M����/���� i������%��I�7� m�[������������� ������EWi{ 5������� �A/eS�w �����/�+/ /O/=/_/a/s/�/�/ �/�/�/�/?'?��?? Q?c??�?�?�?�?�? �?�?O�?5OGOYOkO�)O�O}O�O�O�O�N s �@S V�_R�$TBJO�P_GRP 2,��E� / ?�V	-R4S�.;\��@|�u0{SPU >���UT @��@LR	 �C�� �Vf  C����ULQLQ>�33��U�R����U�Y?~�@=�ZC��P׌�ͥR��P � B��W$o/gC���@g�dDb�^���eeao�P�&ff�e=�7L3C/kaB o�o�P��P�efb-C�p��^g`�d�o��PL�Pt<�eVoC\  �Q@�'p}�`�  A�o�L`�_wC�BrD�S�^�]�_�S~�`<PB��P0�anaa`C�;�`L�w�aQoxp��x�p:��XB$4'tMP@�PCHS��n���=�P����trd<M�gE�2pb ����X�	��1�� )�W���c�������� ����󟭟7�Q�;�PI�w���;d�Vɡ��U	V3.00�RScr35QT�*�QT�A�� �E�'E�i��FV#F"w�qF>��FZ�� Fv�RF�~�MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
�D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt���ٵ=�_t��V �R�p�V9� ]ESTP�ARtp�HFP*SH�R\�ABLE 1%/;[%�SG��Q �W�G�G�GȨ WQG�	G�
G��GȖ�QG�G�8G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ߱���w�S]�CS !ڄ�� �����������&� 8�J�\�n��������� ���� ]\�`��	� �(�:�����
��.��@�w�NUM  ��EEQ�P�	P ۰ܰw�_CFG 0��)r-P�IMEBF_TT�b��CSo�,VER�ڳ-B,R 1=1;[ 8��R��@� �@&   �������/ /)/;/M/_/q/�/�/ �/�/�/?�/?J?%? 7?M?[?m?>�@�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_l_�Y�@cY�MI_CWHAN8 c c�DBGLV��:�cX�	`ETHER_AD ?f�\`��?�_uo�oQ��	`ROUTV!�	
!�d�o�lSN�MASKQhcba255.uߣ'�9ߣY�OOLOF/S_DIb��U;i�ORQCTRL �2		�Ϸ~T �����#�5�G� Y�k�}�������ŏ׏ �����.��R�V��PE_DETAI�/h|zPGL_CONFIG 8�	����/cel�l/$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c� u�����(���ϯ�� ����;�M�_�q��� ��$�6�˿ݿ��� %ϴ�I�[�m�ϑϣ� 2����������!߰� ��W�i�{ߍߟ߱�%}F�������/�A��C�i�H�Eߞ�� ��������?��.�@� R�d�v���������� ������*<N` r������ �&8J\n� �!�����/ �4/F/X/j/|/�// �/�/�/�/�/??�/ B?T?f?x?�?�?+?�? �?�?�?OO�?>OPO�bOtO�O�O�O����User Vi�ew ��}}12�34567890 �O�O�O_#_5_=T�P,��]_���I2�I:O �_�_�_�_�_�_X_j_�B3�_GoYoko}o�o�o o�op^46o�o�1CU�ovp^5 �o�����	�h*�p^6�c�u����� �����ޏp^7R�� )�;�M�_�q�Џ��p^8�˟ݟ���%����F�L� lCamera�J ��������ӯ���E~��!�3��OM�_�`q��������y  e� �Yz���	��-�?�Q� ��uχϙ�俽���������>��e�5i�� c�u߇ߙ߽߫�d��� ���P�)�;�M�_�q� ��*�<��i������� ��)���M�_�q��� ��������������<� û��=Oas�� >����*' 9K]f�Q��� ����/�%/7/ I/�m//�/�/�/�/ n<��^/?%?7?I? [?m?/�?�?�? ?�? �?�?O!O3O�/<׹� �?O�O�O�O�O�O�? �O_!_lOE_W_i_{_�_�_FOXG9+_�_�_ oo(o:o�OKopo�o )_�o�o�o�o�o 
��	g�0�oM_q ���No����o �%�7�I�[�m�& l�n��Ə؏����  ��D�V�h������� ��ԟ柍�g�ڻ}� 2�D�V�h�z���3��� ¯ԯ���
��.�@� R���3uF�鯞���¿ Կ������.�@ϋ� d�vψϚϬϾ�e�w� ��U�
��.�@�R�d� ψߚ߬��������� ��*���w���v� �������w���� �c�<�N�`�r����� =�w��-����� *<��`r�����������  ��1CUgy��������   -/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E_W_i_�  
���(  �%( 	 y_�_�_�_ �_�_�_o	o+o-o?o@uoco�o�o�o�Z* �Q&� J\n������o ���9�(�:�L� ^�p���������܏ � ��$�6�}�Z�l� ~�ŏ����Ɵ؟��� C�U�2�D�V���z��� ����¯ԯ���
�� c�@�R�d�v������ ��п�)���*�<� N�`ϧ����ϨϺ�� ������&�8��\� n߀��Ϥ߶������� ��E�"�4�F��j�|� ����������� �e�B�T�f�x����� ��������+�, >Pb������� ���(o� ^p������ � /G$/6/H/�l/ ~/�/�/�/�//�/�/ ?U/2?D?V?h?z?�?�/�`@ �2�?�?��?�3�7�P��!�frh:\tpg�l\robots�\m20ia\c�r35ia.xml�?;OMO_OqO�O�O�O�O�O�O�O �� �O_(_:_L_^_p_�_ �_�_�_�_�_�O�_o $o6oHoZolo~o�o�o �o�o�o�_�o 2 DVhz���� ��o�
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟�ݟ� �&�8�J�\�n����� ����ȯߟٯ���"� 4�F�X�j�|��������Ŀ־�8.1 ��?@88�?�ֻ�ֿ�3�5�G� iϓ�}ϟ��ϳ����� ���5��A�k�U�w���߿��$TPGL�_OUTPUT �;�!�! ��������,� >�P�b�t����� ��������(�:�L�@^�p�������������2345678901�������� �"��BTfx� �4�����
}$L^p�� ,>��� //$/ �2/Z/l/~/�/�/:/ �/�/�/�/? ?�/�/ V?h?z?�?�?�?H?�? �?�?
OO.O�?<OdO vO�O�O�ODOVO�O�O __*_<_�OJ_r_�_ �_�_�_R_�_�_oo &o8o�_�_no�o�o�o �o�o`o�o�o"4 F�oT|����\��}�����0�B�T�e�@������� ( 	 �� Џ������<�*� L�N�`���������ޟ ̟���8�&�\�J� ��n���������ȯ���"�������*�X� j�F�����|�¿Կ�� C���ϱ�3�E�#�i� {�忇ϱ�S������� ���/ߙ�S�e�߉� ��y߿���;����� ��=�O�-�s���ߩ� ��]��������'��� �]�o���������� ��E�����5G% W}������g� ��1�Ug	 w�{��=O	/ /�?/Q///u/�/� �/�/_/�/�/�/�/)? ;?�/_?q??�?�?�? �?�?G?�?O�?OIO [O9OO�O�?�O�OiO �O�O�O!_3_�O_i_ {__�_�_�_�_�_�R��$TPOFF_�LIM >�op:���mqbN_�SV`  l��jP_MON M<6�dopop�2l�aSTRTC�HK =6�f�� bVTCOMP�AT-h�afVWV_AR >Mm�h.1d �o �oop�`ba_DEFPROG %|j?%ZERO	�o~$qISPLAY`�|n"rINST_M�SK  t| ~^zINUSER�o�dtLCK�|}{QU?ICKMEN�dtoSCRE�p6�~�btpscdt��q��b*�_.�S�T�jiRACE_�CFG ?Mi��d`	�d
?�~u�HNL 2@|i����k r͏ߏ ���'�9�K�]�w�ITEM 2A��� �%$1234567890����  =<��П��  !���p��=��c��^��� �������.���R�� v�"�H�ί��Я��� ���*�ֿ���r�2� ������4�޿�ϰ��� &���J�\�n���@ߤ� d�v��ς������4� ��X��*��@��� ���ߨ�������T� ��x������l��� �����,�>�P����� ��FX��d����� �:�p"� �o�����F 6HZt~��N/ t/�/��// /2/�/ V/?(?:?�/F?�/�/ �/j?�??�?�?R?�? v?�?QO�?lO�?�O�O O�O*O|O_`O _�O 0_V_h_�Ot_�O__ �_8_�_
oo�_@o�_ �_�_Lodo�_�o�o4o �oXojo3�oN�or���o��s�S��B���z�  h��z ��C�:y
 P�v�]�����UD1:\������qR_GRP �1C��� 	 @Cp���$� �H�6�l�Z��|������f���˟���ڕ?�  
���<�*� `�N���r�������ޯ ̯��&��J�8�Z����	�u�����sS�CB 2D� �����(�:�L��^�pς��|V_CONFIG E����@����ϖ�OUT?PUT F�������6�H�Z� l�~ߐߢߴ������� �����#�6�H�Z�l� ~������������ ��2�D�V�h�z��� ������������
� .@Rdv��� ����)< N`r����� ��//%8/J/\/ n/�/�/�/�/�/�/�/ �/?!/4?F?X?j?|? �?�?�?�?�?�?�?O O/?BOTOfOxO�O�O �O�O�O�O�O__+O >_P_b_t_�_�_�_�_ �_�_�_oo'_:oLo ^opo�o�o�o�o�o�o �o $����!�b t������� ��(�:�-o^�p��� ������ʏ܏� �� $�6�G�Z�l�~����� ��Ɵ؟���� �2� D�U�h�z�������¯ ԯ���
��.�@�Q� d�v���������п� ����*�<�M�`�r� �ϖϨϺ�������� �&�8�J�[�n߀ߒ� �߶����������"� 4�F�W�j�|���� ����������0�B� S�f�x����������� ����,>Pa� t��������(:L/x���k}gV� K���//&/8/ J/\/n/�/�/�/W�/ �/�/�/?"?4?F?X? j?|?�?�?�?�/�?�? �?OO0OBOTOfOxO �O�O�O�?�O�O�O_ _,_>_P_b_t_�_�_ �_�O�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����o� ��� �2�D�V�h� z��������ԏ��� 
��.�@�R�d�v��� ������Ϗ����� *�<�N�`�r������� ��˟ޯ���&�8� J�\�n���������Ż��$TX_SCR�EEN 1G�g�}�ipnl/��gen.htmſ�*��<�N�`ϽPa�nel setupd�}�dϥϷ����������ω�6�H� Z�l�~ߐ�ߴ�+��� ����� �2�߻�h� z������9�g�]� 
��.�@�R�d���� �����������}� ��<N`r�� ;1��&8 �\��������QȾUALRM_MSG ?��� �Ȫ-/?/ p/c/�/�/�/�/�/�/��/??6?)?Z?%S�EV  -��6"ECFG �I��  �ȥ@�  A�1 �  B�Ȥ
  [?ϣ��?OO%O7O IO[OmOO�O�O�G�1�GRP 2J�;; 0Ȧ	 �?�O� I_BBL_N�OTE K�:T��lϢ��ѡ�0RDEF�PRO %+ (%N?u_Ѡc_�_�_ �_�_�_�_o�_o>o�)oboMo�o\INU?SER  R]�O��oI_MENHI�ST 1L�9  �(�` ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1�oCUgy�)
13/������p	�vedit(rTG1�I�[�m���� �*pZERO`8�Ώ���� �|o *�<�N�`�r������ ��̟ޟ����&�8� J�\�n����!���ȯ گ����3T�`q�� B�T�f�x��������� ҿ����ϩ�>�P� b�tφϘ�'�9����� ����(߷�L�^�p� �ߔߦ�5������� � �$����Z�l�~�� ���C�������� � 2��/�h�z������� ��������
.@ ��dv����� _�*<N� r�����[� //&/8/J/\/��/ �/�/�/�/�/i/�/? "?4?F?X?C�U��?�? �?�?�?�?�/OO0O BOTOfO�?�O�O�O�O �O�O�O�O_,_>_P_ b_t__�_�_�_�_�_ �_�_o(o:oLo^opo �oo�o�o�o�o�o  �o$6HZl~i? {?������ 2�D�V�h�z����-� ԏ���
����@� R�d�v�����)���П ���������N�`� r�������7�̯ޯ� ��&���J�\�n�����������$UI�_PANEDAT�A 1N����ڱ  	��}  frh�/cgtp/wi�dedev.st�m���%�7�I�Y�)  riρ�@�� �ϫϽ�������Z�� )��M�4�q߃�jߧ� �����������%�7���[�7�� � �   	 
JL�Ϙ����� ����E����:�L�^� p�������������� ��$H/l~ e������o�ܳ7�<N`r ����-���/ /&/8/�\/n/U/�/ y/�/�/�/�/�/?�/ 4?F?-?j?Q?�?�? %�?�?�?OO0O�? TO�xO�O�O�O�O�O �OKO_�O,__P_b_ I_�_m_�_�_�_�_�_ oo�_:o�?�?po�o �o�o�o�oo�o sO $6HZl~�o� ������ �2� �V�=�z���s����� ԏGoYo�.�@�R� d�v�ɏ����П� �����<�N�5�r� Y�������̯���ׯ �&��J�1�n���� ���ȿڿ����c� 4ϧ�X�j�|ώϠϲ� ��+��������0�B� )�f�Mߊߜ߃��ߧ� ��������P�b� t����������S� ��(�:�L�^���� i�����������  ��6ZlS�w�'�9�}���"4FX)�}�� l�����/j '//K/2/D/�/h/�/ �/�/�/�/�/�/#?5?�?Y?��C�=��$U�I_POSTYP�E  C�?� 	 e?�?��2QUICKME/N  �;�?�?��0RESTORE� 1OC�?  �L?��!6OCC1O��maO�O �O�O�O�OuO�O__ ,_>_�Ob_t_�_�_�_ UO�_�_�_M_o(o:o Lo^oo�o�o�o�o�o �oo $6H�_ Ugy�o���� �� �2�D�V�h�� ������ԏ��� �w�)�R�d�v����� =���П������*� <�N�`�r������� �ޯ���&�ɯJ� \�n�������G�ȿڿ������7SCRE��0?�=uw1sc+@u2K�U3K�4K�5K�6K��7K�8K��2USE�R-�2�D�T,�M�k�sUô�4��5��6ʴ�7��8���0ND�O_CFG P�;� ��0PDAT�E ����None�2��_I�NFO 1QC�@��10%�[���I� ��m߮��ߣ������� ���>�P�3�t��i�����<-�OFFSE/T T�=�ﲳ $@������1�^�U� g�������������� ��$-ZQcu����?�
����U�FRAME  ���*�RTOL_ABRT	(�!�ENB*GRP� 1UI�1Cz  A��~��~ ���������0UJ�9MS�K  M@�;N%8�%��/�2oVCCM��V��V�#RG�#Y�9����/����D�BH��p71C����3711?�C0�$MRf2_�*S�Ҵ��	���~XC�56 *�?�6����1$�5���A�@3C��. ��8�?��OOKOx1FOsO�5�51���_O�O�� B����A2�DWO�O 7O_�O8_#_\_G_�_ k_}_�__�_�_�_�_�"o�OFoXo�%TCC��#`mI1�i������� GFS��2�aZ; �| 23�45678901 �o�b�����o�� !5a�4BwB�`56� 311:�o=L�Br5v1�1~1�2�� }/��o�a��#� GYk}�p��� ����ُ�1�C�U� 6�H���5�~���ߏ����	���4�dSEL#EC)M!v1b3��VIRTSYNC��� ���%�SI?ONTMOU�������F��#bU��U�(u FR:\H��\�A\�� �߀ MC��LO�G��   UD�1��EX����'� B@ �����̡m��̡  O�BCL�1�H� ��  =	 �1- n6  G-������[�,S�<A�`=��͗���ˢ��TRAIAN⯞b�a1l�
0�d�$j�T2cZ; (aE2ϖ�i��;� )�_�M�g�qσϕϧπ�������	��F�S?TAT dm~2!@�zߌ�*j$i߾߮�_GE�#eZ;��`0�
� 02���HOMIN� f�U��U� P~�����БC�g�X����JMPERR {2gZ;
  �� *jl�V�7�������� ������
��2�@�q�hd�v�B�_ߠRE� �hWޠ$LEX��i�Z;�a1-e��VM�PHASE  �5��c&��!OFFX/�F�P2n�j�0�㜳E1@���0ϒE1!1?s33�����ak/�k�xk䜣!W�m[�� ���[����o3;� [i {����/ �O�?/M/_/q/� �/��//�/'/9/�/ =?7?I?s?�/�?�/�/ �?�??Om?O%O3O EO�?�?�O�?�O�O�? �O�O�O__gO\_�O E_�O�_�O�O/_�_�_ �_oQ_Fou_�_|o�o �_�oo�o�o�o�o;o Mo?qof-�oI� ����7�[ P���������ˏ ��!�3�(�:�i�[��ŏg�}������TD�_FILTEW�n��� �ֲ:��� @���+�=�O�a�s� ��������֯��� ��0�B�T�f�x����SHIFTMENoU 1o[�<��%��ֿ����ڿ�� ��I� �2��V�hώ� �Ϟϰ�������3�
��	LIVE/S�NAP'�vsf�liv��E��^��ION * Ub�h�menu~߃��`���ߣ���p����	����E�.�5T0�s�P�@� ���AɠB8z�z���}��x�~�P��c ���MEbЩ��<�0���M�O��q���z�W�AITDINEN�D������OK�1�OUT���S�D��TIM����o�G���#���C����b������REL�EASE������T�M�������_A�CT[�����_D?ATA r���%L����xRDI�Sb�E�$XV�R�s���$ZA�BC_GRP 1Ut�Q�,#�0�2���ZIP�u�'�&����[M�PCF_G 1v��Q�0�/� wx�ɤ� 	�>Z/  85�/0�/H/�/l$?��+�/ �/�/?�/�/???r?>�?  �D0�? �?�?�?�?�;����x�]hYLINuD֑y� ��� ,(  *VO�gM.�SO�OwO�O�M i?�O�O^PO1_�O U_<_N_�_�O�_�_�_ _�_�_x_-ooQo8o`�_�o�oY&#2z�� ���oC�e?�a?>N|�oq�����qA�$DSPHE_RE 2{6M��_ �;o���!�io| W�i��_��,��Ï�� �Ώ@��/�v���e� ؏��p���������l�ZZ�� �N