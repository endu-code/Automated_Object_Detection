��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA!R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B!SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C?CFS_UT~p0 "�1�3�#�ؗ`qX"�}R0  4F OIMCM�`O#S�` ��upi �_�p��BA"���M/� h�pIMPEE_F�N��N���@O��r�D_�~�n��Dy�F� dCC_8�r0  T� '��'�DI�n0"���p�P�$I�������F�t �X� GRP0��M=qNFLI�7��0UIRE��$g"� �SWITCH5�A�X_N�PSs"CF�_LIM� w� �0EED��@!��qP�t�`PJ_d=VЦMODEh�.�Z`�PӺ�ELBOF� ������p�  ���3���� FB/���0�>�G� }�� WARNM�`�/��qP��n�NS]T� COR-0b�FLTRh�TRA�T�PT1�� $A�CC1a��N ��r�$ORI�o"V�R�T�P_S� CHUG�0I��rT2��1�I��T�I1�|�� x i#��Q��HDRBJ�; CQ�2L�3L�4*L�5L�6L�7L� �N�9s!��O`S <F +�=�O��#�92��LLECy�>"MULTI�b�"�N��1�!���0T�� ;�STY�"�R`�=l�)2`����*�`T  |� �&$��۱m��P�̱�U�TO���E��EX�T����ÁB���"�2� (䈴![0�������<�b+�� "D"���ŽQ��<� ��kc��'�9�#��與1��ÂM�ԽP��"� '�3�$ L@� E���P<��`A�$JOBn�T���l��TRIG3�% d K�������<���\��+�Y�p�_M��7& t�pFLܐBsNG AgTBA�  ���M��
�!��p� �q��0�P[`��O�'[���0tnah*���"J��_R��CDJ��IdJ
k�D�%C�`�Z����0��P_�P��@ ( @F RO.��&��t�IT�c�NOM��
����S6�CP`T)w@���Z�1P�d���RA�0��p2b"����
$T��.��MD3�T��`QU31���p(5!HGb��T1�*E�7��c�KAb�WAb�cA4#Y�NT���PDBG�D�� *(��PU�t@X��W���AX���a��eTAI^cB�UF��0!+ g� 7n�PIW��*5 P�7M�8M�9
0�6F�7SIMsQS@>KEE�3PATn�^�a" 2`#��"�L64FIX!, ���!d��D�12Bus=CCI�:FgPCH�P:BAD렀aHCEhAOGhA]HW�_�0>�0_h@�f�Ak� ��F�q\'M`#�"�:DE3�- l�p3G@��@FSOES]FgH�BSU�IBS9WC��.� ` ��MARqG쀳��FACLp�SLEWxQ�e�ӿ��MC��/�\pSM_JB M����QYC	g�e�q��Q�0 ā�C�HN-�MP�$G� Jg�_� #���1_FP$�!TC uf!õ#�����d�#a���V&��r�a;�fJ�R���rSEGFR�PIO� STReT��N��cPV5���!41�r��
r>�İ�b�B�O�2` +�[���,qE` &�,q`y�Ԣ}t��yaSIZ%���t�v�T�s� �z�y,qRSINF}Oбc���k ��`��`�`L�ĸ �T`7�CRCf�ԣCC/�9��`a�uah�ub'�MIN��uaDs�T#�G�D�YC��C������e�q0��� �E�V�q�F�_�eF��N3�s�ah��Xa+ep,5!�#1�!OVSCA?� A��rs1�"!3 ��` F/k��_�U��g��]���C�� a�s���R�4� ����N�����5a�R�HANC���$LG��P�f1�$+@NDP�t�AR5@N^��a�q���c���ME�18���}0��RAө�AZ 𨵰:�%O��FCTK���s`"�S�PFADIJ�OJ�ʠ�ʠ�@��<���Ր��GI�p�BMP�d�p�Dba��AES�@	�K�;W_��BAS�� оG�5  M�I�T�CSX[@@�!m62�	$X���)T9�{sC��N�`�a~~P_HEIGHs1�;�WID�0�aVTF ACϰ�1A�P8l�<���EXPg����|��CU�0MME�NU��7�TIT,AE�%)�a28��a��8 P� a��ED�E� ��PD�T��REM.��A�UTH_KEY � ������ �b�Ox	�!}1ERRLH�� �9 \� �q-�O9R�DB�_ID�@l ��PUN_O��Y�$SYS0��4g�-�5I�E�EV�#q�'�PXWO�� �:� $SK7!f2�&�Td�TRL��; �'AC�`��Ġ7IND9DJ.D���_��f1��f���P5L�A�RWAj��"�SD�A��!+r|>��UMMY9d�F�C10d�&���J�<��v}1PR� 
3��POS��J�= l�$V$�q
�PL~�>���SܠK�)?����CJ�@�����ENE�@T��A����S_�RECOR���BH 5 O��@=$LA�>$ ~�r2�R��`�q�b`�3_Du��0RO�@�aT[�Q��b������x! }У�PAUS��>�dETURN���MRU�  CR�p�EWM�b�AGNsAL:s2$LA��!?$PX�g@$P�y A ��Ax�C0 #ܠDO��`X�k�W�v�q�GO�_AWAY��MO��ae���]�CSS�_CCSCB C� �'N��CERI@��гJ`u�QA0�}��@�GAG� R�0�`��{`��{`OF�q�5���#MA��X���&шLL�D� �$���sU�D�)E%!`���OVR310W�,�OR|�'�?$ESC_$`�eDSBIOQ��l q��B�VIB&� �c,�����f�=p�SSW���f!VL���PL���ARMLO
��`����df7%SC �bALspH�MPCh �Ch P�#h �#h 5�UU� ��C�'�C�'�#�$'�d�#C\4�$�pH���Ou��!Y��!�SB ���`k$4�C�P3�Wұ46$VOL�T37$$`�*��^1��$`O1*�$,o��0RQY��2b4~�0DH_THE�����0SЯ4�7ALPAH�4�`���7�@ �0T�qb7�rR�5�8 8� ×���"��JFn�MӁVHBPFUAFLQ"D�s�`�THR��i2dBP�����G(��PVP������������1�J2`�B�E�C�E�CPSu� Y@��Fb3���H�(V �H:U�G�
X0��FkQw�[�Na�'B���C �INHBcFILT���$��W�2�T 1�[ ��$����H YАAF�sDO ��Y�Rp� fg�Q� +�c5h�Q�iSh�Q�PL���Wqi�QTMOU�#c�i�Q\��X@�gmb��vi�h�bAi�fI�aHIG��caB	xO��ܰ��W�"v�AN-u!��	#AVj�H!Pa8$P�(ד#p�R_:�A�a���B�N0�X�M�CN���f1[1�qVAE�p��Z2;&f�I�Q�O�u�rx�wGldDEN{G|d��aF>�!�9��aM:�U�FW	A�:�Ml���X�Lu���$!����!l�ZO ����0%O�lF�s�1&3�DI�W�@���Q���_��!CUgRVA԰0rCR41ͰZ�C<�r�H�v����<�`��<�(�f�CH �QR3�S���t���Xp�VS_�`�ד�IF��ژ�������NSTCY_ OE L����1�tP�1��U��24�2B��NI O7������DwEVI|� F���$5�RBTxS�PIB�P���BY�X����T��HN�DG��G H tn���L��Q��C���5��Lo0 aH��閻�FBP�{tFE{�5�t��T���I�DO���uPMCS�v>�f>�t�>"HOTSW�`s��ІELE��J T���e�2��25�� O� ��HA7�E��3�44�0?��A�K ݬ� MDL� 2J~PE��	A��s ��tːÈ�s�JÆG! ��rD"�ó�����\�TO��W�	��/���SLAV�L  �0INPڐ���`�%ن_CFd�M�� $��ENU��OG��b�ϑ]զPƟ0`ҕ�]�ID�MA�Sa��\�WR0�#��"]�VE�$a�SKI�STs��sk$��2u���J��������	��Q���_SV>h�EXCLUMqJ2NM!ONL��D�Y���|�PE ղI_V>�APPLYZP���HID-@Y�r�_Mz�2��VRFY�0���r�1�cIOC_�f�� 1������O̥�u�LS���R$�DUMMY3�!����S� L_TP�/Bv�"���AӞ�ّ �N ���RTy_u�� չG&r[�O D��Pw_BA�`�3&x�!F ��_5����H������ �� �P $�KwARG�I��� q�2O ���SGNZ�Q q�~P/�/PIGNs�l�$�^ sQ>ANNUN�@�T`<�U/�ߴ�LAzp`]	Z�d~����EFwPI�@ Rk @�F?IT�?	$TOTA%��Pd���!�M�NIY�S+���E��A[�
DAYS\�ADx�@��	�� �EFF_AX�I?�TI��0zCO�JA �ADJ_�RTRQ��Up���<P�1D �r5̀Ll�T�0? ]P�"�p��mtpd��V �0w�G���������SK�SU� ��CTRL_CA��� W�TRAN�S�6PIDLE_�PW���!��A�V曧V_�l�V ��DIAGS���X�� /$2�_SE�#TAC���t!`�!0z*@��RR��vPA���p ; SW�!�!�  ��ol��U��oOH��P�P� ��IR�r��BcRK'#��"A_Ak� ��x 2x�9ϐZs2��%l�W�0t*�x%oRQDW�%MSx��t5AX�'�"��LI�FECAL���10��N�1{"�5Z�3�{"dp5�ZU`}�MO�TN°Y$@FL9A�cZOVC@p�5�HE	��SUPP!OQ�ݑAq� Lj (CL�1_X6�IEYRJZRJWRJ�0TH�!UC|��6�XZ_AR�p6��Y2�HCOQ��MSf6AN��w$��ICTE�Y `>��CACHE�Cp9�M�PLAN��oUFFIQ@�� �0<�1	��6
�N�wMSW�EZ 8䐟KEYIM�p��TM~�SwQq�wQ#�|���OCVIE� ��[ A�BGL���/�}�?����D�?��D\p�ذST��!�R� �T� �T�� �T	��PEMAI�f�ҁ��_FAKUL�]�Rц�1��U�КR�DTR�E�^< �$Rc�uS�% IT��BUFW}�W��9N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTT(����sP��M��Ot�T�LwAX � ��XX~`9#�c_G�3
ЧYN_1�_�D���1 �2M�*��T�F��H@ ~g�`� 0p���Gb-sC_R�AIAK���r�t�RoQ8�u7h�qDSPq��rP��A�IM�c6�\����s2�U�@�A�s�M*`IP���s�!DҐ6�TH�@n�)�OyT�!6�HSDI3��ABSC���@ V`y��� �_D�/CONVI�G��H�@3�~`F�!�pd��psqSCZ"���sgMERk��qFB��Lk��pET���aeR�FU:@DUr`����x�CD,���@p;cJHR�A!��bp�ՔՔ+PSԕC���C��p0�ЕSp�cH *�LX�:cd�Rqa� | ����W��U��U�@�U�	�U�OQU�7R��8R�9R��0T�^�1�k�1x�1��1��1���1��1��1ƪ2RԪ2^�k�2x�2��U2��2��2��2��U2ƪ3Ԫ3^�3k�Bx�3���o���3��U3��3ƪ4Ԣ��EXTk!0�d < � 7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr����\䂴2REM� Fj�N�BOVM��A�oTROV�DT�`6-�MX<�IN��0�,�W!INDKЗ
xw�׀�p$DG~q 36��P�5�!D�6��RIV���2�BGE[AR�IO�%K���DN�p��J�82�P|B@�CZ_MCM�@ȴ1��@U��1�f y,②a? ���P\�"?I�E@��Q�]�am���g� j_0Pfqg RI9e�j�k!UP2_ 3h � �cTD�p�〪�! a���TQ�bB;AC�ri T�P�b��`�) OG��%p���p��IFI�!`�pm�>��	�PT�"���MR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4�@��Uk��� �T�FS#p�Tl �P���e�qP�p$GEX_���1M�2��2� 3�5��9G ���m ��Ѝ��SW�eOe6DEBcUG���%GR���pU�#BKU_�O�1'� �@PO��I5�5MSf��OOfswSM���E�b?��0�0_E �n �0�Y.�D�TERM�o�����ORI�+�p�D�SM�_���b�q�E � �TA�r�y�pe�UP�Rs� -�1�2n$|�' o$SEG,*�> ELTO��$wUSE�pNFIA�U"4�e1���#$p$UFR���0ؐO!��0����OT�'�TqAƀU�#NST��PAT��P�"PTHJ����E�P rF�V"ART�``%B`�a�bU!REL:�aS�HFT��V!�!�(_�SH+@M$���� ���@N8r����OV9Rq��rSHI%0���UN� �aAYLO����qIl����!�@��@ERV]��1� ?:�¦'�2��%��5��%�RCq��EAScYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba��
5aPo��0�p6OR��MY� `GR��t 2b5n� � ��UPaN�Uu Ԭ")���TOCO!S�1POP ��`�pC�����e��Oѥ`REP�R3��aO�P�b�"ePR�%WU.X1���e$PWR��IM�IU�2R_	S�$VI1S��#(AUD���D�v" v��$H|���P_ADDR��H�G�"�Q�Q�QБqR~pDp1�w H� SZ�a��e�ex��e��SE��r��H�S��MNvx ���%Ŕ��OL���p<P��-���ACROlP_!QND_C��ג�1�T �OROUPT��B_�VpQ�A1Q�v��c _��i���i��hx��i����i��v�ACk�I	OU��D�gfsu^d��y $|�P_�D��VB`bPRM�_�b��HTT�P_אHaz (��OBJEr��P��[$��LE�#�s>`{ � ��u��AB_x�T~�S|�@�DBGLV���KRL�YHITC�OU�BGY LO: a�TEM��e�0>�+P'�,PSS|�P��JQUERY_F;LA�b�HW��\!�a|`u@�PU�b�PIO��"�]�ӂ�/dԁ=dԁ�� �IWOLN��}����CXa$SLZ�$INPUT_g�$IP#�P��'���SLvpa~��!�\�`W�C-�B�qIO�p�F_ASv���$L ��w �F1G�U�B0m!���0cHY��ڑ���팒wUOPs� `�� ����[�ʔ[�і"�[PP�SIP�<�іI�2����P_MEMBܿ�i`� X��IP�P�b{�_N�`�����R�����bS�P��p$FOCUgSBG�a~�UJ�Ə� �  � o7JsOG�'�DIS[�J7�cx�J8�7�� Im!�)�7_L�AB�!�@�A��A7PHIb�Q�]�D� J7J\���� �_KEYt� {�KՀLMONa=���$XR��ɀ~��WATCH_����3���EL��}Sy�~���s� �Ю!V8�g� �CTR3�쓥��LG�D� ��R��I�
LG_SIZ���J�q IƖ�I�FDT�IH�_�j V�GȴI�F�%SO��� q �Ɩ���v��ƴ�ǂK�S����w�k�N����E��\���'�*�U�s5��@�L>�4�DAUZ�E�A�pՀ�Dp�f�GH��B?�BOO���� C���PITp���� ��REC��OSCRN����D_p<�aMARGf�`���:���T�L���S��s��W�Ԣ�Iԭ�J{GMO�MNCH�c���FN��R�Kx�PRGv�UF��p0��FWD��HL��STP��V��+������RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28��2��Gh�0PO���������M8�Ģ��EX.��TUIv�I��(�4�@�t�x�J0J�~�P��J0��N�a�#ANA��O"�0�VAIA��dCLE�AR�6DCS_H�I"�/c�O�O&�SI��S��IGN_�vpq�uᛀ�T�d� DEV-�L1LA �°BUW`Ո�x0T<$U�EM��Ł���q��A�R��x0�σ\�a�@OS1�2��3�a�`� �ࠜh�AN%-���-��IDX�DP�2MRO���Գ!�ST��R�q�Y{b! �$E&C+��p.&�A&�p���`� L ��ȟ%Pݘ��T\Q�U�E�`�Ua��_ � �@(��`������# �MB_PN�@ R`r��R�w�TR�IN��P��BAS8S�a	6IRQ6����MC(�� ���CLDP�� ETRQLI��!D�O9=4FLʡh2�Aq3z1D�q7��LDq5[4q5ORG�)�2� 8P�R��4/c�4=b-4�t� �rp[4*�L4
q5S�@TO0Qt�0*D}2FRCLMC@D �?�?RIAt,1ID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCESJ?R�EMhPa�͠��BD4`�B�q`�`�F_A�J�C[��O�H� K��� \ȶ��bTf$� ��LI��q�SREQUIR�E�#MO�\�a�XD�EBU��,1L� M䵔 �p���P�c�AA,1N��
Q�qa�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N�i�PST9� � �4��LOC�RI쀀�EX�fANGx��A,1ODAQ䵍��@$��9�ZMF�����f��"��%8u#ЖVSUP�%�ѻFX�@IGGo�� �rq�"��1��#B��$���p%#by���rx���vbPDAT	AK�pE;����R���M��*� t�`MD�qI��)�v� �tĀA�wH�`��tDIyAE��sANSW�P�th���uD��)�b�ԣ(@$`� PC�U_�V6�ʠ�d�PL�Or�$`�R���B����B�p�����,1R�R2�E�  ���V�A/A d$OCALI�@��G~��2��!V��<$R�SW0^D"���ABC�hD_J2�SE�Q�@�q_J3:M�
G�1SP�,��@PG�n�3m�u�3p
�@��JkC���2'A�O)IMk@{BCS�KP^:ܔ9�wܔJy�{BQܜ������`_AZ.B��?�E�L��YAOCMP0�c|A)��RT�j�ƚ�1�ﰈ��@1�茨����Z��SMG0��pԕ� ER!���#P�INҠACk�p����b�n _�������D��/R��DIU��CD�H�@
�#a�q$�V�Fc�$x��$���`@���b���̂�E�H �$�BELP����!ACCEL���kA°�IRC_R�pG0��T!�$PS�@B2L`���W3��ط9� ٶPAT!H��.�γ.�3���p�A_��_�e�-B�`�C���_MG��$DD��ٰ��$FW�@�p����γ�����DE��PPAB�N�ROTSPE�Eu��O0��D�EF>Q��`$U�SE_��JPQPCD��JY����-A 6qYN�@A�L�̐�nL�MOU�NG���|�OL�y�INC U��a�¢ĻB��ӑ�AENCS���q�B��X���D�IN�I��0���pzC�VE�����23_U ��b�/LOWL���:�O0��0�Di�B�PҠȠ ��PRC����MOS� gTMOpp�@-GPERCH  M�OVӤ �����! 3�yD!e�]�6�<�� ʓA����LIʓdW�ɗ��:p3�.�I�TRKӥ�AY����?Q ^���m�b��`p�CQ�� MOM�B?R�0u��D���y�0Â擰DUҐZ�S_BCKLSH_C�� ��o�n��TӀ���x
c��CLALJ���A��/PKCHKtO0�Su�RTY� B�q��M�1�q_
#Nc�_UMCP�	C�΂�SCL���LMTj�_L�0X����E�� �� ����m�h���6��P	C����H� �P�Ş�CN@�"XT����C�N_��N^C�kCS	F����V6����ϡpj���nCAT�SHs�����ָ1����֙���������PAL���_P���_P0�� e���O1u�$xJaG� P{#�OG�>��TORQU(�p� a�~����Ry������"_W��^�����4t��
5z�
5I;I ;Iz�F�`�!��_8�1���VC��0�D�B�21��>	P�?�B�5JRK��<�2�6i�DBL_�SM�Q&BMD`_D9Lt�&BGRV4
D0t�
Dz��1H_���31�8JCOSEKr�EHLN�0hK�5oDt�jI���jI<1�J�LZ1�5Zc@y��1MYqA�HQB�THWMYTHET=09�NK23z�/Rln�r@CB4VCBn�CqPASfaYR<4gQt�gQ4VSBt��R?U'GTS���Cq��a���P#���Z�C$DUu ��R䂥э2�V�ӑ��Q�r�f$NE��+pIs@�|� �$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b�FP�c�j�FR�VrhVghTd��lV�jV�kV�kUV�kV�kV�kV�iHrh�f�r�m!�x�kUH�kH�kH�kH�kUH�iOclOrhO���nO�jO�kO�kO��kO�kO�kO�FF�.bTQ���E��egSPBALANCE���RLE�PH_'US�P衅F��F��FPFULC�3��3��E��1�l�UTOy_p �%T1T2t���2NW�����ǡ@��5�`�擳�T��OU���� INSE9G��R�REV��R����DIFH��1�l��F�1�;�OB��;C��2� �b�4?LCHWAR��;��ABW!��$ME�CH]Q�@k�q��AXk�P��IgU�i��� 
���!����ROB��CR��ͥ_�� �C��_s"�T � x ?$WEIGHh�9�#$cc�� Ih�.�sIF ќ�LAGK��8SK��K�BIL�?�OD��U��STŰ�P�; ����������
�Ы�Lў�  2�`�"�D�EBU.�L&�n���PMMY9��N8A#δ9�$D&����$��� Q �  �DO_�A��� <	���~��$L�BX�P�N��+��_7�L�t�OH  _�� %��T����ѼT�����TI�CK/�C�T1��%������N��c�Ã�R L�S���S�����_PROMPh�E�? $IR� X�p~ ���!�MAI�0h��j���_9�����t�l�R�0COD捳FU`�+�ID_�" =�����G_SwUFF<0 3�4O����DO��ِ ��R��Ǔن�S����!�{������	�H)�_�FI��9��OR�DX� ����36���X�����GR�9�S��ZDTD�0�t�ŧ4 *�L_NA4���K�>��DEF_I[�K� ��g��_���i��Ɠ��š���IS`i �萚����e����4�0i�Dg����ʍ�D� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{� ��{ԡ�{����}�� v�Ա��g������ ^���K�Փ����!w�N�P'���^����,`�W\�[R����TEFĨ ����OULOMB_tu�0�VISPWITY�A�!OY�A_FRId��(�#SI���R�������3���W�W���0��0_,�EAS%��!�& "����4p�G;� �h ��7ƵCOEFF_Om���$m�/�G!%�S.�߲�CA5����u�GR�` � � �$R� �X]�TM�E�$R�s�Z�/,)�E�R�T;�:䗰� M ]�LL��S�g_SV�($~◰��@���� �"SETU��MEA��Z�x0�u������� � � �� ȰID�"���!*�D�&P���*�F�'����)3��#����"�5;`*��R�EC���!��MS�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I���0�MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X1����MO�R�� H	�CU �A3�z�1Q�
��3���$��FV���2ՠ�AbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų��=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	�����B�s�#�}1� @�@;���O&/�RI#A��
N��xX�s�f�PO_��*�PL}1�,RTv�m��ATUSRBTRC#_T(qR��B ������$ �Ʊ��,�~0�C D��`-CSALl`��SA���]1gqXE@���%���C��J��
���UP(4����P!X��؆�q��3�w�� �PG�5�? $SUB�������t�JMPWAcITO��s��LOyCqFt�!D=�CVF	ш��y���R`�0��CC_CTR�Q�	�IGNR_PLt�/DBTBm�P��z�#BW)����0U@����IG�a��Iy�TNLN��Z�R]aK� !N��B�0�PE�s����r��f�SPD}1� L	�A�`gఠ�S���UN�{���]�R!�BDLY�2������PH_PK��E��2RETRI1Et��2�b���;FI�B� �����8� 2��0DB�GLV�LOGS�IZ$C�KTؑUdy#u�D7�_�_T1@�EM�@C\1A��ℽR��D�FCHE3CKK�R�P�0��e��@&�(bLEc�" PA9�T���P�C�߰PN�����A�Rh�0���Ӯ�PO��BORMATT naF�f1h���2�Sæ�UXy`	��L|B��4�  rE�ITCH��8PL�)�AL_ � �$��XPB�q� C�,2D�!��+2�J3�D��� T�pPD�CKyp��oC� _AgLPH���BEWQo���� ��I�wp� � �b@PA�YLOA��m�_1�t�2t���J3AR���؀դ֏�laTI�A4��5��6,2MOMCP�����������0BϐAD�����\���PUBk`R�Ԑ;���;�����z4�` I$PI\D s�oӓ1yՕ�w�2�w�UZ��I��I��I�〛�p����n���y��e`�9S)bT�SPEED� G��(�Е�� /���Е�`/�e�>���M��ЕSAMP��6V��/���ЕMO�@ 2@�A��QP�� �C��n����������� LRf`kb�ІE9h�EIN09��7S.�В9
yPy�GA�MM%S���D$GGET)bP�cD]Ԛ�2
�IB�q�IN�G$HI(0;A��$LREXPA8)LWVM8z�)��g���C5�C�HKKp]�0�I_��h`eT��n�q���eT,���� ��$�� 1��iPI� RCH_D`�313\��30LE�1��1\�o(Y�7 �t�M�SWFL �M��SCRc�7�@�&��%�n�f�SV���P�B``�'�!�B�sS_�SAV&0ct5B3NO]�C\�C2^�0� mߗ�uٍa��u���u:@e;��1���8��D�P ���������)� �b9��e�GE�3���V�e�Ml�� � �YL��QNQSRlbfqXG�P �RR#dCQp� �S:AW70�B�B[�CdgR:AMxP�KCL�H����W�r�(1n�g�M�!o�� �F�P@}t$WP�u�P r�� P5�R<�RC�R�� %�6�`��� ��qsr %X��OD�qZ�Ug��ڐ>D� ��OM#w�J?\?n?�?�?@��9�b"���]�_��� |��X0��bf ��qf��q`�ڏgzf�ڡEڐ�>j�"�5�t��FdPB��PM��QU�� � 8�L�QCOU!h Q�THI�HOQBpH�YSY�ES��qU�E�`�"�O��� � �P�@\�UN����Cf�O�� P��Vu��!����OOGRAƁcB2�O�tVuITe �q:p/INFO�����{��qcB�e�OI�r�{ (�@SLEQS� �q��p�vgqS����� 4L�ENA�BDRZ�PTION�t�����Q���)�GCuF��G�$J�,q^r�� R����U�g��rS_ED������ �F��PK���E'NU�߇وAUT$1܅COPY�����n�00�MN���PR�UT8R �Nx�OU��$G[rf���_RGADJ���*�3X_:@բ$�����P��W��P��} ���)�}�EX�YCZDR|�NS.��F@�r�LGO�#�NY�Q_FREQR�W`� �#�h�TsLAe#�����ӄ �CRE�� s�IF��sNmA��%a�_Ge#STATUI`e#MAIL�����q �t�������ELE�M�� �/0<�FEASI?�B��n��ڢ�1�]� � I �p��Y!q]�t#A��ABM���E�p<�VΡY�BASR�Z���S�UZ��0$�q���RMS_TR ;�qb ���SY�	�ǡ���$���>C�Q`	~� 2� _ �TM������̲�@ ��A��)ǅ�i$DOUd�s]$Nj���PR+@z3���rGRID�q�M�BARS �TY�@��OTO�p��� Hp_}�!����d��O�P/�� � �p�`POR�s��}�.��SRV��)����DI&0T����� �#�	�#�4!�5!�6J!�7!�8�e�F��2��Ep$VAL�Ut��%��ֱ��/��� ;�1�q��1���(_�AN�#��ⓡRɀ(���TOTcAL��S��PW��Il��REGEN�1�cX��ks(��a����`TR��R��_!S� ��1ଃV�����⹂Z�E��p�q���Vr���V_H��DqA�S����S_Y,1��R4�S� AR�P2�� ^�IG_S!E	s����å_Zp���C_�Ƃ�ENHA�NC�a� T �;�������IN�T�.��@FPsİ_OVRsP�`p�`��Lv��o��7�}���Z�@�SLG�AA�~�25�	��D��YS�BĤDE�U�̦���TE�P���G� !Y��
�J��<$2�IL_MC�x r#_��`TQ�`��q����'�BV�C�P�_� 0�M�	V1V�
V1�2�2�U3�3�4�4�
 �!���� � m�A�2;IN~VIBP����1�2�2�3*�3�4�4�A@p-�C2���p� �MC_Fp+0B�0L	11d���M501Id�%"E� S`�R�/�@KEEP__HNADD!!`$$^�j)C�Q���$��"	��#O�a_$A�!pK��#i��#REM�"��$��½%�!�(U�}�e�$HPWD � `#SBMSUK|)G�qU2:��P	�COLLAB � �!K5�B�� ��g��pITI1{9p#n>D� ,�@FLAP>��$SYN �<�M�`C6���UP�_DLYAA�ErDGELA�0ᐢY�`�AD�Qz�QSKI�P=E� ���XpO�fPNTv�A�0P_ Xp�rG�p�RU@,G�� :I+�:IB1:IG�9JTЀ9Ja�9Jn�9J{�9J9�<��RA=s� AX���4�%1�QB� NFLIC�s�@J��U�H�LwNO_H��0�"?��RITg���@_PA�pG�Q�� �K�^�U��W���LV�d�NGRLT�0_q��O�  " ��OS��T_JvA V	��APPR_WEI{GH�sJ4CH?p�vTOR��vT��LO!O��]�+�tVJ�е��ғA�Q�U�S�XOB�'�'�{�J2P���
7�X�T�<a43DP�=`Ԡ\"<a�q\!��RsDC��L� �рER��R�`� �RV�p�jr�b�RGE��8*��cN�FLG�a�Z����SPC�s�U�M_<`^2TH2�NH��P.a 1�� m`EF11��� lQ �!#� <�p3AT� g�S�&� Vr�p�tMq�Lr���HOMEwr�t2'r�-?Qcu��w3'r���P����w4'r�'�@9�K�]�o����w5'r뤏��ȏڏ����w6'r�!�3�E�W�i�{��w7'r힟��Pԟ����w8'r��@-�?�Q�c�u��uS$0
�q�p�� sF��`ala�!`P����a�`/���-�IO[�M�I֠��*�PO{WE�� ��0Za*��� �5��$DSB G'NAL���0Cp�нlaS2323�� �~`��� / I3CEQP��PEp���5PIT����OPB�x0��FLOW�@T�RvP��!U���CU:�M��UXT�A��>w�ERFAC�� �U��ɲCHN��� tQ  _���>�Q$����OM���A�`T�P#UKPD7 A�ct�T���UEX@�ȟ�U E�FA: X"�1RSP�T�����T ���PPA�0o񩩕`EXP�IOS���)ԭ��_���%��C�WR�A��ѩD�ag֕`Ԧ?FRIENDsaC2�UF7P����TOO�L��MYH C2L�ENGTH_VT�E��I��Ӆ$�SE����UFIN�V_���RG9I�{QITI5B�ױXv��-�G2-�G�17�w�SG�X��_��UQQD=#���AS��d~C�`��q��_ �$$C/�S�`�����S0�0��>��VERSI� ��w�0�5���I��������AAV�M_Y�2 �� 0 � �5��C�O�L@�r� Ȱr�	 ����S0����������������
?�QY�BS���1���� <-������ 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO�jO|O�O�O�OiCC��@XLMT��C��  ��DINp�O�A�Dq�EXE�HiPV_��ATQ�z
��LARMRECOV ��RgLMDG �*�5�OLM_�IF *��`d �O�_�_�_�_j�_'o�9oKo]onm, 
 ��odb��o�o�o�o�^��$� z, A�   2D{�PPINFO u[ �Vw��������`������ �*��&�`�J���n�����DQ����
� �.�@�R�d�v����������a
PPLIC�AT��?�P���`Han�dlingToo�l 
� 
V8.30P/40Cp�ɔ_LI
88�3��ɕ$ME�
F0G�4�-

398�ɘ��%�z�
7D�C3�ɜ
�Non�eɘVr���ɞ@/6d� Vq?_ACTIVU�r�C죴�MODP����C�I��HGAP�ON���OU�P�1*��  i�m����Қ_�����1*�  �@��������Q����Կ�@�
������ ���5��Hʵl�K�HTTHKY_��/�M�S� ����������%�7� ��[�m�ߝߣߵ��� �������!�3��W� i�{���������� ����/���S�e�w� �������������� +�Oas�� �����' �K]o���� ����/#/}/G/ Y/k/�/�/�/�/�/�/ �/�/??y?C?U?g? �?�?�?�?�?�?�?�? 	OOuO?OQOcO�O�O �O�O�O�O�O�O__ q_;_M___}_�_�_�_`�_�_�_kŭ�TOp���
�DO_CLE�AN9��pcNM  !{衮o�o�o��o�o��DSPDgRYRwo��HI��m@�or���� �����&�8�J���MAXݐWdak�H�h�XWd�d���PLUGGW�Xgd���PRC)pB�`"�kaS�Oǂ2^DtSEGF0�K�  �+��o�or�������8���%�LAPOb� x�� �2�D�V�h�z��������¯ԯ�+�T�OTAL����+�U�SENUO�\� �e�A�k­�RGDI_SPMMC.����C6�z�@@Dr\�O�Mpo�:�X�_STRING 1	(��
�M!�S��
��_ITE;M1Ƕ  n�� ����+�=�O�a�s� �ϗϩϻ����������'�9�I/O SIGNAL���Tryout� ModeȵI�npy�Simul�ateḏOu�t��OVER�RLp = 100�˲In cyc�l�̱Prog� Abor��̱~u�Statusʳ�	Heartbe�atƷMH F�aul	��Aler�L�:�L�^�p�����������  ScûSaտ��-�?�Q� c�u������������� ��);M_q��WOR.�û�� ����+= Oas��������//'.PO ����M �6/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�?�?H"DEVP.�0d/ �?O*O<ONO`OrO�O �O�O�O�O�O�O__�&_8_J_\_n_PALT	��Q�o_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o�_GRIm�û9q �_as���� �����'�9�K��]�o�������'�R 	�݁Q����)�;� M�_�q���������˟ ݟ���%�7�I�ˏPREG�^����[� ����ͯ߯���'� 9�K�]�o����������ɿۿ�O��$AR�G_� D ?	����0���  	$�O�	[D�]D���O�e�#�SBN_C�ONFIG 
�0˃���}�CI�I_SAVE  �O�����#�TC�ELLSETUP� 0�%  O�ME_IOO�O�%?MOV_H���ώ��REP��J��U�TOBACK�����FRA;:\o� Q�o����'`��o���{� �� f� o�����*�!�3�`�����f������ ����o�{��&�8�J� \�n������������ ������"4FXj |������\끁  ��_i��_\ATBCKC�TL.TMP 6�.VD GIF PHD_q���N�t#��f�IN�I�P�Օ�c�MESSAG�����|8��ODE_D�����z��O�0�c�P�AUSM!!�0� (73�U/g+(Od/�/x/�/�/ �/�/�/�/???P?�>?t?1�0$: TSK�  @-��T�f�UgPDT��d�0�
&XWZD_ENqB����6STA��0��5"�XIS��U�NT 20Ž�� � 	 ���z��e�ng�-�?���S�o�U@��H����zF�OTo�}Cw�g�^�	���.�O�O�O�O�/_2FMET߀2�CMPTAA��@��$A-�@����@���@����]5���5�(d5��P�5�r�5F*�5�338]SCR�DCFG 1�6/�Ь�Ź�_�_oo(o:oLo��o�Q���_�o�o�o �o�o�o]o�o>P bt���o9�iуGR<@M/�s/N5A�/�	i��v�_ED�1�Y� 
 �%-5�EDT-�'�G?ETDATAU�o��9��?�j�H�o��f�\��A��  ���2�&�!�E���:IB���~�ŏ׏m����3��&۔� �D��ߟJ�����9�ǟ�4���ϯ�(�����]�o�����5 N������(�w��)�;�ѿ_��6ϊ�g� ��(�CϮ���ϝ�+��7��V�3�z�(��@z�����i����8��&���~�]���F����5����9~������]����Y�k�����CR�!ߖ��� W�q���#�5���Y��p~$�NO_DEL���rGE_UNUS�E��tIGALL_OW 1���(*SYST�EM*S	$S?ERV_GR�Vܖ : REG�$8�\� NUM�
���PMUB U�LAYNP\?PMPAL��CYC10#6x $\ULSU0�8:!�Lr��BOXORI�C�UR_��PM�CNV�1�0L�T4DLI�0��	����BN/ `/r/�/�/�/�/�/����pLAL_OUT� �;���qWD_ABOR=f�q�;0ITR_RTN��7�o	;0NONS�0�6 
HCCF�S_UTIL 9#<�5CC_@6Aw 2#; h ?��?�?O#O6]CE_�OPTIOc8�qF@RIA_I�c f5Y@�2�0FF�Q�=2q&}�Ao_LIM�2.�� ��P�]B�T�KX�P
�P�2O��Q��B�r�qF�PQ5T1)TR�H��_:JF_PARAMGP 1�<g^&S�_�_�_�_~�VC�  C�dE�`�o!o`�`U�`�`�Cd��T@ii:a:e>eBa�Gg�C�`� D� kD	�`�w?��2{HE ONFI� �E?�aG_P�1#; ���o�1CUgy�aKoPAUS�1�yC ,����� ����	�C�-�g� Q�w���������я���rO�A�O�H��LLECT_�B�IPV6�EN. QF�n3�NDE>� �G��71234?567890��sB�TR����%
 H�/%)������� W���0�B���f�x��� 㯮���ү+����� s�>�P�b��������� �ο��K��(�:�Г�^�|��B!F� ��I|�IO #��<U%e6�'�9�lK���TR�P2$���(9X�t�Y޼`%��̓ڥH��_MOR֮3&�=��@XB��a��A�$� �H�6�l�~���~S��'�=�r_A?�a�a`D��@K��R�dP��y)F�ha�-�_�'�9�%
�k��G�� ��%Z�%���`�@c.�PDB�+���cpmidbg��	�`C:��@�����p��|N  ��@�9+
���]�­@�s<�^�@ssg�$� �sfl�q��ud1:��:J~��DEF *ۈ���)�c�buf.txt�����_L64FIX ,������l/[ Y/�/}/�/�/�/�/
? �/.?@??d?v?U?�?��?�?�?�?�?,/>#_/E -���<2O�DOVOhOzO�O6&IM���.o�YU>�̱�d�
�IMC��2�/����dU�C��2�0�M�QT:Uw�Cz�  B�i�A����A���Au��gB3�*CG��B<�=w�i�B�.��B���B���5B�$�D?�%B���ezV�C�q�C�v��D���D-lE\D�n`�j��B9"��22o�SD|����� ��U���C�C�����
�xObi�D4,cdv`D��`/�`v`�s]E�D D�`� E4�F*� Ec��FC���u[F���E���fE��fFކ�3FY�F�P�3�Z��@�33 ;��>L���A�w�n,a@��@e�C5Y���a���`A��:w�=�`<#���
���?�ozJRSMO?FST (�,bVIT1��D @3���
д����a��;���bw?����<�M�NTES�T�1O�CR@�4h��>VC5`A�w�DIa+a�aORI`CTP�B�U�C�`4�9��r��:d����q�I?�5��qT_~�PROG ���
�%$/ˏ�t��NU_SER  �U�������KEY_TBOL  ����#a��	�
�� !�"#$%&'()�*+,-./��:�;<=>?@AB�C�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~��������������������������������������������������������������������������������͓���������������������������������耇������������������������LCK�
�����STAT/��s_AUTO_DO ��	�c�INDT_'ENBP���Rpqn��`�T2����STO�r`���XC�� 2�6���8
SO�NY XC-56t�"b����@��F( А�HR50w���>�P�y7b�t�Aff����ֿ� Ŀ���� C�U�0�yϋ�fϯ��π���������-ߜ�T{RL��LETEͦ� ��T_SCR�EEN ��Okcs���U��MMENU 17�� <ܹ��� w���������K� "�4��X�j���� ��������5���k� B�T�z����������� ����.g>P �t����� �Q(:�^p ����/��;/ /$/J/�/Z/l/�/�/ �/�/�/�/�/7?? ? m?D?V?�?z?�?�?�? �?�?!O�?
OWO.O@O�fO�OvO�O�O(y��REG 8�y�����`�M�ߎ�_MA�NUAL�k�DB;CO��RIGY�9��DBG_ERRL&��9�ۉq��_��_�_ ^QNUMSLI�pϡ�pd
��
^QPXWORK 1:���_5oGo�Yoko}oӍDBTB�_N� ;������ADB_�AWAYfS�qG�CP 
�=�p�f_CAL�pR��bbRY��[�
�WX_�P 1<
{y�n�,�%oc��P��h_M��IS�O��k@L��sONT�IMX��
����vy
��2sMOT�NEND�1tRECORD 1B��� ���sG�O�]�K��{�b������ ��V�Ǐ�]����6� H�Z���������#� ؟������2���V� şz��������ԯC� ��g��.�@�R���v� 寚�	���п���c� χ�#ϫ�`�rτϖ� Ϻ�)ϳ�M���&� 8ߧ�\�G�Uߒ�߶� ����I������4�� �p7�n���ߤ�� ��������"���F� 1���|��������[� ����i���BTf����bTOLER7ENC�dB�'r�`�L��^PCSS_�CCSCB 3C$>y�`IP�t}�~ �<�_`r� K�����/�{��5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O`�O�O_�~�LL� D��&qET�c�a� C[C�p�PZP^r_ A� %p� �sp��QGPt[	 A�p�Q�_��[? �_�[oU��p�P�pSB� V�c�(a�PWoio{h+�o�X�o�o�Y��[	r�hLW���N:p����}6ڿ��c��aD�@VB��|��G���+��K� �otGhXGr�So�����eB   =��eͶa>�tYB�� ��pC�p�q�aA"�H �S�Q-��q���ud��v�����AfP ` 0���D^P��pk@�a
�QXT�HQ����a aW>� �a9P��b�e:�L�@^�h�Hc�́PQ�R FQ�PU�z�֟�o\ ^��-�?��c�u���,�zCz�ů�b�2�Щ�RD�����l)*����S̡ 0��]�0�.��@���EQ�p��F�X�ѿU�ҁп�VSȺNS?TCY 1E��]�ڿ��K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}ߏ�����DEVICEw 1F5� MZ �۶a��	� ��?�6�c���	{䰟���_�HNDGD G�5�VP���R�LS 2H�ݠ��/�A�S��e�w����� ZPARAM I�FgHe��RBT 2K��8р<��WPp�C�C��,`¢P¨Z�z��%{�C��2�jMTLU,`"nPB, s���M� }�gT�g��
B��!�bcy�[ 2Dchz�����/��/gT#I{%D��C�` b!��R��A��A,���Bd��A��P��_C4kP�!2��C��$Ɓ�]�ff�A�À��B�
� �| ���/�/�T (��54a5�} %/7/d?/M?_?q?�? �?�?�?�?O�?OO %O7OIO�OmOO�O�O �O�O�O�O�OJ_!_3_ �_�_3�_�_�_�_�_ o�_(ooLo^oЁ=? k_IoS_�o�o�o�o�o �o�o#5G� k}������ �H��1�~�U�g�y� ƏAo�Տ���2�D� /�h�S���go����ԟ ����ϟ���R�)� ;���_�q��������� �ݯ�<��%�7�I� [�m���������}� &��J�5�n�YϒϤ� ���ϣ�ѿ������ F��/�Aߎ�e�w��� �߭���������B�� +�x�O�a����� ������,���%�b�M� ��q����������� ����L#5�Y k}��� �� 61CUg� �������	/ /h/���/w/�/�/�/ �/�/
?�/.?@?I/ [/1/_?q?�?�?�?�? �?�?�?OO%OrOIO [O�OO�O�O�O�O�O &_�O_\_3_E_W_�_ ?�_�_�_�_�_"oo Fo1ojoE?s_�_�om_ �o�o�o�o�o0 f=Oa���� ������b�9� K���o���Ώ��[o� �(��L�7�I���m�������$DCSS�_SLAVE �L���ё���_4D � љ��CFG7 Mѕ��������FRA�:\ĐL-�%04�d.CSV��  m}�� ���A i�+CHq�z�������|�����  ������Ρޯ̩ˡҐ-��*����_CRC_OUT N�������_FSI� ?њ ����k�}������� ſ׿ �����H�C� U�gϐϋϝϯ����� ���� ��-�?�h�c� u߇߽߰߫������� ��@�;�M�_��� ������������� %�7�`�[�m������ ����������83 EW�{���� ��/XS ew������ �/0/+/=/O/x/s/ �/�/�/�/�/�/?? ?'?P?K?]?o?�?�? �?�?�?�?�?�?(O#O 5OGOpOkO}O�O�O�O �O�O _�O__H_C_ U_g_�_�_�_�_�_�_ �_�_ oo-o?ohoco uo�o�o�o�o�o�o�o @;M_�� �������� %�7�`�[�m������ ��Ǐ������8�3� E�W���{�����ȟß ՟����/�X�S� e�w����������� ���0�+�=�O�x�s� ��������Ϳ߿�� �'�P�K�]�oϘϓ� �Ϸ���������(�#� 5�G�p�k�}ߏ߸߳� ���� �����H�C� U�g��������� ���� ��-�?�h�c� u��������������� @;M_�� ������ %7`[m�� �����/8/3/ E/W/�/{/�/�/�/�/ �/�/???/?X?S? e?w?�?�?�?�?�?�? �?O0O+O=OOOxOsO��O�O�O�O�C�$D�CS_C_FSO ?����A� P �O�O_?_:_L_^_ �_�_�_�_�_�_�_�_ oo$o6o_oZolo~o �o�o�o�o�o�o�o 72DVz�� �����
��.� W�R�d�v��������� ����/�*�<�N� w�r���������̟ޟ ���&�O�J�\�n� ��������߯گ��� '�"�4�F�o�j�|��� ����Ŀֿ�������G�B�T��OC_RPI�N_jϳ����� ���O����1�Z�U��NSL��@&�h߱��� ������"��/�A�j� e�w��������� ����B�=�O�a��� �������������� '9b]o�� ������: 5GY�}��� ���///1/Z/ U/g/y/�/�/�/�/�/ �/�/	?2?-???Q?z? u?��ߤ߆?�?�?�? OO@O;OMO_O�O�O �O�O�O�O�O�O__ %_7_`_[_m__�_�_ �_�_�_�_�_o8o3o EoWo�o{o�o�o�o�o �o�o/XS ew������ ��0�+�=�O�x�s� ��������͏ߏ�� �'�P�K�]�o������ �PRE_CHKg P۪�A ��?,8�2�<�� 	 8�9�K���+�q���a��� ����ݯ�ͯ�%�� I�[�9����o���ǿ ��׿���)�3�E�� i�{�YϟϱϏ����� ������-�S�1�c� ��g�y߿��߯���� !�+�=���a�s�Q�� ������������ �K�]�;�����q��� ����������#5� Ak{��� ���CU3 y�i����� �/-/G/c/u/S/ �/�/�/�/�/�/?? �/;?M?+?q?�?a?�? �?�?�?�?�?�?%O?/ Q/[OmOO�O�O�O�O �O�O�O_�O3_E_#_ U_{_Y_�_�_�_�_�_ �_�_o/ooSoeoGO �o�o=o�o�o�o�o �o=-s�c �������'� �K�]�woi���5��� ɏ��������5�G� %�k�}�[�������ן �ǟ����C�U�o� A�����{���ӯ���� 	��-�?��c�u�S� ������Ͽ῿��� ��'�M�+�=σϕ�w� ����m������%�7� �[�m�K�}ߣ߁߳� �߷����!���E�W� 5�{��ϱ���e��� ����	�/��?�e�C� U������������� ��=O-s��� ��]����' 9]oM��� ����/�5/G/ %/k/}/[/�/�/��/ �/�/�/?1??U?g? E?�?�?{?�?�?�?�? 	O�?O?OOOOuOSO eO�O�O�/�O�O�O_ )__M___=_�_�_s_ �_�_�_�_o�_�_7o Io'omoo]o�o�o�O �o�o�o!�o1W 5g�k}��� ���/�A��e�w� U�������я��o� ���	�O�a�?����� u���͟�����'� 9��]�o�M������� ��ۯ��ǯ�#�ůG� Y�7�}���m���ſ�� ���ٿ�1��A�g� E�wϝ�{ύ������� 	�߽�?�Q�/�u߇� e߽߫ߛ�������� )���_�q�O��� �����������7� I���Y��]������� ��������!3W iG��}��� �%�A�1w �g������ /+/	/O/a/?/�/�/ u/�/�/�/�/?�/ 9?K?�/o?�?_?�?�? �?�?�?�?O#OOGO YO7OiO�OmO�O�O�O �O�O_�O1_C_%?g_ y__�_�_�_�_�_�_ �_o�_+oQo/oAo�o �owo�o�o�o�o�o );U__q�� ������%�� I�[�9����o���Ǐ �����ۏ!�3�M?� i��Y�������՟� ş����A�S�1�w� ��g����������ӯ��+�=��$DCS_SGN QK��c��7m� �16-MAY-�19 09:20�   O�l�4-J{ANt�8:38}������ N.DѤ���������h��x,rWf*�o��^M��  O��VERSION �[�V3.�5.13�EFLOGIC 1RK���  	���P�?�P�N��!�PROG_EN/B  ��6Ù��o�ULSE  �TŇ�!�_ACC�LIM�����Ö��WRSTJ�NT��c��K�E�MOx̘��� ���I?NIT S.�G��Z���OPT_SL� ?	,��
 ?	R575��YЫ74^�6_�7_�50��1��2_�@ȭ�|�<�TO  H�跿��V�DEXҚ�dc����PA�TH A[�A�\�g�y��HCP�_CLNTID y?��6� @�������IAG_G�RP 2XK� ,`� ��� �9�$�]�H������1234567890����S�� |�������!�� ��H���@;�dC�S���6 �����.� Rv�f��H ��//�</N/� "/p/�/t/�/�/V/h/ �/?&??J?\?�/l? B?�?�?�?�?�?v?O �?4OFO$OjO|OOE� �Oy��O�O_�O2_���_T_y_d_�_,
�B^ 4�_�_~_`O o�O&oLo^oI��Tjo �o.o�o�o�o�o �O '�_K6H�l� ������#�� G�2�k�V���B]��� Ǐُ�������(���L�B\Drx�@���PC����4�  79֐�$��>���:�����ߟ�ʟܟ���CT_C�ONFIG Y���Ӛ�e�gU���STBF_TTS��
��b����Û�u�O�MAU���|��MSW_CuF6�Z��  伿OCVIEW��[ɭ������-� ?�Q�c�u�G�	����� ¿Կ������.�@� R�d�v�ϚϬϾ��� ����ߕ�*�<�N�`� r߄�ߨߺ������� ��&�8�J�\�n�� ��!����������� ��4�F�X�j�|����KRC£\�e��!*� B^������C2�g{�SBL_FA?ULT ]��ި>�GPMSKk���*�TDIAG �^:�աI���UD1: 6789012345�G�BSP�-?Q cu��������//)/;/M/� �
@q��/$��TRECP��

 ��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOi/{/�xO�/UMP_OP�TIONk���AT�R¢l��	�EPM�Ej��OY_TEM�P  È�33B�J�P�AP�D�UNI��m�Q��Y�N_BRK _�ɩ�EMGDI_�STA"U�aQSUN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 J�#!�,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;��A����O ���� � I ߵ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$
T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����裆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7����; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  C��0����(7�?�<B�?B����2�ٸ*9�N SMTT#t�[)��X�4�$HO�STCd1ux����?�� MC�x��;zOx��  27.0�@1�O  e�O�O	_ _-_;Z�O^_p_�_�_��LN_HS	anonymous�_�_�_�oo1o yO��Fh Fk�O�_�o�O�o�o�o �oJ_'9K]�o �_�����4o �XojoG�~�o^��� ����ŏ����� 1�T���y������� ����,�>�@�-�t� Q�c�u���������ϯ ���(�^��M�_� q�����ܟ� �ݿ� �H�%�7�I�[Ϣ�� �ϣϵ����l�2�� !�3�E�Wߞ���¿Կ ����
�������/� v�S�e�w������ �������+�r߄� ��s�����߻����� �����'9K]�� �������4� F�X�j�l>��}� �����// 1/T��y/�/�/�/��/.D\AENT 1=v
; P!J/?  ��/3?"? W??{?>?�?b?�?�? �?�?�?O�?AOOeO (O�OLO^O�O�O�O�O _�O+_�O _a_$_�_ H_�_l_�_�_�_o�_ 'o�_Koooo2o{oVo �o�o�o�o�o�o5 �oY.�R�v���zQUICCA0���3��t14��"����t2��`�r��ӏ!ROUTE�Rԏ��#�!P�CJOG$���!�192.168�.0.10��sC�AMPRTt�P�!�d�1m�����RT�폟�����$NAM�E !�*!R�OBO���S_C�FG 1u�) ��Aut�o-starte�dFTP& ��=?/֯s���� 0�B��f�x������� ��S������,�� �������ϼ�ޯ���� �����ʿ'�9�K�]� oߒ�ߥ߷�������8��SM%y� {�U�ό������� ����
��.�@�c����v������������z �%�7�I�K�8�\ n���k���� �3�FXj|�����a��7 /M*/</N/`/ r/9�/�/�/�/��/ �/?&?8?J?\?�m? ���?�//�?�?O "O4O�/XOjO|O�O�O �?EO�O�O�O__0_ w?�?�?�?�O�_�?�_ �_�_�_o�O,o>oPo boto�_o�o�o�o�o �oK_]_o_L�o�_ �o�����o� � �$�6�Y�Y�~���𢏴�ƏZ�_ERR� w3�я�PDUSIZ  g��^�p���>�W�RD ?r�Cq��  guestb�Q�c�u��������`�SCDMN�GRP 2xr�;���H�g��\�b�K� 	P01.00 8`��   � ��   B  ���� ���_H���L��L�}�L�����O8�`����l�����a4�U  �Ȥ� �8����\���)�`�;��������d�.�@�R�ɛ_GWROUېy������	ӑ���QU�PD  ?u�����İTYg�����TTP_AUT�H 1z�� <�!iPenda�n��-�l���!�KAREL:*8-�6�H�KC]�m���U�VISION SET���ϴ�!�����R�0�� H�Bߏ�f�x��ߜ߮����CTRL {�����g�
��?FFF9E3��At�FRS:DEF�AULT;�F�ANUC Web Server;� )����9�K��ܭ����������߄WR_�CONFIG �|ߛ ;��I�DL_CPU_P5CZ�g�B�I�y�w BH_�MINj��)�}�GNR_IO���g���a�NPT?_SIM_D_������STAL_S�CRN�� ���T�PMODNTOL8������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMAST�E��ɾeSLAV�E ~��c�O�_CFGٱBU�O�O@CYCL�En>T�_ASG� 1ߗ+�
  ����//+/=/ O/a/s/�/�/�/�/���NUM��
�@IPCH�^R?TRY_CNZ��@�@��������1 @kI�+E��z?E�a�P_MEMBERS 2�ߙ�� $���2����ݰ7�?�9a�SDT�_ISOLC  �����$J23�_DSM+�3J?OBPROCN���JOG��1�+��d8�?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSRE�QO��KANJI_����a[�MONG ����b�yN_ goyo�o�o�o�Y�`3	�<� ��e�_ִ���_L���"?`EY�LOGGINL�E�������$L�ANGUAGE Y��<T� {q��LGa2�	�b����g�xP��  *��g�'��b����>�MC:�\RSCH\00�\<�XpN_DISP �+G�H��O��O߃LOCp�D�z���AsOGB?OOK ����`��󑧱����X� ����Ϗ����a�*��	p������!�m��!���=p_B�UFF 1�p��2F幟���՟�D� Collaborativǖ ���F�=�O�a�s��� ����֯ͯ߯����B�9�K���DCS ��z� =��� '�f��?ɿۿ���H@�{�IO 1��# ~?9Ø��9�I� [�mρϑϣϵ����� �����!�3�E�Y�i� {ߍߡ߱��������-E��TMNd�_B� T�f�x�������� ������,�>�P�b��t�������L��SE�VD0��TYPN1�$6���Q�RS"0&��<2FLg 1�"�J0��� �����G�TP:pOF�NGNAM1D�mr�t7UPS�GI"5�a�O5�_LOAD�N@G %�%�TI�pZUZAU�N#�(MAXUALRM�'���(��'_PR"4F0d��1��B_PNP� V� 2�C	M�DR0771ߕz�BL"8063%�@ �_#?�ߒ|/�C��z�6��/􈃟/Po@P 2���+ �ɖ	~T 	t  ��/ �%W?B?{?�k?�? g?�?�?�?O�?*OO NO`OCO�OoO�O�O�O �O�O_�O&_8__\_ G_�_�_u_�_�_�_�_ �_o�_4ooXojoMo �oyo�o�o�o�o�o �o0B%fQ�u �������� >�)�b�M�����{��� �����Տ��:�%��^�p�S�������D�_LDXDISA�pB�MEMO_{APjE ?C
 �,�(�:��L�^�p������� ;1�C ���� 4�������4��X����C_MSTR ����w�SCD 1���L�ƿH�� տ���2��/�h�S� ��wϰϛ��Ͽ���
� ��.��R�=�v�aߚ� �ߗ��߻������� <�'�L�r�]���� �����������8�#� \�G���k��������� ������"F1j Ug������ �B-fQ��u���h�MKCFG ����/�#�LTARM_��
7"0�0N/|V$� METPUᐶ�3����ND� A�DCOLp%A {.C7MNT�/ �%� ����.E#>!�/|4�%POSCF�'=�.PRPM�/9�ST� 1��� {4@��<#�
1 �5�?�7{?�?�?�? �?�?�?)OOO_OAO SO�OwO�O�O�O�O_��A�!SING_C�HK  �/$M/ODAQ,#�����.;UDEV 	���	MC:o\HOSIZEᝢ��;UTASK %���%$123456�789 �_�U9WT�RIG 1���l3%%��9o��"ocoFo�5#�VYP�QNe���:SEM_INF �1�3' �`)AT&F�V0E0po�m)��aE0V1&A3�&B1&D2&S0&C1S0=�m)ATZ�o;"t�H?g�a[o�xA���z����  �o>��o'��K �������я:� L�3�p�#�5���Y�k� }������$�[�H�� �~�9�����Ưد�� ������ӟ�V�	�z� ������c�Կ����
� �.���d��)�;� �Ͼ�q�������˿ <���`�G߄ߖ�IϺ� m�ϑϣ����8�J� ��n�!ߒ�M�����|��h_NITOR� �G ?�[   	EXEC1��/�25�35�45�5�5��P7�75�85�9�0�Қ�4��@� ��L��X��d��p��|�������2���2��2��2��2���2��2��2��2�23��3��3�@�;QR_GRP_�SV 1��k �(�A�z�4�~��K�������K:z�j]��Q_D��^�PL�_NAME !�3%,�!De�fault Pe�rsonalit�y (from �FD) �RR2�� 1�L6(�L?�,0	l d������ ��//(/:/L/^/ p/�/�/�/�/�/�/�/ZX2u?0?B?T?f?@x?�?�?�?�?\R<? �?�?O O2ODOVOhO�zO�O�O�OZZ`\R�?�N
�O_\TP�O:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHo_)_~o�o�o�o �o�o�o�o 2D Vhz�[omo�� ��
��.�@�R�d��v���������Џ�� Ef  Fb�� F7���  G ��!��d� �@�R�6�t����獀�l���ʝ����� ݘ����"�@� F�d���� "𩯹�ݐA�  ϩU[�$n�B�oE �� �� @D�  �?��� �?�@��A@��;f��FH� ;��	l,�	 �|��j�s�d�>���� ��� K(���Kd$2K ���J7w�K�YJ˷�Ϝ�J�	�ܿ�� @I����_f�@�z���f�γ��N������	X�l������W�S�ĽÔ��I �����5����  ����A?o�i#�;����� ���l� �Ϫ�-���ܛG�G�jѲ��@n�@�a   � � ��ܟ*�͵	�'� � H��I� �  y�Рn�:�Èl�?È=��̈́�в@�ߚЕ����D/�����̷NP�  ',���-��@
�@���?=�@A���B��  Cj�a�B�e�Ci��#�B�и�ee��^^ȹBР��P�����̠�����ADz ՟�n�3��C�i�@��R�R�Y����  ��@� ���  <���?�ff������n� ɠ#ѱ@y9G
(���I�(�@uP~����t�t����>����;�Cd;���.<߈<��g�<F+<AL�������,�d�|,�̠?fff?���?&&��@���@x��@�N��@���@T� H�ِ�!-�ȹ�| ��
`������ �//</'/`/r/]/�/��eF���/�/ �/�/m?��/J?�(�E��G�#�� FY�T?�?P?�?�? �?�?�?O�?/OO?O eOk��O�IQOG�? �O1?�OmO_0_B_T_"������A_�_@	_�_�_�_ o��A��aAn0 bФ/o C�_pUo�_�Op��؃o��o�o�o���W������oC�E�  q�H�d��؜a@q���e�F�BµWB�]�NB2�(A���@�u\?��D�������b��0�|�uR�Ｃ�
x~������Bu*�C��$�)`��$ ���GC�#���rA�U����1��eG�D�I�m�H�� I:��I�6[F����C�I��J��:\IT�H
~QF�y���p�*J�/ �I8Y�I��KFjʻCe�o�� s�����Џ���ߏ� *��N�9�r�]����� �������۟���8� #�\�G�����}����� گů���"���X� C�|�g�����Ŀ��� ����	�B�-�f�Q� ��uχ��ϫ������ ��,��P�b�M߆�q� �ߕ��߹�������(� �L�7�p�[����������s($���33:����$���3���d�,�4���@�R�wa����l�~�wa���ex����wa4 �{�� ����(L:ue%P�P~�A�O�������	����G2W} h������/����O�O7/m/[(d =�s/U/�/�/�/�/�/ ?�/1??U?C?y?�=  2 Ef9g�Fb��77�9fBX)aa)`C9A`�&`w`@-o�?w`e�O)O�?MO�Ow`�?�?�O�O�O�O9c?�0�A7h�t4w`w`!:w`xn
 �O9_ K_]_o_�_�_�_�_�_��_�_�_o#ozzQ ���h��G����$MR_CABL�E 2�h ��a�T� @�@�0�Ae��a�a�a�%�`��0�`C�`�a�O8�tB�nׇd��`�aE�4�E�#�o�f-�#��0��0�D�O��By`���Š��bED4E�c,��o�go8  ���C�0�7�d4
vے��0 �b��XE'�Z&�l�`y`r
qC�p�bHE�
v�#g�5D�Ү(�qz�lҠ`��0�q��p�b0�
v�%�c���b=%	E;h��u/o�c-��4 tH�\�?�9�K�]�o� ԏϏ��
�ɏۏ@���t?��eo �a����������b����� �����`�	 ����@������_% �*�0��6 ��ݐ����`��	�����@�������*,� ,�-�\cOM� �ii��3�� � /���%% 2345?678901i�{�! f�����������15����
��`��not se�nt3�����;��TESTFE�CSALGR  �e�qiG�1d.�š
:�� �DCbS��Q�c�u��� 9U�D1:\main�tenances�.xml��ֿq�� =��D?EFAULT-�i4~\bGRP 2�M��  =��a��{p  �%F�orce�sor� check  ���b�z��p����h5-[ �ϻ����������D�%!1st �cleaning� of cont�. v�ilat�ion��}�Rߗ+���[�ߔߦ߸����mech�caYl`������0��h5k�@�R�d��v�����(�rollAe_Ƶ����/����(�:����B�asic qua?rterly�������,�����������M��M��:C@"@GpP�a�b`i4��@�����#C���M"��{Pb�t���Sup�pq�grease���?/&/�8/J/\/��C+ ge���. batn�y`/��/h5	/�/�/��/? ?_�ѷenB'�v��/�/��/����?�?�?�?�?�G(=?O�qp"CrB1O��0�/`OrO�O�O�O��t$��Lf��C-m��A�O:�OO$_6_�H_Z_l_�t*ca�bl�Om���S<m��Q�_:�
_�_�_ oo0oo)(Ӂ/�_�_���_�o�o�o�o�ov�O@hau16�l�2r xm�<qC:��op���|���ReplaW�AfUȼ2�:�._@4�F�X�j�|�m�$%� ��o�������#���
� �.�@���d���ŏ׏ ����П����U�*� y�����r��������� 	�q��?�߯c�8�J� \�n���ϯ�����ڿ )����"�4�Fϕ�j� ��˿����������� �[�0�ϑ�fߵϊ� �߮�����!���E�W� ,�{�P�b�t����� ������A��(�:� L�^���������� ���� $s�H�� ����q����� 9]o�Vhz ���U�#�G /./@/R/d/��/�/ ��//�/�/??*? y/N?�/�/�?�/�?�? �?�?�???Oc?u?JO �?nO�O�O�O�O+J�r	 H�O�O__6M 2_@OBE:_p_>_P_�_ �_�_�_�_ o�_�_o Hoo(oZo�o^opo�o �o�o�o�o �o :z� �bA?�  @�q _����Fw�� �H;* �** @q>v �p2T�f�x�:�������ҏ��eO^C7� Տ#�5�G�	�k�}��� ُ���c�����W� �C�U�g���ß)��� ��ӯ���	��-�w� ����9�������m�Ͽ���=�O�E	A��$MR_HIST� 2�>uN�� �
 \$�Force s�ensor ch�eck  1234567890q��3����ß��N}SB� -�319.8 ho�urs RUN �9.�Y�!1st� cleanin�g of con�t. venti?lation0ÄϨ�Ϩ�-�Y���mwech��cali��%Ό4��o�D7N�t��95��1�����rolle�h�+�=�O��Y��Basic quarterly� �ߤ߶�
O4�F��(� ����b�t����� ������M�_�����:�����p���:�SK�CFMAP  .>uQ��r5��������ONR�EL  .��3���EXCFE�N��:
��QF�NCXJJOGO/VLIM8dNá ���KEY8��_PAN7����������SFSPDTYPxC��SIG�:��T1MOT�G���_CE_GRP� 1�>u\ �D�����/Ⱥ ��/�/U//y/ 0/n/�/f/�/�/�/	? �/???�/c??\?�? P?�?�?�?�?�?O)O�OMO,���QZ_E�DIT5 )TC�OM_CFG 1����[�O�O�O }
�ASI �yB3�
__+[_�O_��>O�_bHT__ARC_U���T_MN_MO�DE5�	UA�P_CPL�_gN�OCHECK ?��� ��  o.o@oRodovo�o�o �o�o�o�o�o*�!NO_WAITc_L4~GiNT�A����EUwT_E�RRs2���3��@ƱJ�����>_�)��|MO�s��}x�:Ov���8�?������ l��rP�ARAM�r�����j���5�5�G� =  r�b�t� s�X������������`֟�0����b��t�����SUM_RSPACE�����A�ѯۤ�$ODRD�SP�S7cOFFSET_CARt@��_�DIS��PEN_FILE:��7�AF�PTIO�N_IO��q�M_PRG %���%$*����M�WO_RK �yf ��춍����   ������	 �������It��RG_DSBL  ���C�{u��RIE�NTTO7 ��Cɴ A��UT�_SIM_Dy����V�LCT ��}{B �٭�ď_PEX�P=��R[AT�W dc�>�UP ���`���e�w�]ߛߩ���$�2r�L�6(L?���	l d������ &�8�J�\�n���� �����������"�4�F�X���2�߈����� ��������*�<w�Tfx��������J`�ˣG���Tz�Pg���� ��/"/4/F/X/j/ |/�/�/�/���/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?�/�/ ,O>OPObOtO�O�O�O �O�O�O�O__(_:_��O��y_�]2����_�^�_�_�W^]@^]��/ooSog�� Hgrohozo�o�o�o�o��oF`�#|`�AG�  9y����OK��1�k�����<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	 '|�Q�s�r�q/>��u �sF`�H<zH~��H3k7GL�z�HpG�9�9l7�k_B�T�F`C4T��k�H���t��-��Ae���k������s���  ��ሏ����EeBVT����dZ��g���ڏ ����q-�Fk�y�{FbZU���n@6�_  ���z��Fo��Be	'� �� ��I� ��  �:p܋=����ڟ웆�@���B�,���B��g�AgN��� � '|���g��B�*��p�BӀC׏�����@  #�B�u�&�ee�^^މB:p2���>�m�6p�Z���Dz ?o}�܏������׿�������Ǒ��� f� � � �M���*�?�ff�_8�Jφܿ 3pϑ�ñ8@�Чϵʖq.·�(����P���'��s�tL��>��/�;�Cd;���.<߈<��g�<F+<AL ��^oiΚrd@�|�r6p?fff?��?&�п�@���@x��@�N��@���@T� ��Z���ћtމ�u�� �w	�x��ti�>�)�b� M��q��������� ����:�%�^��������W���S�E�  �G�aF�� Fk���������1 U@yd���� ��q��	��{�A ��h�����a��ird��A{/w�/J/5/n/vAG�A0���":t�/ C^/�/xZ/ ލ?���/��/1??���W���t�g��pE� ~1��?04�0
1�1@�IӀ��BµW�B]�NB2�(�A��@�u\�?����������b�0�|�uR�����
�>��ؽ��Bu�*C��$�)`��? ���G�C#���r�AU����1��eG���I�m�H�� I:��I�6[F����C4OI���J�:\IT��H
~QF�y��Ol@�*J�/� I8Y�I��?KFjʻC��-? �O�O__>_)_b_M_ �_�_�_�_�_�_�_o �_(oo%o^oIo�omo �o�o�o�o�o �o$ H3lW�{� ������2�� V�h�S���w�����ԏ �������.��R�=� v�a�������П���� ߟ��<�'�`�K�]� ��������ޯɯ��&�8�#�\��3(J��g�3:a������J�3��c4�������������1��㚅ڿ��1����e���14 �{ 2�2�r�`ϖτϺϨ�J�%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ��� �������3��W�B� {�f�4���������d�A����!��1�3� E�{�i��������������  2 Efn�7Fb�7��6�B�!�!� C9� �� �0@�/`r������#x��+=�3?, V�8�v��0�0�:�0�.
 D� ����//%/7/�I/[/m//�/�:� ���ֻ�G����$PARAM_M�ENU ?2���  �DEFPUL�SE�+	WAI�TTMOUT�+�RCV? S�HELL_WRK�.$CUR_ST�YL� 4<OP9TJJ?PTB_?Y2�C/?R_DECSN 0�Ű<�?�?�?�? �?OO?O:OLO^O�O��O�O�O�O�!SSR�EL_ID  �.�����EUSE_PROG %�*q%�O0_�CCCR0��B���#CW_HOSoT !�*!HT�_=ZT��O_�Sh_zQ��S�_<[_TIM�E
2�FXU� GD�EBUG�@�+�CG�INP_FLMS�Ko5iTRDo5gP+GAb` %l�tk�CHCo4hTYPE
�,� �O�O�o# 0Bkfx�� �������C� >�P�b���������ӏ Ώ�����(�:�c��^�p�����7eWOR�D ?	�+
 �	RSc`��P�NS��C4�JO�v1��TE�P��COL�է�2��gLVP 3�����Oj�TRACECTL� 1�2��!{ ��� ��Қ�q�DT Q�2�Ǡ��D �� :��f��Ԡ�Ԡ���}�ׯ���;�4��4��4� ��;�u:�q:���;�U8�	8�
8�8�U8�8�8�8�T�@:�8�8����� ���ٱ޴���ؿ�$�6��� 
�l�~�@�R�dϞϰ� ��������
��V�h� zߌߞ߰��������� 
�,�>�P�*�<�v���*�����˶; ]+8� (��)��*������%�7�I� [�m������������ ����!��5�G�Y� k�}�������ſ�� С�*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6@ubt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀�V�߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h?�z?�?�?�?�?�1�$�PGTRACEL�EN  �1  ���0���6_UP �/���A@�1�@�1_CFG7 �E�3�1U
@�<D�0<D�ZO<C�0uO$BDEF�SPD �/L��1�0��0H_C�ONFIG �\E�3 �0�05d�D��2 �1�AaPpDsA�A�0��0�IN'@TRL ɽ/MOA8pEQPEv�E��G�A�<D�AILID(C��/M	bTGRP 1}ýI l�1�B  ������1A�33FC�� F8� E�� @eN	�A�AsA�Y��Y�A�@� 	 �vO�Fg�_ ´8cokB;`baBo,o�>oxobo�o�1>о�?B/�o�o~��o =%<��
C@yd ��"������  Dz@�I�@A 0�q� �������ˏ�� �ڏ���7�"�4�m��X���|���Ú)ґ�
V7.10be�ta1HF @�����Aq�ܢQ  �?�� �BܠP�p �C���&�B�EQ�A���Q�P�Q�� @ß[�m����<CA���0�b�@���f�������ҡ�R�ܣ�R����1�i������t<B!CeQ�KNOW_M  �lE7FbTSV ĽJ�BoC_�b� t�������������1��]aSM�SŽK ���	NB�0����ĿK���-�bb��A�R� �P����0�Ŗ��bQ+MR�S��T�iN�`��d���V]ST�Q�1 1�K
 4aMU�iǨj� K� ]�oߠߓߥ߷����� ��2��#�h�G�Y�� }�������
������,�27�I��1�#<t�H��P3^�p�����,�4���������,�5(:,�6 Wi{�,�7����,�8�!3n,�MAD�6 F�,�OVLD  �KD�xO.�PAR?NUM  �MC\/%�SCH� E�
9'!G)�3Y%UP�D/��E�/P�_C�MP_��0@�0'�7E�$ER_CH�K�%5H�&�/�+RqS���bQ_MO��+?=5_'?O�_RES_G6��:�I�o �?�?�?�?O�?O7O *O[ONOOrO�O�O�{4]��<�?�Oz5�� �O__|3 #_B_G_ |3V b_�_�_|3� �_ �_�_|3� �_�_o|3�Oo>oCo|2V 1��:�k1!�@c?��=2THR_IN�Rc0i!}�o5d�fM�ASS�o Z�gM�N�o�cMON_QUEUE �:ը"�j0��O�N� U�1Nv�+DpEND8Fqd?`yEXEo`uƅ BEnpPAsOP�TIOMwm;DpPR�OGRAM %�$z%Cp}o(/BrT�ASK_I��~O?CFG �$���K�DATA��&T���j12/ď ֏������+�=�O� a����������͟���INFO�͘�� 3t��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����
�Θ� '��FJ�a K_N��T��˶�ENBg ڽw1��2���GN�2�ڻ� P(O�=�{��]ϸ�@���v� �u�uɡd�Ʒ_EDIT ��T�����G�WER�FL�x�c)�RGA�DJ Ҷ�A�  $�?j00��a��Dqձӆ5'�?��ʨ�<u�)�%e������FӨ�2Y�R��	H;pl�G��b_�>�pAodɻt$�*�/� **:�j0�$�@�5Y�T���^��q�߈b~�L��\� n���������� �����4�F�t�j�|� ������������b LBT�x�� ��:��$, �Pb���/� ���/~/(/:/h/ ^/p/�/�/�/�/�/�/ V? ??@?6?H?�?l? ~?�?�?�?.O�?�?O O O�ODOVO�OzO�O _�O�O�O�O�Or__ ._\_R_d_�_�_�_�_�_�_�f	g�io�pWo �o{d�o�~o�ozo�B�PREF S�Rږp�p
�?IORITY�w[�}��MPDSP�q���pwUT6����OoDUCT3������OG��_T�G��8��ʯrTOE�NT 1׶� �(!AF_IN�E�p,�7�!t�cp7�_�!u�dN���!ic�mv��ޯrXYK��v����q)� ,�����p��&�	� �R�9�v�]�o����� П������*��N�`�*�sK��9}�ߢ�\��Ư ,�/6�H�������خ�At�?,  �Hp���P�b�t����u�w�HANCE �R��:�wd��连�2s��9Ks��POR_T_NUM�s�p����_CAR�TREP{p�Ω�SoKSTA�w dʷLGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_a_seiban�o \��olߒ�}߶ߡ��� ������"���X�C� |�g���������� ���	�B�-�f�Q��� u������������� ,<bM�q� ������(|L�VERSIyp��w} di�sabledWS�AVE ߾z	�2600H76%8S?�!ؿ����/ 	5(�r)og+^/y�e{/�/�/��/�/�*�,/? ��p���_�p 1��Ћ� ������Wh?z?�W*pURGE��B�p}vgu6,�WF�0DO�vƲ©vW%��4(�C�WR�UP_DELAY� �\κ5R_HOT %Nf�q׿�GO�5R_NORM�AL&H�r6O�OZGS�EMIjO�O�O(qQ/SKIPF3��W3x=_98_J_\_] �_�_{_�_�_�_�_�_ �_	o/oAoSoowoeo �o�o�o�o�o�o�o +=aOq�� ������'���7�]�K�������)E�7$RA{���K/��zĀÁ_PARA�M�A3��K @�.�@`�61�2C�<��y��C��6$�BÀBTIF��4`�RCVTMO�Uu�c��ÀD�CRF3��I ��+UC�AqD���2=\�(�?��]�
�ޅ���4��+_����;�Cd;���.<߈<�g��<F+<L�A��Ѱ��d�u�L� ������ϯ�����)�;�M�_���RDI�O_TYPE  �M=U�k�EFPO�S1 1�\�
 	x4/�����+� $/<��$υ�pϩ�D� ��h��ό��'����� �o�
ߓ�.ߤ�Rߌ� ������5���Y��� i��*�<�v���r��� �������U�@�y�� ��8���\������������?��c����2 1�KԿX��T�x��3 1� ����nY�S4 1�'9K��/�'/�S5 1���/�/�/|�/:/S6 1�Q/�c/u/�/-??Q?�/S7 1��/�/
?D?��?�?�?d?S8 1�{?�?�?�?WOBO{O��?SMASK 1�L��O�D�GXN�O���F&�^��MOCTEZ�Ż��Q_ǁ��%]pA݂��PL_RANG!Q]�_QOWER �ŵ��P1VSM_DRYPRG %ź�%"O�_�UTART� �^�ZUME_PRO�_�_4o���_EXEC_EN�B  ��#�e�GS�PD`O`WhՅjbT3DBro�jRM�o�h�INGVERSI�ON Ź�#o�)I_AIRPURhP �O(�M�MT_�@T�P#_�ÀOBOT_ISOLC�NTV@A'q�huNAME�l���o�JOB_ORD_NUM ?�X�#qH76�8  j1Zc@n�r
�rV�sw��r�?�r�?�r�pÀPC�_TIMEu�a�x�ÀS232>R1��� LTE�ACH PENDcANw�:GX��!O Maint�enance C�onsj2����"���No UseB�׏������1�8C�y�V�NPO�P@��YQ�cS�C7H_L`�%^ ��	ő��!UD�1:럒�R�@VA#IL�q@�Ӏ�J�Q�SPACE1 2�ż ��YRs�i�@Ct�YRԀ'{��?8�?��˯ ����"���7�2�c� u�����G���߯ѿ� ���(��u�AC�c� u�����Ͻ�߿���� ���(��=�_�qσ� ��C߹������߱�� $��9�[�m�ߑߣ� Q������߭��� ��� 	�W�i�{���M��� ����5���.S� e�w�����I����� ��*?as ��E����� /&//;/]o�� ����/2/�/?"? �/7?Y/k/}/�/�/O? �/�/�?�?�?O0OO~KA��*SYPp�M*�8.302�61 yB5/21�/2018 A� �WPfG|�H�_�TX`� !$C�OMME��$USAp �$ENABLED�Ԁ$INN`QpI�OR�B�@RY�E_�SIGN_�`�AP��AIT�C�BWRKz�BD<�_TYP�CRINDXS�@W��@%VFRI{�_G�RPԀ$UFR�AM�rSRTOOL�\VMYHOL�A�$LENGTH_�VTEBTIRST��T  $SE�CLP�XUFINV�_POS�@$�MARGI�A$�WAIT�`�ZX2l�\�VG2�GG1�AAI�@�S�Q	g�`_WR��BNO_USE_�DI�BuQ_REQ��BC�C]S$CUR_TCQP�R"a^f� �GP_STA�TUS�A @ ��A3`�BLk�H$�zc1�h�P@���@_��FX �@E_MLT_CT�C�H_�J�`CO�@O�L�E�CGQQ$W��@w�b#tDEA�DLOCKuDELAY_CNT�a�3qGt�a$wf �2 R1[1T$X<�2[2�{3[3$Zwy�q%Y�y�q%V0�@�c�@�b$V�`�R�V�UV3oh>b�@� � �d�0arMSKJ�LgWaZ�C`�NRK�PS_RATE�0$���S
`�Qv�TAC��PRD����e�S*��a4�b u �DG�A 0�P��flp bquS2�ppI�#`
`�P �
�S\`  }�A�R_ENBQ� �$RUN?NER_AXI�<`�ALPL�Q�RU�TH�ICQ$FLI�P7��DTFERE�N��R�IF_CH�SU�IW��%V)�G!1����$PřA�Q�P�ݖ_JF�PR�_P�	�RV_D�ATA�A  {$�ETIM����$VALU$��	�OP_  � �A  2� �SC*��	� �$ITPa_!�SQ]PNPOU}��o�TOTL�o�DS}P��JOGLIb�N�PE_PKpc�Of�ji��PX]PTAS��$KEPT_M#IR��¤"`M�b�APq�aE�@�y�`q�g@١c�q�PG��BRK6�x���L�I��  ?�SJ�q��P�ADEz�ܠBS{OCz�MOTNv�DUMMY16Ӂ�$SV�`DE_�OP��SFSPDO_OVR
���@�LD����OR��T-P8�LE��F����6��OV��SF��F����bF�d�ƣ&c)��fQc�LCHDLY>��RECOV���`���W�PM��gŢ�R�O������_F�?�� @v�S �NVE�R�@�`OFS�PC,�CSWDٱc�ձ��X�B����TRG�š��`E_FDO��MOB_CM}���B���BLQ�¢	�Q�̄V�za�BUP�g��G
��AM���@`K�̊�e�_M!�d�AMxf�Q��T$CA����DF���HBKXd�v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�3�A��ATIO�0��͠��US����WaAB��R+c�`tá`xDؾA��_AUXw�?SUBCPUP���S�`����3Եжc���3�FLA�B�HW_Cwp"�Ns&�]s�Aa��$UNI�TS�M�F�ATT�RIz�Z�CYC=L�CNECA����FLTR_2_F�I��TARTUP`Jp����A��LP�������_SCT*cF�_F�F_P���b�FqS��+�K�CHA/Q���*�d�RSD���Q����Q���_T�H�PROr���հE#MPJ���G�T�� �Q�DI��@y�RAILAC4/�bMX�LOf�xS��ځ���拁���+PR#�S`app��C� 	��F�UNC���RIN�`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ng�DAQ�B�rkL�D�र&q�M�K���TI���j���$�@RIA_S�W��AF��Pñ�#��%%�p9r1��MsOIQ���DF_~P�(�PD"LM-�F�A�PHRDY�DORG�H; _QP�>s%MULSE~Pz�T��*�� J��Jײ���FAN_AL�MLVG��!WRN�%HARDP��Uc�O�� K2$SHADOW]�kp�a02���� STOf�+�_,^�w�AU{`R��eP_SBR�z5����:F�� �3MPINF?�\�4��3gREGV/1DG�b+cVm �C�CFL(��?�DAiP��ҌZ`�� �����Z�	� �P(Q$�A�$Z�Q V�@�[�
o� ��EG߀o���kAAR���㌵�2�axG��AXEROB��RED���W�QD�_�Mh�S�YA��AF��FS�GW�RI�P~F&�STRP����E�˰EH�)�$�D�a\2kPB6P��t=V��Dv�OTO�19)���ARYL�tR0�v�3���FI&�ͣ?$LINKb!\�J�Q�_3S���E���QXYZ2�Z5N�VOFF���R�RJ�XxPB��d0s�G�cFI�03g��������_J ��'�ɲ�S&qR0LTV[6���aTBja�"�b�C���DU�F7.�TUR� X��eĂQ�2XP�ЊgFL��E���x@�`�U9Z8����� 1	)�K��Mw��F9��劂����ORQj��G;W3���#�Ґd ���uz����1�tOVE�q_�M��ё?C�uEC �uKB�v'0�x-�wH� �t���& `��qڠ �B�ё�u�q�wh�EC�h����ER��K	B�EP����AT�K�6e9e�W����AXs�'��v�/� �R ����!�� � �P��`��`�3p�Yp�1�p�� ��  �� (�� 8�� H��  X�� h�� x�� ����ޙ�DEBU�$�%3�I��·RAB����ٱ�sV��� 
d�J、��@� ��������Q���a�� �a��3q��Yq+$�`%"\<�cLAB0b�u�'�GRO���b<��B_s��"Tҳ *`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθ0uݸ��PNT0��?�SERVE �Z@� $`EAV�!�PO����nP�!�P@�$!Y@ � $>�TRQ"�b
=��BG�K�%"�2\��� _ � l��5�D6ER)RVb(�I��V0`;�N��TOQ:�7�L�@P
�R��e G�%�Q����<�50F� ,h�`�z�>�RA�? 2 d!�����S�  M��phxU �� <�OCu�G�  ��C�OUNT6Q9�P@F�ZN_CFGF�# 4#��6��TG4�_�=�����ӎ�VC ���M �"��`$6��q ��FA E� &��X�@�����H��A����AP���P@HEL�0��� 5b`B_B;AS��RSR�6E�CSH����1�Ǫ��2��3��4��5*��6��7��8��}�ROO����P�PNLEA�cAB)ë ��ACKu�INO�T��(B$UR0� =��_PU��!0��OU+�Pd�8j��� V���TPFWD_KcAR��� ��RE(�� P�P�>QUE�:RO�p�`r0P1I� x�j�P�f��6�QSEM��0��� �A��STYL�SO j�DIX�&������S!_TMCMA�NRQ��PEND�It$KEYSWITCH���k�HE�`BEATM683PE{@LE��>�]��U��F��S~pDO_HOM# �O�@�EF�pPR�aB�A#PY�C� Ox�!���OV_M|b<<0 IOCM�dfFQ���k�HKYAG D�Q�7��UF2���M���p�cFO;RC�3WAR�"��OM|@  @�S�#o0U)SP�@1*�2&3&4E���*T�O��L���8OUNLOv�D4K$�EDU1  �S�Y�HDDNF� �M�BLOB  �p�SNPX_;AS�� 0@�0|��81$SIZ�1�$VA{���MU/LTIP-��# �A� � A$��� /4`�BS���0�C���&FRIF�BO�S���3� N=F�ODBUP߰�%@3;9(�^ы�Z@� x��SI��TqEs�r�cSGL�1	T�Rp&�Н3B��@��0STMTq�3P�g@VBW�p�4SHsOW�5@�SV���_G�� 3p$PaCJ�PИ���FB�-PHSP AW�E�P@VD�0WC�; ���A00��PB  XG XG XG$ XGU5VI6VI7VI8VI9VIAVIBVI�XG�YF@`XGFVH��X�bI1oI1|I1�I1��I1�I1�I1�I1��I1�I1�I1�I1��I1Y1Y2UI2�bI2oI2|I2�I2��I�`�X�I2p�X�I2��I2�I2�I2�I2BY2Y�p�hbI3oIU3|I3�I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3YU3Y4�i4bI4oIU4|I4�I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4YU4Y5�i5bI5oIU5|I5�I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5YU5Y6�i6bI6oIU6|I6�I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6YU6Y7�i7bI7oIU7|I7�I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7YY7T�VP� UD�#y"ՠ��
<A62���t�R��CSMD� ��M5�Rv�,]��Q_h�R���pe����<�YSL��>�  � �%\2 ��+4�'��W�BVALU��b��'�z��FH�ID_L����HI��I���LcE_��㴦�$0�C�SAC�! h� �VE_BL�CK��1%�D_CPU5ɧ 5ɛ ������C�� ��R " � PWj���#0��LA�1S�Bћì���RUN_FLG�Ś����ĳ  ����������H����ХĔ�TBC2���# � @ B ��e �S�8=�F'TDC����V���3d�Q�THF�����R�L�ESERCVE9��F��3�2��E��Н�X -$��LEN9��F���f�RA��W"G�WI_5�b�1��д2�MO-�T%S60U�I�k�0�ܱF����[�DyEk�21LACEi�0�CCS#0�� _M�A� j��z��TCV����z�T�������.Bi�'A�z�'AJ$h�#EM5���J��@@Ri�V�z���2Q `�0&@o�h��JK��VK9��{���щ�J0����JJ��JJ��AAL���������4��5�ӕ NA1������.�LD��_�1* �CF�"% `�GRO�U���1�AN4�C��#m REQUIR��EBU�#��6�7$Tk�2$���pzя #�& \�/APPR� C� 0��
$OPEN�C'LOS�St��	ri�
��&' ��MfЩ���W"-_M	G�7CB@�A�ܸ�BBRK@NO�LD@�0RTMO!_5ӆp1J��P��������������6��1�@� m1�#�(�# �����'��+#PATH''@!6# @!�<#� � '��1�SCA���6I�N��UCJ�[1� C0@UM�(Y ��#�"������*���*��� P�AYLOA~J2=LؠR_AN^�3�L��91�)1AR?_F2LSHg2B4LO4�!F7�#T7�#ACRL_�%�0ȏ'�$��H��.�$yHA�2FLEX�u�J!�) P��2�D߽߫���0��* :����z�FG�]D����z���%�F1]A�E�G4�F�X�j�|���BE������ ������(��X�T*� A���@�XI�[�m�\At�T$g�QX<�=�� 2TX���emX������ ������������t+	�J>+ �-�`K]o|�٠AT�F�4�ELFPѪs��J� *� JEmC3TR�!�ATN�v�zHAND_VB�.��1��$, $�8`F2Av���S�W�
"-� $$M*0.�]W�@lg��PZ����A�� � 1����:AK��
]AkAz��LN��]DkDzPZ G��C�ST_K�lK�N}DY��� A�� ��0��<7]A<7W1�' ��d�@g`�P��������"
"J"�. M�2D%"��xH����ASYMj%0�� j&-��-W1�/_�{8� �$���@��/�/�/�/ 3J<��:9�/�89�D_V�I�v����V_�UNI�ӛ��cD1J ����╴�W<��n5Ŵ �w=4��9��?�?<Œuc�4�3��%�H���/�j��0�SDIzuO�Ćќk�>0 �`��I��A��#���@ģ����@��IPl� 1o � /�ME.Q�p��9�ơT}�P�T�;pG �+ Gt � ���'��T�0� $DUMM�Y1��$PS_f�@RF�@;�$b��'FLA@ YP�(c|��$GLB_TP�ŗ���9 8P�q��2 X� z�!ST9�� SB}RM M21_V�T$SV_ER*01O�p����CL����eAGPO��f�GL~�;EW>�3 4H �W$YrZrW@�x�A1+�A���";�"�]U&�4 8`NZ��"�$GI�p}$&� -� �Y�>��5 LH {��}$�F�E��NEAR�(PN�CF��%PTAsNC�B	!JOG�@� 69�$J�OINTwa?pd�MwSET>�7  x�E��HQtpS{r��up�>�8� �pU�.Q?�� LOCK�_FOV06���BG�LV�sGLt�TE�ST_XM� 3�EMP�����_��$U&@%�w`24� Y��5��2�d��3��CE- ���� �$KAR�QM��T�PDRA)�����VcECn@��IU���6��HEf�TOOiL�C2V�DRE 'IS3ER6��@�ACH� 7?O�x �Q�29Z�H I��  @$RAIL_BOXEwa��ROBO��?���HOWWAR�1�_�zROLM j��:qw�jq� �@� O_Fkp! �d�l>�9�� �R O8B: �@�	""�OU�;��Һ�3ơ�r�q_�/$PIP��N&`H��l�@��#@CORDEDd�p >f��fpO�� < D ��OB⁴sd����Kӕ���qS;YS�ADR�qf���TCHt� =� ,8`ENo��1A
k�_{�-$Cq7�f��VWVA��> Ǥ  &��PR�EV_RT�$�EDITr&VSHWRkq�֑ &R:�%v�D��JA�$�a?$HEAD�6�4� �z#KE:�E��CPSPD�&JM%P�L~��0R*P�ģ?��1%&I��S�rC�pNE; �q�wOTICK�C��M�1�3�3HN��@ �@� 1Gu�!_GP8p6��0STY'"xLO��O2l2?�_A t 
m G3%S%$R!{�=��S�`!$��w`���ճ�r��Pˠp6SQU��x�E��u�TERC��0��TSUtB ����hw&`gw�Q)b�pO����@IZ��4{��^�PR�kј�B1XPU���E_�DO��, XS�KN~�AXI�@���UR�pGS�r� ^0�d&��p_) �ET�BQPm��o��0Fo�2�0A|���Rԍ���aOSR�Cl>@P��b_�yU r��Y��yU��yS��yS ���UЇ�U���U���U �]��Ul[��Y�bXk�]Cm�����YR�SC�� D h��DS~0��Q�SPL���eATހ���A�]0,2N�ADDRE�S<B} SHIF�{s��_2CH�pr�I��=q�TVsrI��E"���a�Ce�
��
;�VW�A��'F \��q��0l|\A@�rC�_B"R{z�p�ҩq�TXSCWREE�Gv��1TINA���t{�����A�b?�H T 1�ЂB�����I��Ap��BE�y RRO������� B��D1UE4I �g�!p�9S��RSM]0�GUNEX(@~Ƴ�j�S_S�ӆ��Á։�ģ��ACY�0� [2H�pUE;�J�¸���@GMT��L�ֱ�A��O	�BB�L_| W8���K ���0s�OM��L1E/r��� TO!�s��RIGH��BRD<
�%qCKGR8л��TEX�@����WIDTH�� �B[�|�Z<��I_��Hi�� L 8K���_�!=r���R:�_���Yґ��O6q�M�g0紐U��h�Rm��LUMh��FpGERVw �P����`�N��&�GEKUR��FP)�)� �LP��(RE%@�a)�ק�a�!��f �5*�6�7�8Ǣ#B@�É@���tP�fW��S@M�USR�&�O <����U8�Qs�FOC)��PRI;Qm� :����TRIP�m�SUN����Pv��0���f%��'���@�0 �Q����AG ��0T� �a>q�OS�%�RPo���8�R/�A�H�L4����	U¡�SU�g��¢�5��OFF���T��}�O�� 1�R�����S�GU�N��6�B_S�UB?���,�SRT�N�`TUg2��mCO9R| D�RAUrPE�yTZ�#'�VCC���	3V AC36�MFB1�%d�PG� �W (#��ASTEM�����0�PE��T3G�X y�\ ��MOVEz�A��AN�� ���|M���LIM_X�� 2��2��7�,�����0ı�
�BVF�`EӐ��~��04Y��IQB�7���5S��_Rp� 2��� WİGp+@��}СP��>3�Zx ����3���A�ݠCZ�DRID���ѡVy08�90� De�MY_UBYd���6��@��!��X��GP_S��3��L�K�BM,�$+0DE�Y(#EX`�����U/M_MU� X����ȀUS�� ���G0`PACI���а@ ��:��:,�:����CRE/�3qL�+���:[��TARG"��P�r��R<��\ d`��A��$�	4��AR��SW2 ��-��@Oz�%qA(7p�yREU�U�01�X,����HK�2]g0��qP� N� �E9AM0GWOR��ާMRCV3�^ U���O�0M�C�s�	���|�REF _���x(�+T� �� �������3_RCH4(a�P�Ѐ��hrj�NA�5��0�_ ��2����L@��n�@@OU~7w6���Z��a2[��R1E�p�@;0\�c�a�'2K�@SUL��]2��C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��PQ5I�]7q�}�Tg`�4D`�0.`0�APg_HUC�5SA��CMPz�F�6�5�5
�0_�aR��a�1I�\!X�9�qVGFS���ad ��M8��0p�UF_x��B� �ʼ,RO��Q��'l����UR�3GR�`.�3IDp���)��D�;��A��~�IN"��H{D���V@AJ���S͓UWmi`=�����TYLO*��5����bt� +�cPA� �cCACH�vR�U@vQ��Y��p�#CF�-I0sFR�XT���VNn+$HO����P !A3�XBf�(1 ����$�`VPy� ^b_'SZ313he6K3he12J�eh chG�ch�WA�UMP�j��IkMG9uPAD�i�iIMRE�$�b_SIZ�$P����0 ���ASYNBUF��VRTD)u5tq~ΓOLE_2DJ�(Qu5R��C��U��vPyQuECCUl�VEMV �U�r�WV�IRC�aIuVTP G���rv1s��5qMP#LAqa��v�V0��cm� CKLA�S�	�Q�"��d ! �ѧ%ӑӠ@}¾�q$�Q���Ue |�0!�rSr�T�#0! ���r�iI��m�vK�BG��VE�Z�P�K= �v�Q�&�_H�O�0��f � �>֦3�@Sp�SLO�W>�RO��AC�CE���!� 9�VR`�#���p:���AD������PAV�j�� D:����M_B"���N^�JMPG ��g:�>#E$SSC��F��vPq��hݲvQS��`qVN��LEX�c�i T`�sӂ�ܗQ�FLD �DEsFI�3�02����:|"P2�Vj'� �A��V�4[`MV_PIs��t`���A�@��FI��|�Z��Ȥ�����A����A��~�GAߥ1 LsOO��1 JCB�इXc��^`�#PLA!NE��R��1F�c�����pr�M� [`������S����f����A@f��R�Aw�״tU�΁pRKE��d�VA{NC�KL�V��.�� k���ϲ��BR_AA� l���2� ��p�#Hć�m# h���O K�$��d����kЍ0OU&Aʞ"A�
p�pSK��TM@FVIEM 2�l ��P=���n� <<��dK�UMKMYK1P��`mD��ACU��z#AU��o $���TIT�$P�R����OP����VSHIF�r�p`J�Qsԙ�fO�xE$� _R�`U �#����s��q����@��G�"G�޵'�T��$�SCO{D7�CNTQ i�l�>a�-�a� ;�a�H�a�V���1�*+�2u1��D�����  � SMO"�Uq��a�JQ���K��a_�R[�r�n�*@LIQ�AA/`/�XVR��s�n�yTL���ZABC�Ct�t�c�
|!�ZIP��u���L�VbcLn"�Z�MPCFx�v:��$�� ���DMY_LN�������@y�w Ђ(a�u� M�CM�@CbcCAR�T_�DPN� O$J71D���=NGg0Sg0�BU�XW� ��UXEUL|ByX����	�����xC 	���m�YH�}Db  y 80<���0EIGH�3n�#?(� H����$�z ���|�����$%B� Kd'��_��L3�RVS�F`���OVC�2'�$|Ј>P&��
q���5D&�TR�@ �VD���SPHX��!{ ,p� *<�$R�B�2 2 ����C!�  �@V+| b*�c%g!��b)g"�`�V*�,8�?� V+�/V.�/�/?�/�/V(7%3@/R/d/v/�/ 6?�/�/�?�?�?O4OOION;4]?o?�?�? �?SO�?�?�O_�O0_Q_8_f_N;5zO�O�O �O�Op_�O_o8o�_ MonoUo�oN;6�_�_ �_�_�_�oo%o4U@j�r�N;7�o �o�o�o�o� BQ��r�5���������N;8 �����Ǐ=�_� n���R���ş��ڟN;�G � џ�
����?��� W�i�{�������ï� .�������A��dW�<�N�|������� Ŀֿ�ޯ���0� B�_�R�d�꿤϶��� ����������*�L� ^��rτ�
������� �����&�8�J�l��~� `ҟ @ �з����ߩ��-����&�,���9� {�����a��������� ������A'Y �������@��a#1�
����N;_MODE � ��S "��[�Y�B���
/\/*	|/�/R4CWORK_AD��	��DT1R  ����� �/� _?INTVAL�+$���R_OPTI[ON6 �q@�V_DATA_G�RP 27���D��P�/~?�/�?�9 ��?�?�?�?OO;O )OKOMO_O�O�O�O�O �O�O_�O_7_%_[_ I__m_�_�_�_�_�_ �_�_!ooEo3oioWo yo�o�o�o�o�o�o �o/eS�w �������+� �O�=�s�a������� ͏���ߏ��9�'��I�o�]�����$S�AF_DO_PULS� �~������CAN_TIM�����ΑR ��Ƙ�E��5�;#U!P"�Z���� �?E�W� i�{�����.�ïկ篰����'(~�"T"2F���dR�I�"Y��2�o+@a얿 ����)�u��� k0ϴ���_ ��  T� � �2�D�)�?T D��Q�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ�x/V凷������߽��R�;��o �W�p��
�t��Diz$�� �0 � � T"%!������� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FX ��࿁����� ��/`4�=/O/a/ s/�/�/�/�/�/�/�!!/ �0޲k�ݵu�0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o k$o6oHoZolo~o�o �o�o�o1/�o�o  2DVhz�/5? ��������&� 8�J�\�n��������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c�u��� ���`Ò� ϯ����)�;�M� _�q���������˿ݿ�� ����3� ����&2,��	�12345678�v�h!B!���2�Ch��� 0�ϵ���������� !�3�9ѻ�\�n߀ߒ� �߶����������"� 4�F�X�j�|�h�K߰� ��������
��.�@� R�d�v����������� ���*<N` r������� &��J\n� �������/ "/4/F/X/j/|/;�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�/�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_�?L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o=_ �o�o�o�o�o�o  2DVhz�����h������u��o.�@�R���Cz�  B��   ����2&� �� _�
���  	�_�2�Տ�X���_�p������ďi�{������� ß՟�����/�A� S�e�w���������N� �����+�=�O�a� s���������Ϳ߿�@��'�9�K�_��丁��<v�_��$S�CR_GRP 1�
� ��� �t ���� ��	 /������� ���������_����8��)�a����&�?DE� DW8����l�&�G�CR-�35iA 901�23456789}0��M-20���8��CR35 ���:�
��������������:֦����G���&������	��]�o����:�?��H���>������������&���ݯ:��j�����g������B�t�Ɛ��������A���� c @�`��@� N( ?�=��Ht��P
��F@ F�`z�y���� �� �$H���Gs^p��B��7��/�0/ /-/f/Q/�/u/�/�/ �/8���P�� 7%?�����"?W?-2?<���]? H�1�?t�ȭ7�������?-4A, �&E@��<�@G�B-1  3OZOlO-:HA�H�O\�O|O P�B(�B��O�O_��EL_D�EFAULT  ������`SHOTST�R#]JA7RMIPO�WERFL  �i�/UYTWFDO�$V /URRVE�NT 1�����NU L!D?UM_EIP_-8��j!AF_I�NE#P�_-4!FIT�_->�_;o!���`o �*o�o!�RPC_MAINĈojh�vo�o�cVI�S�oii��o!�TPpPU�Yd�k!
PMON?_PROXYl�VAeZ�2r��]f���!RDM_S�RV��Yg�O�!#R��k��Xh>���K!
�`M��\i����!RLSYN�C�-98֏3�!�ROS�_-<�4�"��!
CE4pMOTCOM���Vkn��˟!	��CONSd̟�Wl���!���WASRC��Vm��c�!��USBd��XnR���Noӯ� ������!��E��i��0���WRVICE�_KL ?%�[� (%SVCPGRG1��-:Ƶ2ܿD�˰3�	�˰4,�D1�˰5T�Y�˰6|���˰7�ϩ�˰�����9����ȴf�!� ˱οI�˱��q�˱� ��˱F���˱n���˱ ���˱��9�˱��a� ˱߉��7߱��_� �������)�� ��Q����y��'�� �O����w����� ����˰��İ d�c������ =(as^� �����/�/ 9/$/]/H/�/l/�/�/ �/�/�/�/�/#??G? 2?k?V?}?�?�?�?�? �?�?O�?1OCO.OgO RO�OvO�O�O�O�O�O�	_�O-_��_DEV� �Y�M{C:5Xd�GTGRP 2SVK ���bx 	� W
 ,�PK 5_ �_�T�_�_�_o�_'o 9o o]oDo�ohozo�o �o�o�o�o�o5{ �_g����� �����?�&�c� u�\�������Ϗ��� J\)���M�4�q��� j�����˟ݟğ�� %���[�B��f��� ���ٯ�������3� �W�i�P���t���ÿ ���ο���A�(� e�L�ί��RϿ��ϸ� ����� ��O�6�s� Zߗߩߐ��ߴ���� ��'�~ϐ�]���h� ������������� 5��Y�@�R���v��� ������@�	��? &cu\���� ����;M4 qX������� /�%//I/[/B// f/�/�/�/�/�/�/�/ �/3??W?�L?�?D? �?�?�?�?�?O�?/O AO(OeOLO�O�O�O�O��O�O�O�O_iV ��NLy�6 *� 		S=>���+c"_VU@Tn_Y_B����B�2�7J�j~Q´~_g_��_�Q%JOGGGING�_�^7T(?VjZ�Rf��Y���/e�_%o7e�Tt�]/o�o{m�_�o �m?Qi�o�o;)Kq%��o�}o s������9� {`��)���%���ɏ ���ۏ�S�8�w�� k�Y���}���ş��� +��O�ٟC�1�g�U� ��y�������'��� �	�?�-�c�Q���ɯ ����w���s���� ;�)�_ϡ���ſOϹ� ����������7�y� ^ߝ�'ߑ�ߵߣ��� �����Q�6�u���i� W��{������=� �M���A�/�e�S��� w������������ =+aO���� ��u���9 ']���M�� ����/5/w\/ �%/�/}/�/�/�/�/ �/=/"?4?�/?�/U? �?y?�?�?�??�?9? �?-OO=O?OQO�OuO �O�?�OO�O_�O)_ _9_;_M_�_�O�_�O s_�_�_o�_%oo5o �_�_�o�_[o�o�o�o �o�o�o!coH�o {������ ; �_�S�A�w�e� ������я���7��� +��O�=�s�a����� �П�����'�� K�9�o�������_��� [�ɯ���#��G��� n���7���������ſ ����a�Fυ��y� gϝϋϭϯ�����9� �]���Q�?�u�cߙ� �ߩ���%���5���)� �M�;�q�_���߼� �߅������%��I� 7�m������]����� ������!E��l ��5������ �_D�we �����%
// ���=/s/a/�/�/ �/��/!/�/??%? '?9?o?]?�?�/�?�/ �?�?�?O�?!O#O5O kO�?�O�?[O�O�O�O �O_�O_sO�Oj_�O C_�_�_�_�_�_�_	o K_0oo_�_co�_so�o �o�o�o�o#oGo�o ;)_Mo��� �o����7�%� [�I�k��������� �ُ���3�!�W��� ~���G�i�C����՟ ���/�q�V������ w��������ѯ�I� .�m���a�O���s��� ����߿!��E�Ͽ9� '�]�Kρ�oϑ��� ��Ϸ����5�#�Y� G�}߿Ϥ���m���i� �����1��U��|� ��E���������	� ��-�o�T������u� ����������G�, k���_M�q�� �����% [Im���	 ���//!/W/E/ {/��/�k/�/�/�/ �/	???S?�/z?�/ C?�?�?�?�?�?�?O [?�?RO�?+O�OsO�O �O�O�O�O3O_WO�O K_�O[_�_o_�_�_�_ _�_/_�_#ooGo5o Wo}oko�o�_�oo�o �o�oC1Sy �o��oi���� �	�?��f�x�/�Q� +���Ϗ�����Y� >�}��q�_������� ˟���1��U�ߟI� 7�m�[�}����ǯ	� �-���!��E�3�i� W�y�ϯ��ƿ����� ���A�/�eϧ��� ˿UϿ�Q�������� �=��dߣ�-ߗ߅� �ߩ��������W�<� {��o�]����� ����/��S���G�5� k�Y���}��������� ������C1gU ������{��� �	?-c��� S������/ ;/}b/�+/�/�/�/ �/�/�/�/C/i/:?y/ ?m?[?�??�?�?�? ? O??�?3O�?COiO WO�O{O�O�?�OO�O _�O/__?_e_S_�_ �O�_�Oy_�_�_o�_ +oo;oao�_�o�_Qo �o�o�o�o�o'io N`9��� ���A&�e�Y� G�i�k�}�����׏� ��=�Ǐ1��U�C�e� g�y����֟���	� ��-��Q�?�a���ݟ ��퟇��ϯ��)� �M���t���=���9� ��ݿ˿��%�g�L� ����mϣϑϳ��� ����?�$�c���W�E� {�iߟߍ߯������ ;���/��S�A�w�e� ������������� +��O�=�s������ c�����������' K��r��;��� ����#eJ� }k����� +Q"/a�U/C/y/ g/�/�/�//�/'/�/ ?�/+?Q???u?c?�? �/�?�/�?�?�?OO 'OMO;OqO�?�O�?aO �O�O�O�O__#_I_ �Op_�O9_�_�_�_�_ �_�_oQ_6oHo�_!o �_io�o�o�o�o�o)o Mo�oA/QSe�����%{,p��$SERV_M�AIL  +u�!��+q�OUTP�UT�$�@��RV 2�v  $� (�q�}���SAVE7�(�TOP10 2W�� d 6 	*_�π(_����� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ�ݷ��YP��'�FZ�N_CFG N�u$�~���~�GRP 2��D� ,B   �A[�+qD;� B}\��  B4~��RB21��H7ELL��u���j�k�2�����%RSR�������
� C�.�g�Rߋ�v߈��� ������	���-�?�Q��  �_�%@Q���_���,p1����ޖ�g��2,pd����HKw 1�� �� E�@�R�d��������� ��������*<�e`r���OMM� �����FT?OV_ENB�_����HOW_REG�_UI�(�IMI_OFWDL� ��^�)WAIT� ��$V1�^�NwTIM����VA�_)_UNcIT����LC�TRYB�
�M�B_HDDN 2W� 2�:% 0 �pQ/�qL/^/�/�/��/�/�/�/�/�"!O�N_ALIAS k?e�	f�he� A?S?e?w?�:/?�?�? �?�?�?OO&O8OJO �?nO�O�O�O�OaO�O �O�O_"_�OF_X_j_ |_'_�_�_�_�_�_�_ oo0oBoTo�_xo�o �o�o�oko�o�o ,�oPbt�1� ������(�:� L�^�	���������ʏ u�� ��$�Ϗ5�Z� l�~���;���Ɵ؟� ���� �2�D�V�h�� ������¯ԯ���
� �.�ٯR�d�v����� E���п���ϱ�*� <�N�`�r�ϖϨϺ� ��w�����&�8��� \�n߀ߒߤ�O����� ������4�F�X�j� |�'���������� ��0�B���f�x��� ����Y������� ��>Pbt�� ����(: L�p����c �� //$/�H/Z/ l/~/)/�/�/�/�/�/��/? ?2?D?V?]3��$SMON_DE�FPRO ����1� *SYST�EM*0m6RECALL ?}9� ( �}0c�opy mdb:�*.* virt�:\tmpbac�k\=>147.�87.149.4�0:10296 <�6�95172]?O�+M}4x�2fr:\�?I@�?�1�?O�O.�O }5?EaGOYO��6uO�O_*_}
x�yzrate 61 �O�O�O _�_�_�6E?W__192  �_q_�_o&o9^�_�_ �_ o�o�o6E�_�59308 ^opo�o�%8C8�2�3ou�tput\tcp�serv3.pc��0: over �=>370278��0357235 ��o��.ACs:o�rderfil.dat�?�ox	��.M/�?��i������7D3?OR_�ms��� �(�;I�O؏�f�� ����<N`r��� '���U�p������ 8�J�e�n����#��� I�[��������4�F� W�j�|���2�D�ͯ h����ϝϰ�¯]�� x�	��.�@�ӿd��� ߙ�,߾�O�a�t߆� �)�<�N������� ���U���p���%� 8�����n� ������� G�Y���~�!4oF_ ���������_�o�17516�no��$7Dtpdisc 0�������7Dtpconn 0InXj|//��9?�Q�G� ��/�/���?Y/�p/ �/?%?8OK]��/ ?�?�?�OM?_?� u?؇?O*O}<��te�st_ԑerٜ1�62791424�:263469  �?�O�O2/D/�/�zO __�/�/�O�/�O�_ �_.?@?�?d?v_�_o �_�?�_�_�2�_�o�o �O�O�Oaowo�o-_�?_�oc_�o����$SNPX_AS�G 2�����q� P� 0 '%�R[1]@1.1,��y?��s%�!� �E�(�:�{�^����� ��Տ��ʏ���A� $�e�H�Z���~���џ ����؟�+��5�a� D���h�z�����ů� ԯ���
�K�.�U��� d�������ۿ���� ��5��*�k�N�uϡ� ���ϨϺ������1� �U�8�Jߋ�nߕ��� �����������%�Q� 4�u�X�j������ �������;��E�q� T���x��������� ��%[>e� t������! E(:{^�� ����/�/A/ $/e/H/Z/�/~/�/�/ �/�/�/�/+??5?a? D?�?h?z?�?�?�?�? �?O�?
OKO.OUO�O dO�O�O�O�O�O�O_ �O5__*_k_N_u_�_ �_�_�_�_�_�_o1o oUo8oJo�ono�o�o��d�tPARAM ��u�q W�	��jP�d9p��ht��pOF�T_KB_CFG�  �c�u�sOP�IN_SIM  �{vn��p��pRVQSTP_DSBW~r"t��HtSR Zy� � & RO�B195_SERgV M���v�TOP_ON_ERR  uCy8��PTN Zu�k�A4�RI�NG_PR�D���`VCNT_GP� 2Zuq�!px 	r��ɍ���׏���wVD��RP 1�i p�y�� K�]�o���������ɟ ۟����#�5�G�Y� ��}�������ůׯ� ����F�C�U�g�y� ��������ӿ��	� �-�?�Q�c�uχϙ� ������������)� ;�M�_�qߘߕߧ߹� ��������%�7�^� [�m��������� ����$�!�3�E�W�i� {��������������� /ASew� ������ +=Ovs��� ����//</9/ K/]/o/�/�/�/�/�/ �/?�/?#?5?G?Y? k?}?�?�?�?�?�?�?��?OO)�PRG_�COUNT8v�8k�GuKBENB��FE�MpC:t}O_UPD� 1�{T  
4Or�O�O�O__ !_3_\_W_i_{_�_�_ �_�_�_�_�_o4o/o AoSo|owo�o�o�o�o �o�o+TO as������ ��,�'�9�K�t�o� ��������ɏۏ��� �#�L�G�Y�k����� ����ܟן���$�� 1�C�l�g�y������� ��ӯ����	��D�?� Q�c���������ԿϿ ����)�;�d�_��q�=L_INFO {1�E�@ �2@����������� �ٽ`y*�d�h'��¬��=`y;MYSDEBUGU@ʶ@���d�If�SP�_PASSUEB�?x�LOG  *���C��*ؑ��  ��A��U�D1:\�ԘΥ�_MPC�ݵE&�8�A���V� �A�SAV !������ҶX���SVZ�T�EM_TIME �1"���@ 0/  cX��ч�������$T1SV�GUNS�@VE'��E��ASK_OPTIONU@�E�A:�A+�_DI��qO�G�BC2_GRP� 2#�I�����@�  C���<Ko�?CFG %z���� �����` ��	�.>dO� s������� *N9r]�� �����/�8/#/\/n/v$Y,�/Z/ �/�/H/�/?�/'?? K?]�k?=�@0s?�?�? �?�?�?�?O�?OO )O_OMO�OqO�O�O�O �O�O_�O%__I_7_ m_[_}__�_�_�X�  �_�_oo/o�_SoAo co�owo�o�o�o�o�o �o=+MOa �������� �9�'�]�K���o��� ������ɏ���#��_ ;�M�k�}�������� ß�ן��1���U� C�y�g����������� ����	�?�-�c�Q� s����������Ͽ� ���)�_�Mσ�9� �ϭ�������m��� #�I�7�m�ߑ�_ߵ� ������������!� W�E�{�i������ ��������A�/�e� S�u�w����������� ��+=O��sa ������� 9']Kmo� ������#// 3/Y/G/}/k/�/�/�/ �/�/�/�/??C?�� [?m?�?�?�?-?�?�? �?	O�?-O?OQOOuO cO�O�O�O�O�O�O�O __;_)___M_�_q_ �_�_�_�_�_o�_%o o5o7oIoomo�oY? �o�o�o�o�o3! CiW���� �����-�/�A� w�e����������я ���=�+�a�O��� s�������ߟ͟��o �-�K�]�o�ퟓ������ɯ���צ��$�TBCSG_GR�P 2&ץ��  �� 
 ?�  6� H�2�l�V���z���ƿ��������(�_d�E+�?��	 HC���>Ǚ��G����C��  A�.�e�q�C;��>ǳ33��SƑ/]϶�Y��=Ȑ� ?C\  Bȹ��{B���>����,P���B�Y�z��L�H�0�$����J�\�n�����@�Ҿ�� �������=�Z�%�7���?3������	V3.00~.�	cr35��	*����
��������� 3��4��   {�CT��v�}��J2�)�������CFG [+ץ'� *�V�����I����.<
� <bM�q��� ����(L7 p[����� �/�6/!/Z/E/W/ �/{/�/�/�/�/.�H� �/??�/L?7?\?�? m?�?�?�?�?�? OO $O�?HO3OlOWO|O�O ����Oӯ�O�O�O!_ _E_3_i_W_�_{_�_ �_�_�_�_o�_/oo ?oAoSo�owo�o�o�o �o�o�o+O= s�E���Y�� ���9�'�]�K�m� ������u�Ǐɏۏ� ��5�G�Y�k�%���}� ����ßşן���1� �U�C�y�g������� ӯ������	�+�-� ?�u�c���������� Ͽ���/�A�S��� ��qϓϕϧ������ ��%�7�I�[���m� �ߑ߳������߷�� 3�!�W�E�{�i��� �����������A� /�e�S�u��������� ������+a O�s��e��� ��'K9o] ������� #//G/5/k/}/�/�/ [/�/�/�/�/�/?? C?1?g?U?�?y?�?�? �?�?�?	O�?-OOQO ?OaO�OuO�O�O�O�O �O�O___M_�e_ w_�_3_�_�_�_�_�_ oo7o%o[omoo�o Oo�o�o�o�o�o! 3�o�oiW�{� ������/�� S�A�w�e�������я �������=�+�M� s�a���������ߟ� �_	���_ן]�K��� o�������ۯɯ��� #���Y�G�}�k��� ��ſ׿������� �U�C�y�gϝϋ��� ���������	�?�-� c�Q�s�u߇߽߫��� �����)��9�_�M� ����/����i���� ��%��I�7�m�[��� ���������������� EWi{5�� ������A /eS�w��� ��/�+//O/=/ _/a/s/�/�/�/�/�/ �/?'?��??Q?c?? �?�?�?�?�?�?�?O �?5OGOYOkO)O�O}Op�O�O�O�N  �@�S V_R��$TBJOP_G�RP 2,�E��  ?��V	-R4S.;\=��@|u0{S~PU >��U�T @�@LR	� �C� �Vf?  C���ULQ�LQ>�33�U�R�����U�Y?�@=��ZC��P�����R��P  Bȸ�W$o/gC��@g��dDb�^�㙚eeao�P&ff~�e=�7LC/kFaB o�o�P��P��efb-C�p�B�^g`�d�o�PL�P�t<�eVC\ � �Q@�'p�`��  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�anaaF`C�;�`L�w��aQoxp�x�p:���XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb����X �	��1��)�W��� c������������ 󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSc7r35QT*�QT��A�� E��'E�i�F�V#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG��G#
�D���E'
E�MKE���E��ɑE�ۘE���E���F���F��F���F(��F�5��FB��F�O��F\��F�i��Fv��F���vF�u�<#�
<t����ٵ=�_��V �R�p�V9�~ ]ESTPARtp��HFP*SHR\�A�BLE 1/;[$%�SG�� �W�
G�G�G� WQG�	G�
G�GȖ�QG�G�G�ܱv�'RDI~�EQ�ϧ� ��������W�O_�q�@{ߍߟ߱���w�S]�CS !ڄ������ ������&�8�J�\� n������������� ] \�`��	��(�:� ����
��.�@�w��NUM  �EUEQ�P	P ۰�ܰw�_CFG �0��)r-PIMEBF_TTb��CSo�,VERڳ-B�,R 11;[' 8��R�@� �@&  ��� ����//)/;/ M/_/q/�/�/�/�/�/ ?�/?J?%?7?M?[? m?>�@�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_��_l_�Y@c�Y�MI_CHAN�8 c cDBGLV��:cX�	`�ETHERAD �?f�\`���?�_uo�oQ�	`RO�UTV!	
!��d�o�lSNMAS�KQhcba255.uߣ'9ߣY��OOLOFS_D�Ib��U;iORQCTRL 2		�Ϸ~T��� ��#�5�G�Y�k�}� ������ŏ׏�����.��R�V�PE_�DETAI/h|zP�GL_CONFI�G 8�	����/cell/$�CID$/grp1V�̟ޟ�������o?�Q�c�u����� (���ϯ������ ;�M�_�q�����$�6� ˿ݿ���%ϴ�I� [�m�ϑϣ�2����� �����!߰���W�i� {ߍߟ߱�%}F��� ����/�A�C�i�H�Eߞ�������� ��?��.�@�R�d�v� ������������� ��*<N`r� ������& 8J\n��!� ����/�4/F/ X/j/|/�//�/�/�/ �/�/??�/B?T?f? x?�?�?+?�?�?�?�? OO�?>OPObOtO�O��O�O���Us�er View ���}}1234567890�O�O�O�_#_5_=T�P��]_���I2�I:O�_�_�_@�_�_�_X_j_�B3�_ GoYoko}o�o�o o�op^46o�o1CU�ovp^5�o������	�h*�p^6 �c�u����������ޏp^7R��)�;�M� _�q�Џ��p^8�˟ ݟ���%���F�L�� lCamera�J���� ����ӯ���E~�� !�3��OM�_�q��������y  e��Yz��� 	��-�?�Q���uχ� ��俽���������>��e�5i��c�u߇� �߽߫�d������P� )�;�M�_�q��*�<� �i���������)� ��M�_�q�������� ��������<�û��= Oas��>��� �*'9K] f�Q������ �/�%/7/I/�m/ /�/�/�/�/n<�� ^/?%?7?I?[?m?/ �?�?�? ?�?�?�?O !O3O�/<׹��?O�O �O�O�O�O�?�O_!_ lOE_W_i_{_�_�_FOXG9+_�_�_oo(o :o�OKopo�o)_�o�o@�o�o�o ��	g�0�oM_q��� No����o�%�7� I�[�m�&l�n�� Ə؏���� ��D� V�h���������ԟ 柍�g�ڻ}�2�D�V� h�z���3���¯ԯ� ��
��.�@�R���3u F�鯞���¿Կ��� ���.�@ϋ�d�vψ� �ϬϾ�e�w���U�
� �.�@�R�d�ψߚ� ������������*� ��w���v���� ����w�����c�<� N�`�r�����=�w�� -�����*<�� `r�������x���  �� 1CUgy��������    -/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_�i_�  
��( � �%( 	 y_�_�_�_�_�_�_ o	o+o-o?ouoco�o�o�o�Z* � Q&�J\n ������o��� 9�(�:�L�^�p�� �������܏� �� $�6�}�Z�l�~�ŏ�� ��Ɵ؟���C�U�2� D�V���z�������¯ ԯ���
��c�@�R� d�v�����᯾�п� )���*�<�N�`ϧ� ���ϨϺ������� �&�8��\�n߀��� �߶���������E�"� 4�F��j�|���� ��������e�B� T�f�x����������� ��+�,>Pb ���������� (o�^p� ������ /G $/6/H/�l/~/�/�/ �/�//�/�/?U/2?�D?V?h?z?�?�/�`@� �2�?�?�?�3��7�P��!frh�:\tpgl\r�obots\m2�0ia\cr35?ia.xml�?;O MO_OqO�O�O�O�O�O�O�O ���O_(_ :_L_^_p_�_�_�_�_ �_�_�O�_o$o6oHo Zolo~o�o�o�o�o�o �_�o 2DVh z������o� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟�ݟ��&�8� J�\�n���������ȯ ߟٯ���"�4�F�X� j�|�������Ŀ־�8�.1 �?@8?8�?�ֻ� ֿ�3�5�G�iϓ�}� ���ϳ��������5߀�A�k�U�wߡ߿���$TPGL_OUTPUT ;�!��! �� ������,�>�P�b� t����������� ��(�:�L�^�p������������2345678901�� �������"�� BTfx��4�@����
}$ L^p��,>� �� //$/�2/Z/ l/~/�/�/:/�/�/�/ �/? ?�/�/V?h?z? �?�?�?H?�?�?�?
O O.O�?<OdOvO�O�O �ODOVO�O�O__*_ <_�OJ_r_�_�_�_�_ R_�_�_oo&o8o�_ �_no�o�o�o�o�o`o �o�o"4F�oT�|����\��} �����0�B�T�e��@������� ( 	 ��Џ��� ���<�*�L�N�`� ��������ޟ̟�� �8�&�\�J���n��� ������ȯ���"�������*�X�j�F��� ��|�¿Կ��C���� ��3�E�#�i�{�忇� ��S����������/� ��S�e�߉ߛ�y߿� ��;�������=�O� -�s���ߩ��]��� �����'����]�o� �����������E��� ��5G%W}�� ����g��� 1�Ug	w�{ ��=O	//�?/ Q///u/�/��/�/_/ �/�/�/�/)?;?�/_? q??�?�?�?�?�?G? �?O�?OIO[O9OO �O�?�O�OiO�O�O�O !_3_�O_i_{__�_�_�_�_�_�R�$T�POFF_LIM� >�op:�y�mqbN_SV`�  l�jP_�MON <6�)dopop2l�a�STRTCHK �=6�f� bVTCOMPAT-h��afVWVAR �>Mm�h1d ��o �oop`b�a_DEFPRO�G %|j%R�OB195_SE�RV	�j_DIS�PLAY`|n"rI�NST_MSK � t| ^zINqUGp�odtLCK�|�}{QUICKMEyN�dtSCRE�p�6��btpscdt�q��b*��_.�ST�jiRA�CE_CFG U?Mi�d`	�d�
?�u�HNL �2@|i����k  r͏ߏ���'�9��K�]�w�ITEM �2A�� �%$�12345678�90����  =<�П��  !���p��=��c�� ^����������.� ��R��v�"�H�ί�� Я������*�ֿ�� �r�2ϖ�����4�޿ �ϰ���&���J�\�n� ��@ߤ�d�v��ς��� ���4���X��*�� @�����ߨ��� ����T���x���� ��l��������,�>� P�������FX��d ������:� p"��o��� ��F6HZt~ ��N/t/�/��//  /2/�/V/?(?:?�/ F?�/�/�/j?�??�? �?R?�?v?�?QO�?lO �?�O�OO�O*O|O_ `O _�O0_V_h_�Ot_ �O__�_8_�_
oo �_@o�_�_�_Lodo�_ �o�o4o�oXojo3�o N�or��o���s�S�B���zψ  h��z 8��C�:y
 P�v��]����UD1:�\�����qR_G�RP 1C��?� 	 @Cp� ��$��H�6�l�Z��|�����f���˟��<�ڕ?�  
�� �<�*�`�N���r��� ����ޯ̯��&��0J�8�Z���	�u������sSCB 2D� ����π(�:�L�^�pς��|V�_CONFIG E���@����ϖ��OUTPUT yF������� 6�H�Z�l�~ߐߢߴ� �����������#�6� H�Z�l�~������ ��������2�D�V� h�z������������� ��
�.@Rdv ������� )<N`r�� �����//% 8/J/\/n/�/�/�/�/ �/�/�/�/?!/4?F? X?j?|?�?�?�?�?�? �?�?OO/?BOTOfO xO�O�O�O�O�O�O�O __+O>_P_b_t_�_ �_�_�_�_�_�_oo '_:oLo^opo�o�o�o �o�o�o�o $�� ��!�bt���� �����(�:�-o ^�p���������ʏ܏ � ��$�6�G�Z�l� ~�������Ɵ؟��� � �2�D�U�h�z��� ����¯ԯ���
�� .�@�Q�d�v������� ��п�����*�<� M�`�rτϖϨϺ��� ������&�8�J�[� n߀ߒߤ߶������� ���"�4�F�W�j�|� ������������� �0�B�S�f�x����� ����������, >Pa�t���� ���(:L>/x���k} gV�K���/ /&/8/J/\/n/�/�/ �/W�/�/�/�/?"? 4?F?X?j?|?�?�?�? �/�?�?�?OO0OBO TOfOxO�O�O�O�?�O �O�O__,_>_P_b_ t_�_�_�_�O�_�_�_ oo(o:oLo^opo�o �o�o�o�_�o�o  $6HZl~�� ��o���� �2� D�V�h�z�������� ԏ���
��.�@�R� d�v���������Ϗ� ����*�<�N�`�r� ��������˟ޯ�� �&�8�J�\�n����������Ż�$TX_�SCREEN 1}Gg��}ipnl/���gen.htm�ſ�*�<�N�`Ͻ�Panel soetupd�}�d�@�Ϸ����������� ��6�H�Z�l�~ߐ�� ��+�������� �2� �߻�h�z������ 9�g�]�
��.�@�R� d������������� ��}���<N`r ��;1�� &8�\��������QȾUA�LRM_MSG k?��� � Ȫ-/?/p/c/�/�/�/ �/�/�/�/??6?)?�Z?%SEV  �-�6"ECFoG I���  ȥ@�  }A�1   B�Ȥ
 [?ϣ��?O O%O7OIO[OmOO�O��O�G�1GRP 2�J�; 0Ȧ	 ��?�O I_BB�L_NOTE �K�:T��#lϢ�ѡ�0R�DEFPRO %+ (%N?u_Ѡ c_�_�_�_�_�_�_o �_o>o)oboMo�o\�INUSER  �R]�O�oI_ME�NHIST 1L��9  (_P� ��)/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,1133,1�oDVLhz~�(
50�������zed;it(rONE�I��[�m���	#�OP�EN8�Ώ���� 3�'���~71��P��b�t����0���R�OB195t0RV�?�ݟ����� z37̟X�j�|����/�)r95G�ݯ��� 6Q�`q|oB�T�f�x� ������1�ƿؿ��� � ϯ�D�V�h�zό� ��-���������
�� �Ͻ�R�d�v߈ߚ߬� ;���������*�� N�`�r����7�I� ������&�8�#�\� n��������������� ��"4F��j| ����S�� 0BT�x�� ���a�//,/ >/P/�t/�/�/�/�/ �/�/o/??(?:?L? ^?I��?�?�?�?�?�? �?�/O$O6OHOZOlO �?�O�O�O�O�O�OyO _ _2_D_V_h_z_	_ �_�_�_�_�_�_�_o .o@oRodovoo�o�o �o�o�o�o�o*< N`r�o?�� ����8�J�\� n�����!���ȏڏ� �������F�X�j�|� ����/�ğ֟���� ���B�T�f�x����� +�=�ү�����,� ��P�b�t��������z��$UI_PAN�EDATA 1N����ڱ�  	�} � frh/cgt�p/widedev.stm���%��7�I�Y�)  ri ρ�@�밙ϫϽ��� ����Z��)��M�4� q߃�jߧߎ������߀���%�7��[�7��� �     H�d�� ����������E�� ��:�L�^�p������� ����������$ H/l~e������o�ܳ7� <N`r���� -���//&/8/� \/n/U/�/y/�/�/�/ �/�/?�/4?F?-?j? Q?�?�?%�?�?�? OO0O�?TO�xO�O �O�O�O�O�OKO_�O ,__P_b_I_�_m_�_ �_�_�_�_oo�_:o �?�?po�o�o�o�o�o o�o sO$6HZ l~�o����� �� �2��V�=�z� ��s�����ԏGoYo �.�@�R�d�v�ɏ�� ��П������ <�N�5�r�Y������� ̯���ׯ�&��J� 1�n�������ȿڿ ����c�4ϧ�X�j� |ώϠϲ���+����� ���0�B�)�f�Mߊ� �߃��ߧ�������� ����P�b�t���� ������S���(�:� L�^����i������� ���� ��6Z�lS�w�'�9�}���"4FX)�}��l��� ��/j'//K/2/ D/�/h/�/�/�/�/�/ �/�/#?5??Y?��C��=��$UI_PO�STYPE  �C�� 	� e?�?�2QUI�CKMEN  �;�?�?�0RESTORE 1OC��  �L?��6OCC1O��maO�O�O�O�O�O uO�O__,_>_�Ob_ t_�_�_�_UO�_�_�_ M_o(o:oLo^oo�o �o�o�o�o�oo  $6H�_Ugy�o ������ �2� D�V�h�������� ԏ����w�)�R� d�v�����=���П� �����*�<�N�`�r� �������ޯ�� �&�ɯJ�\�n����� ��G�ȿڿ�����7oSCRE�0?�=u1sc+@Wu2K�3K�4K�U5K�6K�7K�8K��2USER-�2�D�SksMì�3��4��U5��6��7��8����0NDO_CFG� P�;� ��0P�DATE ���None�2���_INFO 1eQC�@��10%� [���Iߊ�m߮��ߣ� ���������>�P�3��t��i���<-�OFFSET T�=�ﲳ$@������ 1�^�U�g��������� ��������$-Z@Qcu���?�
�����UFRAME�  ����*�R�TOL_ABRT8	(�!ENB*?GRP 1UI�1Cz  A�� ~��~�����!���0UJ�~9MSK  M�@�;N%8�%x��/�2VCCM�³V�ͣ#RG�#Y��9���/����D��BH�p71Ce���3711?�C06�$MRf2_�*S��Ҵ�	���~XC56 *�?d�6���1$�5��m�A@3C��.' ��8�?���OOKOx1FOsO�5��51��_O�O��? B����A2 �DWO�O7O_�O8_#_ \_G_�_k_}_�__�_ �_�_�_"o�OFoXo�%TCC�#`mI1�i������� GF�S��2aZ; ��| 2345678901�o�b���� �o��!5a�4Bw�B�`56 311:�o=L�Br5v1�1 ~1�2��}/��o�a� �#�GYk}� p�������ُ� 1�C�U�6�H���5�~� ��ߏ���	���4�dSELEC)M!v1�b3�VIRTS7YNC�� ����%�SIONTMOiU������F���#bֳ����(u FRk:\H�\�A\��� �� MCLOG��   oUD1��EX�����' B@ ����̡m��̡_  OBCL�1��H� �  =�	 1- n?6  -�������[�,S�A�`=�̩͗��ˢ��TRAIN⯞b�a1�l�
0d�$j�T2cZ; (aE2ϖ� i��;�)�_�M�g�q� �ϕϧ��������	���F�STAT 	dm~2@�zߌ�*jq$i߾��_GE�#�eZ;�`0�
�� 02��HOMI�N� f־��ֿ ~�����БC��g�X���JMPE�RR 2gZ;
  ��*jl�V�7��� ������������
��@2�@�q�d�v�B�_ߠ�RE� hWޠ$LE�X��iZ;�a1-e���VMPHASE'  5��c&��!�OFF/�F�P2*n�j�0�㜳E1@��0ϒE1!1�?s33�����a k/�kxk䜣!W�m[�䦲�[���p�o3;�  [i{��� �/�O�?/M/ _/q/��/��//�/ '/9/�/=?7?I?s?�/ �?�/�/�?�??Om? O%O3OEO�?�?�O�? �O�O�?�O�O�O__ gO\_�OE_�O�_�O�O /_�_�_�_oQ_Fou_ �_|o�o�_�oo�o�o �o�o;oMo?qof- �oI����� 7�[P����� ����ˏ��!�3�(� :�i�[�ŏg�}�������TD_FILTuEW�n�� �ֲ:���@���+�=� O�a�s��������� ֯�����0�B�T��f�x���SHIFTMENU 1o[�<��%��ֿ���� ڿ����I� �2�� V�hώ��Ϟϰ��������3�
�	LIV�E/SNAP'�?vsfliv��E�����ION �* Ub�h�menu ~߃�����ߣ���p���	����E�.�50�s�P�@j� ��AɠB8z��z��}��x�~�P�� ���KMEb���<�0���MO��q����z�WAITDI/NEND�������OK1�OUT����SD��TIM.����o�G��� #���C���b������RELEASE�������TM�������_ACT[������_DATA 	r��%L����x�RDISb�E��$XVR�s����$ZABC_GR�P 1t�Q�,�#�0�2���ZIP�u'�&�����[MPCF_G' 1v�Q�0�/�� w�ɤ�� 	�Z/  8�5�/�/H/�/l$?��+�/�/�/?�/�/�???r?�?  �D0�?�?�?�?�?�;����x�]hY�LIND֑y�� ��� ,(  *VOgM.�SO�OwO�O�M i?�O�O^ PO1_�OU_<_N_�_�O �_�_�__�_�_x_-o oQo8o�_�o�oY&#s2z� �� �oC�e?a?>N|�o�q����qA�$DS�PHERE 2{6M��_�;o��� !�io|W�i��_��,� �Ï���Ώ@��/� v���e�؏��p�����`�����ZZ�� �N