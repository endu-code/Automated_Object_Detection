��   ,��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2R �$�$CLASS  �������Pz��P� VERS?��  ��5�IRTUAqL��' 2 ��P @ e����  B� ��� K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{����������_C_CCL� ?��  �	All pa�ram��
Ba�se!�Pos�./Speed �checkF�Sa�fe I/O c�onnect�}R���,�>�P�b�t�SEI��@���� � ,�>�g�b�t������� ��Ο�����?�:� L�^���������ϯʯ ܯ���$�6�_�Z� l�~�������ƿ�� ���7�2�D�V��z� �Ϟ����������
� �.�W�R�d�vߟߚ� �߾��������/�*� <�N�w�r������������O���� C�l�g�y��������� ������	D?Q c������� �);d_q �������/ /</7/I/[/�//�/ �/�/�/�/�/??!? 3?\?W?i?{?�?�?�? �?�?�?�?O4O/OAO SO|OwO�O�O�O�O�O��O__�N�   7�_b_�_�_�_�_�_ �_�_�_oo(o:oco ^opo�o�o�o�o�o�o �o ;6HZ� ~�������0� �+_�SI��6� F�;�}�������ŏҏ �����,�>�U�b� t���������Ο�� ��-�:�L�^�u��� ������ʯܯ��� $�6�M�Z�l�~����� ��ƿݿ����%�2� D�V�m�zόϞϵ��� ������
��.�E�R� d�vߍߚ߬߾����߀����*�<�G�Y�P�C_6�SFDI1$N��2���3���I4���5���6����7���8-�e�Q� c�u������������� ��);Mdq ������� %<I[m�� ������/!/ 3/E/\/i/{/�/�/�/ �/�/�/�/??4?A? S?e?|?�?�?�?�?�? �?�?OO+O=OTOaO$l�~�O���O��C ��C��C��C��C ��C,��CD�@�o_�_ �_�_�_�_�_�_�_o :o5oGoYo�o}o�o�o �o�o�o�o1 ZUgy���� ���	�2�-�?�Q� z�u�������Ϗ� 
���)�R�M�_�q� ���������ݟ�� *�%�7�I�r�m���O�}�S���BVOF�F��FENCE~ۯEXEMG�|���NTED"��OP�2�AU;TO:�T�Oy�<�O�MCC��3��CSBP�����O�@}�ׯ ����t����DIS��OC_6�²_~�qė� 