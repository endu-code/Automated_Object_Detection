��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk" 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&�B4��_sC3���r7�"�A_p�d`U��@VA}DCMVROU
b��1PERIO�sF31P���2D-��32%T��1_D��2H�ĺ3��T����K�95K��K�7CL����0�ADJ����_Uvdr[PAUX�@��	 4�@C�P?a$� A�&�n@� qUX_AXS>� \
LD��� 
 h �D�rӠ�Cd��C�t�C �F�@�H�G1P�FOXp4�XAXISU� Tj��D͡�q�E��yAP@M@ 	BQ܀HR
$IDX\PRVڹQSa�GRT��L $F�E_�Uנ���TTOOL�R�p;�A��p�y1;DOf` \��0�R_PKG�RQ= BQ NR�P�BQS�P[Q #2	hQ�P�S�P�2�Q�Qba�	�1ad�o$VFLw0IM�,�LT�r�:a��Tc��6Tb����$DIYG��C$d0JgGUg	�d�4�d�cMPSWP�  �$ @�� � ����a �  &�` &�`V�ERSION�h�I@�5�aIRTUAL�o�avS�?�h&�  �aL|J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x��a+u|P�11 29{q\�`I@�� ֓�Ә��  ?�a @�`����A�  �����#�����3��-�?�Q�?��g�U����  D�  Bp  =���Ϳ�?333C?�a�̠�̤@��vߥA ��/  &� G�P ?ff=fˡ>��ߥ�� �����0�ܙD���̤ ˡ��k�C�Z�[���`�0�����ӿٲ��B�ђǟI�ÿ��<;���F@ K���������Dz��l�W� I��ٺ��ܑ�P`B��w���ēV��'� 9�K�]�o�5ߓ���_� q�ۿ�������#� 9�G�y�7�I�j�߳� ����������a��!���y�3����ϋ� 9�K�]�oρϓϙ��� x���D���������� �,>�b��`����� ������ɤ����� ��Đؓ���2/d����L����^/\�Ϣ�@]�ĐW��"�`�"��'B���������/"  $đƚ�$1>!B,4_��(����1?��?�?�8>��� �ā�//@/�?T/f/ ?O�/�/�/�/�/�/�O ??,?>?P?b?;_�? __�?�?�?�?�?OO (O�_o^OpO�O�O�O �O�O�O�O __$_�o H_Z_3~_�W��fx���2�����$	���o2�2-�V� h�z�������ԏ� �������Dqdd���� �l��ߩߩ�b�����o�����ğ���cd��p(������qT�@� a>Ho�
}��[��c|�>LŠ���_v����<#�
�Qsbp�|��X��o�C��� a?e?a��3�T`��@ �G_�
�T���_����x�2bo%{B ta�������1��U�g�k�`>X�ؤ�����ϑ�It$ ��$�$�>�٢
���A���߭�'�����4�+����s�.����Ճa$敕��(�4$ܛ�S�e�;�{�.��>��H��ރa5����8M�Y��;�=���3��a�B�	9�R�=�v� a�ߡ�����������m����  �b\'������`k� S�K�X�,�w�������P/�����C��Q�??333;�s�<�|�saD/  C``�G�P ?fff/a>$���?_	W�_ ��0��_g�;�5c ?�4'e��xu�j� F@ �0�[�� DzI ����w5���y ܃�����/ ���/�/7I�_I/ [/m//�/�/�/�?�? �?�/?!?3?E?W?i?�{?�?kO}O�?�?�L� Oq�O����� ��O���O�O�_
__ ._@_R_d_o�_�_,o �_o�_�_oobo%�`&/ $.(� �?��>�"��o���� }��o��E+̰�B�� +��ȴC��8����� {j4�~gĠ{t��"�� �����$�3t7�q�x����>���3t �cu����� �����)�W���_� q�����������ݏ� ȯ�%�7�I�k�%�� ��j���ǟٟ��� Ϳ3�E�W�i�{�a��� ����կ�L�o0��������2Q/�A�S�e�v�Uώ�2�߲��� ��������0�B�T� [Ru��������� 7M;	;	/�DO*GT�V@� �M�D�i���Op@�����Ѱ����A>�a��f��B�BH���>L! H���g�O<#�
�ϲp���w�E�v�������A��7������@ \A�b�f��D?B,�@�7J���_���Bб ���Z{�p��N���>�4_�U�/^��It$ //$��K>�5
/a'A���a/	/�/-/?&��+�{���%.����%ޏ�$敕�%(4�$��%�/�+;��=.#5>��H/5���5��?58M�	YK5��= g5��8�x?�+	�/�?�?�?�7 ?�?O$O6OHOZO��o�GnlG   ;¸`�X���E�E ��A��O�O�O	_�2( _^����`=�e?333���B�����D/  C��G�P ?fff��>���e�Y�Q�i� �OVb�m����W�i� ]ooo�o��k��_wo�o<�`F@ uawU�`Dz�P$to��o�j"���� ��_�_oo'o�Ko U�)��o�oﯥ� ����1���"� Y�k�}�������ŏ׏@�ǟٟX�1��̸k� �oC��o'9K Q���0�B���f�x��� ������z������� l�>�P�b�t���lu��`�\�nπϊx�O� ������4����� C�<���R(���� c�$�C� ���׺ ��ڷ  �Ę�~Jk���_V�؏��/�?�<Q�]�>�����]� ����������+�� O�a�s߅߳�U����� ��������9�K�$ o���������� ��#�5�G�u�k�) ������������� �1ǼZό�/0/B/X%2�l�/�/�/�/�-	��"2�/? ?2? D?V?h?z?�?�?�?�d �n�>�GYGZ<�� �Y�Y�������ijO |O�O�O�FK �G�LO^Ib!W�#�>� �'_����4U�>L}PdQ�.B�<'#�
K+p4_�Bp�t�FB���@��SU�RkU@�� lT��o�δ���ζ ��0o��eB,TU Po�o�o�o�o��P>a�T�O�OrIC�It$ �$�&>%��R
k�wAHD��e���v�@+��=�+�.���7��A�$敕G�(4$��S���;��.��>��H���A5�����8M�Y���==dPÅ�B�ԏ�{	�
���.��g� Y�n���������%o�=|��ȗ  B ��R�T_b�P#��J ��X/�A�S�e��|��j�B�	��S��?333�E+��D7Ica�D/  CGÿP ?fff�A> �Q8D����O=X� ���M�O���o�� ˿���?Y�ӿ-�Kl�F@ _�k�ӥbl�Dz���k�]��/��~!^/P) � ;�M�_�q���Iߧ��� s߅���K��%� 7�M�[ߍ�K�]�~�� ���������!�3�u� #�5����Sl���)� ��M�_�qσϕϧϭ� GR����X�������� 
�@R�v� ������/��0�����ȫ��  viڗ�N.k_=C� �/o�㢄`s���U�" �d�Q�f�PcEci3�/ 6|P3$�ښ�$E>�Us��(��)o�<�?�8>�����:/ -/?/Q/c/u/�/`O�/ �/�/�/?�O?)?;? M?_?q?J_�?�?�_�? �?�?O#O�_7OIO"o mOO�O�O�O�O�o�O �O_!_3_oW_i_B �_{���z���u�2	�����.�F�2A�j�|����� ��ď֏�����
� -�Xqxd�����l��� ��b�����Ɵ؟���!�wd�p<���P���qh�T�_a>\���}z�o� s��>�L٠�� o��y<#�
�Q�bp��/�l�8�o.�c���_aSe Wa��G�h`ǥ@�Ȥ [s��T���_�V����Fbo9{B�a���� �3�E�(�i�{�.k��>l�����ϥ�I�t$ ��$8�>��
���A������;�����H�+��̞��.�����G�$�敕��(4$�x��g�y�;��.���>��H��G�5{����8M�Y�O�=���G��a0�V�	M�f�Q��u��ߵ� ������ ����'��>$�  �bp ;������g�_�l� @���������C������c��e��S?3�33O���P���ñD�/  Ct`G�P_ ?fffO�>8� ��Ss	k�_!xD� s{�O�IwS�' H;e#��/��j� F@ ��/o�� Dz] ����pI�q��y ܗ �����//�/ �/K]�_]/o/�/�/ �/�/�/�?�?�??#? 5?G?Y?k?}?�?�?O�OO�?g|�#O��O �����/	_�� �O�O�__0_B_T_f_ x_2o�_�_@o�_$o�_ oo,ovo$%t:/&8B(�OPp\c ҹ6��o�~ǯ���o� �E?��BPp?��ܴ W���L������jH��g ؠ�tPq6�#������8�GtK߅���	��>���Gt�w� ��������� +�=�k��s������� ��͏����ܯ'�9� K�]��9�����~�ɟ ۟���-�#��G�Y� k�}���u���ů��鯀lD�������2@eC�U�g�yߊ�i���2�����������  �2�D�V�h�of�� ��Դ������KMO	O	 C�XO>Gh�j"�4�a�X�}�ӴИ���(�����p�>�a���z��B�B\���>L�5 \���{�<#�	
��p�����E,�������p������İ#@pA$�b �z�B�SB@�KJ���s���B�n��������t >��Hs�i�*/�Itk$ C/$��>�I	
#/u'A �u//�/xA/S&��+����%�.����%��$�{���%(4$�5��/�+;��.75>���HC5��5�=�S58M�Y_5��= {5��L��?�+	 �/�?�?�?�7?O&O�8OJO\OnO}K�$C�CSCH_GRP�12 2�����A&� �\��Xo��  O��`�l t �E�E���A�__@,_>_�2U_C^����`yQ�e?333���R����#D/  �CаG�P ?fff��>���e�Y �Q�}��Ojb�m��� �W�i��o�o�o����2o�o�E`F@� 8uDa�U�E`Dz �PYtDo6�j6��� �o&o8oJo \o"��o�L�^��o�o �����&�4�f� $�6�W�������ď֏ ����N������f����x�&8J \n�����e�w�1� ������ѯ������ +���O���s������� �u�Ϸ�ϣϵϿxȄ���ٳ.��i� '�#��x�q�H��R< L������8�W�  �����4 �����J���sLV�����/�t���>����Ē�����*�<� N�`�9��ߖߨߺ��� ������&�8�J�# n��Y��������� ��"��F�X�j�|� ����^�������� �0B/f�����S/e/w/�%2�l�/�/H�/�/=�22? C?U?g?y?�?�?�?�? �?�?�d�nN1!Q|Y |Zqȝ�Y�Y�՟�� ��i�O�O�O�O�FP� W�O�I�!AW-3�>5�\_�S�H��iU>L�P�Q�<cB�<#�
�`�pi_RE��V<B���,0�U bA�U@푡T4�Lo�� В�fȚeo��Ba�U�o�oBT�P>Ea�T�Ox�O�~CIt$ �-$6>��R
��wA}D�����v!P�+���`�.��y�l� Q$敕|��(4$܈�@�R�;���.��>��H��� Q5��Ѕ8'M�Y܅(M=�P�� R�	�/�	&�?�*� c�N���������ǟٟ��Zo Mؾ��  �I�b�T�b�P X�@�8JE�hd�v�����������<B�>�<�S,�?333(U`��)TlI�aD/  C�MG�P ?fff(Q>amD,�L�D� ����L�TM(_"� P�,� �!��?����bπ��F@ `�Š��Hb��Dz6� �Ġ���d�"ʳ!�/�) �p��������� ~�ܿ�Ϩߺ�$�6π 6�H�Z�l߂ߐ��߀� �������� �2�D� V�h��X�j���������^����ϔϦϸ� ������|R������� 	-?Qu� �����O���M/���/����) 5�i���. �_nC��/����`�� ) e�"�d0a�f%`�E �ih!?k�Ph$)!�@�$z>�U��8 $$��^o�<�?�8>���  $�:P/b/t/�/�/�/ �/�O�/�/??D?�O L?^?p?�?�?�?_�? �?�_ OO$O6OXOo lO~OWo�O�O�O�O_ �O�o _2_D_V_h_No �_�_w�_l�/����u2>��.�@�$R�c�B{�2v��� ��ÏՏ�����/� A�H�?�b��q�dةت �l$�(�(�r1��A�C����:�1�V��d��pq�ݟ��q����Ia>���S}���5sť>L���5o���Ty<#�
�Q�bp�ůd���c�����Ia�e�a�|��`��@I������Sd,�o۶$���{bLon{B �a��G�h�z�]Ϟ���ckM�>��!�L�B���ړIt$ �$�m�>�"�
��N�A�ٔN���p��,�}�+���̼�.������|�$敕��(�4$��՜߮�;�{�.�>��H��|�5��,�8M�Y8儝=��T�|�%qe��	�ߛ��� ���������#�5�G��\�4Y�  (r�p�E��M��� ������u���������Px�������*��?333����|ș��D/  C�`�G�P ?fff��>m�ɔ��	��_ Vxy�C�����~� ��J\}peX��dx��j� F@ �0�d��� Dz� $����~���y �����/ 8B/??���_�/ �/�/�/�/�/?�?�? OF?X?j?|?�?�?�?��?O�O�OEOO�L� XO�0_��//&/ 8/>_آ_/_�_S_e_ w_�_�_�_go�_�_uo oYo+o=oOoao�oY%��o/I[mw(� <O�p�c�k�!�~�� Γ0)� Ut�R�p t�P�Č�0Ɓ����� �j}��g��t�qk�X� ֎L�m�|t�ߺ�x,�>�J�>���|t J�������� �<�N�`�r���B��� ��̏ޏ���ۯ&�8� �\�n�������n�ȟ ڟ�����"�4�b�X� �|�������į��� �����p�Gy��/�E�2�xߊߜ߮�������2����� �1�C�U�g�y��� ������	�4	4
)� �M�	�	xOsG�ϟ@W�i��������8�@��9�K�O����� Q>�a��R R��!>Lj Q����O<#�
8��p!����EaϿ������ Q��@���X@ �AY�b��w��Bu�@7�Jײ����B� A=�����/��� >�}����_/^6�It$ x/$��K>�~
X/�'A5���/R/�/v/�&��+�{��5.���$5���$敕45(4�$�@5�/
;;��=.l5>��Hx5���5���58M�	Y�5��=Q �5����?�+	�/�?�?OG T?FO[OmOO�O�O���n�G   ��p��L� U�E ���A�_._@_R_�2(i_W^����`��e?333��R��$��XD/  C�G�P ?fff��>�-��ei�Q<��� �O�b}����Wy� �o�o�o̵��Fo�o<8�Y`F@ LuXa�U Y`Dz�PmtXo�J�jk�K�=� �(o:oLo^opo6��o �`�r��o�o8�� � �$�:�H�z�8�J�k� ����Ə؏���� �@b��"���z�4���� ��:L^p�� ��4y���E�����ӯ ���	�ÿ-�?�ѿc� ����������ϵu�`��Ϸ����xȘ� ���c�G}�;�X&� �υ�\��Rq`���� ��m��� P�P � ��#�i  ����J��2��`V�����/��<���>����Ħ� ��,�>�P�b�t�M� �ߪ߼����ߞ��� (�:�L�^�7���m ����������$�6� Z�l�~�������r ������ DV //z�����g/y/�/�%2�l�/�/�/
?=	�322.?W?i?{? �?�?�?�?�?�?�? t �nNE!e�Y�Z�ܝ �Y�Y��ϗ��i�O �O�O�OVd� )W��O�I�!UWA3L>�I�p_-g�\��}U�>L�P�Q�wB)<'#�
�tp}_RpY��VPB��L@@D�U4bU�U@� �TH�`o/����f ܚyo3&+Bu�U �o�o 2Vh`>Ya�T_�O��C�It$ �$%6>%��R
��A�D��(���v5P+��=�t�.�����4Q�$敕��(4$�ܜ�T�f�;��.�ȅ>��Hԅ4Q5����8M�Y��<M=�P�4R��C�	:�S�>�w�b��� ����ɟ۟���noM|��  � ]�(b�T�b`l�T�LJ Y�-hx�������0�ů���PB�R��S@�?333<Ut�=T�I�a�D/  CaGÿP ?fff<Q> %a�D@�`�X��(1� ��`�hM<_6�d�@� �5�(O���vϔ��F@ �Ŵ��\b��DzJ��Ĵ����x�6��!�/�) � ��������̿����� ����8�JϔJ�\�n� �ߖߤ��ߔ������ �"�4�F�X�j�|�� l�~��������r� ���ϨϺ��������� �R�����/A Se��-� ��c�a/'�0//%//����=  I�i#���.�_~C� �/��,��`��= ,e2 �dDa�f9`�E�i|5? �P|$=!#�4�>e��%84$8�ro�<�?H>���4$Jd/ v/�/�/�/�/�/�O�/ ??*?X?�O`?r?�? �?�?�?�_�?�?�_O &O8OJOlO&o�O�Oko �O�O�O�O__�o4_ F_X_j_|_bo�_�_� �_(l�1/����u�2R�0�B�T�f�w�V��2����ŏ׏� ����1�C�U�\�S� v��q�d���l8�<� <�0rE�+�UW��!�N�E�j��d�p���P������]a>��̯g}���Is٥>�L"�	�IoӒhy<#�
�Q�bpٯx���8w�����]a�e �a�����`�@]�� ���g/d@�-o�8�տ�b`o�{B�a���� [�|ώ�qϲ���wka��>��5�`�V���I�t$ 0�$��>�6�
�b�A�b�
����.�@֑�+��̞��.����Ր�$�敕��(4$�x�հ���;��.$��>��H0吡5{��@�8M�YL���=	�h吢9qy��	�߯����������%�7�I�[�j��$�CCSCH_GR�P13 2������&�� \�~E�y  <r���Y� �a������������+��B0����>��?333�����ܙ�D/ � C�`G�P ?fff��>��ᔜ �	��_jx��W�ĝ ���������e�l����j2F�@ %%1���2Dz� F$1#/��#���y �% 7I?mw/9?K?� ��_�/�/�/�/?!? S?O#ODO{?�?�?�? �?�?�?�?;O�O�OzOSO\��O�e_/%/ 7/I/[/m/s_�R_d_ o�_�_�_�_�_�_�o oo�o<o�o`oro�o �o�o�%��/~���(�qO�p�cɠ� V��ޓe^�5U� )�9R�p����%Ġ�D� �����j���g!��t �q�����`�9���t���οa�s��>����t����� )�;�M�&�q������� Տw�ݏ���%�7� �[�m�F�������ǟ 韣�����3�E�W� i�����Kϱ�ïկ� ��߿�/��S���| �@�R�d�z�2��ߐ�����������2 �0�B�T�f�x��� �����������>� i	i
^̵M�	�	���O �G�������������=�m�n�����.
�ڱ>"qI��@R85R��V>L� �xƿP���<#�
m�M�pV��2U����)���ڱ��u.��@�A�!r9�� ���B��l�JR�ݿ��BN�vr��/ �//A/��� >2�������/k�It$ Z�/$��>��
�/�'Aj��/�/?�/�&� +���M5.����Y5$敕i5(4$�u5-??;�;��.�5>��yH�55���5O8M�Y�5�=�  �5���?;	?,O OPO;G�?{O�O�O�O��O�OG���n�G  ��6p�� � EU-U%�2QQ_c_@u_�_	B�_�^)��+py�u?333�MRY��D/  �C:�G�P ?fff>�Z�u9i 1aq���
_�b9}A� g=y/�o�o����{o�oOmʎ`F@� �u�a�U5�`Dz #`�t�oQz�р�r� �]ooo�o�o �ok��o�����# m�#�5�G�Y�o�}��� m����׏����� 1�C�U���E�W�֟��i���K��o�� ���ϯi����z� �����,�>���b� t�Ϙ�꿼�ο�� <��u:� ���������͟�"Ø�G�� pލW��Ϻߑ�b� ����Ң� ���U��XǞ U�р�J��g���V����?K������>������=�O�a�s߅� �ߩ߂��������1� ��9�K�]�o���l ���������#�E� �Y�k�D�������� �����1CU ;y�d/���
��/�/�/�%2+|	??H-???P=//h22c? �?�?�?�?�?�?�?
O O.O5t,~ONz!��Y �Z��ii	"�� ./0y�O�O'__CV�� ^W�O�I�!�Wv3��>~��_@-����"#�U>L�P�Q"<�BA)<#�
���p�_QR���PV�B����uy�Uib��U@6��T}o@/ ��f��oh9[+B��U�o4UgJ��P:`>�ad9_x/_��CIt$ 	�-$Z6>�b
�;�A�D;��]���jP�+��̩�.��y���iQ$敕Ņ�(4$�х����;���.��>��H�	�iQ5���8'M�Y%�qM=�PA�iR!R�x�	o���s� �����ן����"��4��oIM!�F�  "��]b2d�b:` �����J��bh����ѯ��e���讅B���<cu�?333qU���rT�I�aD/  C��G�P ?fffqQ>Za�Duŕ��� �C(f�0͝Mq_k� ��u7�I�j�]EO׿�Qϫ���F@ `���Q��b�Dz� ����ϭ�k��!�/�) ܹ�˿ݿ�� ��%�/����m��� ߑߣߵ�������� ����3�E�W�i�{�� ��������2�����E���������� �%�+�R
�@ Rdv��T�� b�F*<N��FՖ/\�6/H/Z/d��)�r ~�iX�/�. �_�C/?��a�p�� r ae=2�dyavn`�E �i�j?��P�$r!X�@E4�>9e�Z8i$m��oL+O7H>��� i$7J�/�/�/�/�/�/ ?�O)?;?M?_?�?/_ �?�?�?�?�?�?�_O %O�_IO[OmOO�O[o �O�O�o�O�O_!_O_ E_i_{_�_�_�_�o �_�_�o]l4/f/�
��2�2��e�w���$�����Ă2��� ����0�B�T�f�x� ���ĈΫ��q�d!�!� |m�q�q�erz�`�����D�V���z����d�%���&�8�<��҃��>���}����~s�>LW�>�~o���y<#�
%arp������N��������e�a-�Ų�`E�@��F���ddu�bo$�m�
��b�o�{B q.�*ϐϱ��Ϧ����Ϭk��>�j������L�#�It$ e�$���>�k�
Eߗ�A�"���?߹�c�u�Ơ+�����.�����š$敕!�(�4$�-�����;�{�.Y�>��He��š5��u�8M�Y��͝=>���Ţnq����	������� ��A�3�H�Z�l�~��������}��  qr�����9��� ��ݚ��	-?P��VD���s��?333ͥΤ|�E�D/  C�`�G�P ?fff͡>�����	�)o �x������ͯ�� �ϓ���e��3�x/%zFF@ 9%0E��FDz� Z$�E7/	/�X�8�*� �'9K]#? ��/M?_?��%o�/ �/�/?'?5?g?%O7O XO�?�?�?�?�?�?�?�OOO�O_�OgO!\� �O/y_'/9/K/]/o/ �/�_!�f_x_2o�_�_ �_�_�_�_�oo,o�o Po�oto�o�o�o�o�%���/����(� �O�p�cPɴ�j(�E� �yr�IU�^�MR�p ����Z�ձy�ʰ=�=� zƏwV���q���� ���M���t���xu�����>����t �����+�=�O�a� :���������鏋�� ��'�9�K�$�o��� Z�����ɟ۟����� #���G�Y�k�}����� _�ůׯ�����1� C��g�����T�f�xߎ�2������������ �2�D�V� h�z���������� ���2�R�}	}
r� �M�	�	���O�G���@����������Q���@������B.�9�>6q]��TRIR��j>L� �ڿd���O<#�
��a�pj�	FU��=����9�-�1��!B��@ �A�5rM�����B��@��Jf ���Bb� ���///C/U/�� >F������/^�It$ �/$�K>��
�/�'A~���/�/?�/�&" +�{��a5.���m5�!$敕}5(4�$܉5A?S;;��=.�5>��H�5!�5���58M�	Y�5)�=� �5!��
O0;	'?@O+OdOOG �?�O�O�O�O�O�O[���n�G   ��Jp��� YUAU 9�FQe_w_�_�_B(�_�^=��?p�-u?333)aR*m���D/  CN�G�P ?fff)>n�-uMiEa���� _�bM}U�)#gQy-/ �o"���o	c<�ʢ`F@ �u�a	eI�`Dz7`�t�o��e#z�є߆� �qo�o�o�o�o��o �����%7��7�I� [�m�����Ï������ ����!�3�E�W�i�@��Y�k��ß}���� _կ������ �}¯ԯ����
�� .�@�R��v���Ϭ� ��п����P��uN�`��� ����� *�6ìW�τޡk� ���ߥ�b���*� �Ҷ1�&���i� "�lǲ i�*�Z��{���V�!�%?_��<����>���!��� Q�c�u߇ߙ߽߫ߖ� ������E���M�_� q�������� ��%�7�Y�m�� X����������� !3EWiO�� x/���߰/�/�/�%2?|?/?A?S?d=	C/|22w?�?�?�? �?�?�?OO0OBOIt @~cN�!��Y�Z�%� )i)i"2��B/Dy�O _;_2_WV�� rW��O�I�!�W�3J>����_T-����6#�U�>L`�Q6�BU)<'#�
��p�_eRp��/dV�B��J@���U}b��U@J� �T�©oT/-��f %��o|Mo+B��U �oHi{^��dN`>�a"dM_C_��C�It$ �$n6>%�#b
�O�A�DO���q��-�~P+��=̽�.���Ʌ}Q�$敕م(4$��兝���;��.��>��H�}Q5���-�8M�Y9��M=�PU�}R&!f���	�������������� ��$�6�H�W���$CCSCH_G�RP14 2����y�&� \m.2�p)  )"��qb Fd�bN`֥���Jávh �����y�/���B����+c��?33�3�Uޢ�T�I�aD/�  C�G�P /?fff�Q>na�D ��ʹ±�W(��D©� �M�_���ɉl�~ϟπqYOφ�����F@ �����b�Dz��3����Ϡ�81�/�) �� � �$�6���Z�d�&�8� �ϴ���������� � �@����1�h�z�� ���������(�����g�@����z���R � �$�6�H�Z�`�R? Qu����� ���){M_ q��{ժ/��k/}/�/���^�� �y ��C/>�_�CR/K?" ��p&� uer2t�a 1v�`�E�i��?�` �$�!��z4�>Me&��8��$���oNL`OlH>����$lJ�/�/�/ ??(?:?_^?p?�? �?�?d_�?�?�? OO $O�_HOZO3o~O�O�O �O�O�o�O�O�o _2_ D_V_�_z_8�_�_�_ �_�_�o
oo�@o�l@i/�/-�?�Q�g�2�� ������Џ����2��/�A�S�e�w� ���������Ľ���� +tV�V�K|�������r �������y�������Ԧ*tZ��[�m�q����a>!6��}p-"�sC�>L���s��o=��y<#�
Za:rpC��������au
qb���pz�@��{�"&� ��d��oYƢ�?��b�o�{B;qc�_�����@�����.��k˰>����ʯ����X�It$� ��$�>���
z���AW���t��ߘ߼����+���:�.����F���$�=�V�(4$�b���,�;��.��>���H����5�����8M�Y���=@s������q��	�	 � ��=�(�v�h�}����������4�ڝ���  �r# �ô n�˰2��>�Pbt��y��� ��%?333��:�F�z�D/ � C'pG�P ?fff�>�G�% &^o�x���&-.� ��*)�����e�֟h�</Zz{F�@ n%z�"�{Dz�$zl/>/���m�_� �J\n ��X?��/�?�?� /Zo?"?4?F?\?j? �?ZOlO�O�?�?�?�? OO0OBO�O2_D_�O�OV\��O8/�_\/n/ �/�/�/�/�_V��_�_ go�_�_�_oo+o�o Ooao�o�o�o�o�o�o �o)�%'��/����(ȺO�s���� �]�z�H����~U� ���R��΂��
��� ��r�r�Bz��Ew��B� ���քT�ʵ���t���8Ϫ���Ș>����tȚ*�<�N�`� r�����o���̏ޏ�� ���&�8�J�\�n��� Y�������ڟ���� 2��F�X�1�|����� ���֯������0� B�(�f�x�Qߜ��� ��ߛ߭���2,�ߐ��,�=��U�2 P�y���������� ��	��"$.<�gч� �	�
���M��_ �G�)����0����K������w
c�#�>kq�-݉R8~Rӟ>L� �xϙ�.�<#�
����p�>{U��=r���#�b�f��Vw��@#Q�jr�-� ��R��J�U�&�H�B����!/B/T/ 7/x/�/=�'>{��&�/��It$ Z�/$G�>��
�/(7A��(?�/J?�/6�W +��̖5.�����5V$敕�5(4$ܾ5v?�;�;��.�5>��yH�5V5��EO8M�YE^�=�  .EV��?Oe;	\?uO `O�O�G�?�O�O�O�O�_!_�6�~3W  �pJ� '�UvUn�{QO�_�_@�_�_RB�_�^r��tpybu?333^�R_���D/  �C��G�P ?fff^>G��bu�i za��0�S_r�}��^ Xg�yb/$6WJ�2���o>����`F@� �u�a>e~�`Dz l`�t�o��Xz������ ܦo�o�o�o �o���ޏ��Zl ��l�~�������Ə�� ��ȟ� �2�D�V�h� z�����������������2��
���� � ������	�ÿ -�?�Q�c�u���Aϫ� ��O��3���)�;� ��3���I�#�5�G�Q���_�k��EW�� �����
��ڥNb� ޢ_�N*��f
&[ �����W��� ��_рEZ2��&�VG�V��Z?���$�>���V�$��ߘߪ߼��� �������(�:�L�z� ���������  ���6�H�Z�l��� H����������� <2�Vhz�� ����/�J!�S��/�/	?52t|R?d?Hv?�?�=x/�22�? �?�?�?OO/OAOSO eOwO~tu~�N�!�i j,Z�^i^iR"g�M� w/yy1_C_p_g_�V�0�W_%Y)1�W�3>���_�-�ڢk#�U>LD`+ak<�B�)<#�
��p�_�Rץ;/�V�B����e�b�2e@�3d���o�/Q b�OvZ��o���+B�e}�������`>�aWd�_xx_9�SIt$ R�-$�6>�Xb
2���AT��,���P�b��P�+����.��y����Q$敕��(4$��ҏ�;���.F�>��H�R��Q5��b�8'M�Yn��M=+`���R[!����	��џ�� ����.� �5�G�Y�k��}��o�MjΏ�  ^"���b{d&r�` �ҥ�Jס�h�����,���C�1��B���<`c��?333�U���T�I2qD/  C��G�P ?fff�Q>�a�D��޹ֱ �(��y����M�_�� �ɾ�ϒϳϦ�O �����*3�F@ `&�2����b3�DzȰ G�2�$��ϴ�E1%?9 ���&�8�J� �n�x�:�L���� ���������"�T�� $�E�|�������� ����<�����{�T������f�&�8�J� \�n�tbSe� ������ �=�as�������/��/�/�/���r�� �=y��W/> 2o�Cf/_?6��Kp: � �e�2Gt�afv�`*U *y��?�C`�$�!��@�4N�e:��8�$����obLtO�H>��� �$�J�/�/??*?<? N?'_r?�?�?�?�?x_ �?�?OO&O8Oo\O nOGo�O�O�O�O�O�o �O_�o4_F_X_j_�_ �_L�_�_�_�_�_�o o0o	�To�l}/�/A�S�e�{�2�̮���ҏ$�����2�1� C�U�g�y��������� ӟ�������?tj�j� _|�������r�������ɍ���̯ï�>t�n��o�����/���a>#!J��}A6�sW�>L�����oQ���y<#�
naNrp�W���3���*����auqv��/p��@��"":���d��omƶ�S�r�o �B Oqw�s��������0�B��k߰>3���ޯԯ���l�It$ ��$���>���
����A�k��߈��߾��+����N�.����Z��$敕j�(�4$�v�.�@�;�{�.��>��H����5����8M�Y���=������q���	�-��Q� <���|������������H�����  �r7 �״��߰F .&�3�Rdv�P
��*��, ��%?333�N�|Z���D/  C;p�G�P ?fff�>��[�%:2ro �x�:-B��>) ���/u�|�xP/nz�F@ �%0��6Dz$�$���/R/*����s� �^p���l? ��/�?�?/$/no$? 6?H?Z?p?~?�?nO�O �O�?�?�?O O2ODO�VO�OF_X_�O�Oj\� �OL/�_p/�/�/�/�/ �/�_j��_�_{o�_�_ 	oo-o?o�ocouo �o�o�o�o�o�o=�%�;�?���	8� �O�#s�����q��� `�����U���R� �₣��������� Vz�Yw��V����� h�޵�����L�x��Пܘ>���� ܚ>�P�b�t������� ��Ώ����2�ԯ:� L�^�p�����m���ʟ ��� ��$�F� �Z� l�Eϐ�����Ư��� ��� �2�D�V�<�z� ��e߰�����߯�����2,,
��.�@�Q�0�i�2d��� ������������/� 6$-.P�{ћ��	�
�� ]
�_W/�1)@����(D����@_�����ыw�7�>q�AݝR�R#ӳ>L� �#ϭ�B�O<#�
ʱ��p��R�U��Q�����7�v�z��j���@ 7Q�~r�A�	�R�@�Z�i�:�\�B�� ��5/V/h/K/�/�/Q�;>�:0�/^��It$ 
?$[�K>�
�/<7A���<?�/^??6k +�{�̪5.����5�j$敕�5(4�$��5�?�;;��=.�5>��H
Ej�5��E8M�	Y&Er�=� BEj�SOy;	p?�OtO�O�G �?�O�O�O_#_5_D[��$CCSCH_�GRP15 2����fQ?&� \Z�>]�  ғp ^3�;�U�U���Q c�_�_�_ofBo
nʆ���pvu?3�33r�Rs���D�/  C��G�P_ ?fffr>[ ��vu�i�aοD؈_1r �}��r�g�yv/Yk �^�F��os���pF@ �uqse�pDz�` ���p�z������ ��o �o�o#�GQ�� %���ʿ����ŏ׏ ���-�����U�g� y���������ӟ�ïկT�-�笸g��?� ���#�5�G�M�� ,�>���b�t������� ��v�����h�:� L�^�pϺ�h���~�X�j�|߆��K��Р� �zW0������?�8� ��b ���b_�� z&o����ʌ��� � �Ԕ�zZg���:f|��n?�;�M�Y�>�����Y����� ������'� K�]� o���Q�������� ����5�G� k�}� ������}����� 1Cqg%/�� �����	�/-�V߈�?,?>?T52@�|�?�?�?�?�=�/�22�?
OO.O@ORO dOvO�O�O�O�t�~�N �!$CiCj8,���i�i �"�����/�yf_x_�_�_�V$G0�WH_ZY(^1g�3�>��#o�-���#0e>L�y``a�*R�)<#�	
G'"p0o�R�p/�VR�����Oe�b ge@��hd�� �/����Fv��,���+B(!PeL�����	����`>�q�d�_�_n�ESItk$ ��$�6>��b	
g���ADT��a�ۏx�����P+���'��.���3��Q$�{��C�(4$�O����;��.{�>���H���Q5�=���8M�Y���M�=``���R�!П��	 ���*��c�U�j� |�������!�M��ħ  �"��b �d[r�`���J��h +�=�O�a��x�f�R����c��?33�3�U'��T3YgqD/�  C G�P /?fff�Q>�a4T ����K�(䯮�� ]�_��������π��OU���)�G*h�F@ [�g�ϵrh�Dz��|�g�Y�+���8z1Z?L9 �7�I� [�m��E�ϭ�o�� ����G���!�3�I� W��G�Y�z������� ������/�q�1����C���%ߛI� [�m�ߑߣߩCb� �T���� �<N�r��� ��/��?�ߴ/�/�/��ȧ�� �ry ֧�/J>go1S�/�?k ߲�po� �e�2|t�a �v�`_U_y/*�?2'x` /4�!֪�4AN�eo��8��$�%�L�O�H>����$�J?)?;? M?_?q?�?\_�?�?�? �?O�_O%O7OIO[O mOFo�O�O|o�O�O�O �O_�o3_E_i_{_ �_�_�_�_��_�_o o/oSoeo>��o�l@�/�/v�������2� �����*�	�B�2=�f�x��������� ҟ������)�T� tt�����|�����r �����
�¯ԯ����st��8�������d�P�q>X!��pvk�s��>Lհ��o���<#�
�a�rp��+�h�*�_���qOuSq��C�dpõ@ĴW"o� ��d���o������Br5�B�q�����/�@A�$�e�w�*{�>h����	��ߡ�It$� ��$4�>��
���A����7��߼��D�+��̃�.������C�$�=���(4$ܫ�c��u�;��.��>���H��C�5�����8M�Y��K�=@���C��q,�R�	I� b�M���q�������������}�#��   �rl 7�� ���{c[�h<ȇ����?���_���a �O%?333�K��L�����D/ � CppG�P ?fffK�>4���O% og�o�@
"o-w� K�Es)O�/#/D/7u���+/�/�z�F�@ �%�+k��DzY�$��/�/E*ց���� ܓ�� ���?�	?�?�?G/ Y/�oY?k?}?�?�?�? �?�O�O�OOO1OCO UOgOyO�O�O{_�__�O�\�_�/�_�/�/ �/�/�/�/o���_�_ �oo,o>oPoboto. �o�o<�o �o (r 5p�6?�"�4�>8�_L�Xs��2 ���ÿ������U; ���RL�;����S��� H����ɋzD��w԰�� L�2
�����4�C��G�����>���C��s������� ��͏ߏ����'�9� g�	�o���������ɟ �����ؿ#�5�G�Y� {�5Ϗ���z�ůׯ� ��)����C�U�g�y� ��qϯ������7�� @��������2a,?�Q�c�u��eߞ�2 ����������
��.� @�R�d�k$b.������ �	�
��G]KK?�T_ :Wd�f)0]Ty���Д 	��
��l�>�q�v��R8�RX��>L1xX���w�<#�
����p���U(߆����l��ů����@lQ �r�v� >�OR<��GZ���o���B��/j/�/�/ �/�/�/��p>�D�oe&?��It$ Z??$��>�E
?q7A��q??�?=?O6ޠ +����5.�����5�$敕�5(4$�E�?�;�;��.3E>��yH?E�5��OEO8M�Y[E��= wE�HшO�;	�?�O �O�O�GO_"_4_F_�X_j_��W~|W  K��p�h" p�U�U���Q��_�_@oo�B0on����pyM�u?333���R���!D/  �C��G�P ?fff�>����u�i �a�y؜_fr�}��� �g�y�/m���{������ pF@� �q�e� pDz �`4����z2��� ��o% 7��[e�'�9��� ����Ǐُ���A� ���2�i�{������� ß՟�)�ׯ�h�A����{��S���%� 7�I�[�a��@�R�� v���������п���� Ϙ�*�|�N�`�rτ� ��|��ߒ�l�~ߐߚ��_��д�*)�WD� ���S�L�#��b8  '��Зs�4$�S&� )�ʠ���0�Ԩр�Z{���o'f����?�O�a�m�>�����m��������� )�;�_�q����� e��������%�� I�[�4��������� ������!3EW �{9/����� ��/A�jߜ�.?@?R?h52�|�?�?H�?�?�=�/�22�? O0OBOTOfOxO�O�O �O�O�t�~�N1,$Wi WjL,���i�i�"���� �/�yz_�_�_�_�V+$[0�W\_nYr1gC�>�7o�-.�#��#De>L�`ta�<>R�)<#�
[;"�pDo�R ��/�VR���%!ce�b {e@ȡ|d�'�/� ���Zv��@���+B<!de`�����/���`> q�d�_x�_��YSIt$ ��-$�6>��b
{�͇AXT͏u�����P�+���;�.��y�G��Q$敕W��(4$�c��-�;���.��>��H����Q5����8'M�Y��]=t`ӕ�R�!�
�	��� >�)�w�i�~��������Ư5�M��ا  �"$��b�dor�` 3��Z ��h?�Q�c��u�����z�R��<�c�?333e;��dGY{qD/  C�( G�P ?fffa>�aHT�'�� _�(����'�/]o�� +����������Oi����=�[*|�F@ `o�{��#r|�Dz� ��{�m�?��ʎ1n?`9 �K�]�oρϓ� Y���߃�����[ �#�5�G�]�k��[� m������������� 1�C���3E����W���9߯]�o߁ߓ� �߷߽Wb��h� ��,�Pb �������*/���(?���/�/�/��Ȼ�0#�yꧠ/^> {oES�/�?�p� 0�e�2�tq�v psU syC*�?F'�`C41�@�4UN�e���8�$���9�L�O�H>��� �$�J+?=?O?a?s?�? �?p_�?�?�?�?O�_ 'O9OKO]OoO�OZo�O �O�o�O�O�O_3_�o G_Y_2}_�_�_�_�_ �_��_oo1oCo) goyoR��o�l�/�/������ą2���	��$-�>��V�2Q�z� ������ԟ���
� �#��=�h��t���� �|�����r�����֯���1��t���L���ʩ΁x�d�$q>l!��.�����>L�б���/�<#�
�a�rp���?�|�>�s���$qcugq��W�xp׵@$شk"��.��d��o������Vr'I�B �q����"�C�U�8�y���>{(�>|���'����ߵ�It$ ��$�H�>���
��)�A���)���K����X�+���̗�.������W�$敕��(�4$ܿ�w��;�{�.��>��H���W�5���8M�Y�_�=а/�W� �@�f�	]�v�a��� ������������"�1�$CCSCH�_GRP16 2����S&� \G�|/J�  � � K� ���(���o� �Pȼ���S�	��s��u �c%?333_��`������D/  C�pGÿP ?fff_�> H���c%���o1�u "�-��_�z�)c�F/ X/y/Ku3��`/�/�z�F@ �%�`��Dz�4��/�/z*�ʏ�� � ����/�?4/>?  OO|/�/�o�?�?�? �?�?�?O�O�O_BO TOfOxO�O�O�O�O_ �_�_A__�\�T_�/ ,o�/�/�/?"?4?:o ��o+o�oOoaoso�o �o�oc�o�oqU '9K]�U5��k?0E�W�i�s8�8_�� �s��g�ێ׿��,� %��Up�� b��O�L� ��g��\�ϥ���zy� �w�����g
T�Ҟ'� i�x�[��(�:�F�>���x�F��� ��̏ޏ�����8� J�\�n���>�����ȟ ڟ���׿"�4��X� j�|�����j�į֯�� ����0�^�T��x� ��������������� �l�C�u���+�A�2�,t���������2����	��-� ?�Q�c�u������$�. �����00%�|]� �t҉_oW�ߛ)Se����4��5PG	K������>�q���b�R��>�LfM����<#�
4��p��U8]߻�������� ��<���T@�QU �r /��sĄRq�3&|Z/�¤���B�=9/ �/�/�/�/�/?�˥�>�y��[?2I�t$ t?$��>�z
T?�7A1�?N?��?r?�6� +��̞E.��� E�$�敕0E(4$�x<E�?K;��.hE�>��HtE�5{���E8M�Y�E��=M�E�}ѽO�;	�?�O�O_WPOB_ W_i_{_�_�_/���~>�W  ���p ��H"�e�U���Q �o*o<oNo�BeoSn�����p��u?3�33�b� 	T!D�/  C�G�P_ ?fff�>� !�u y�a8Ϯ��_�r  ���g��/�� ��Ű�B��4�UpF@ H�Tq�e�UpDz�`i�TF��p�zg�G�9� �$ 6HZl2����\� n���4����� � 6�D�v�4�F�g����� ԟ���
��^�����v�0������� 6�H�Z�l�~�����0 u���Aϫ���Ͽ�� Ͽ�)�;���_ϱσ� �ϧϹ�߱��Ǐ������ψȔ����� _)�Wy�7�T�߁� X��bm \������i$ ��&�LL)���� e����Z��.��\f�����?/������>����Ԣ��� (�:�L�^�p�I��� ������ ��$�6� H�Z�3~���i���� ����� 2/V hz���n/�� �
/@R+?v������c?u?�?�52@�|�?�?�?OM�//B2*OSOeOwO�O�O �O�O�O�O�O�t�~^ A1a$�i�j�,ح�i�i �"�˧�/�y�_�_�_�_
f`$�0%g�_�Y(�1Qg=C�>E�lo�=c�X��#ye>L��`�a�sR9<#�	
�p"pyobU��/fLR���<%@!�e0rQ �e@���dD� \?����vتu/" /";Bq!�e����.��R�d�+p>�Uq�d o�_���SItk$ Џ$!F>��b	
���A�T���$�xΏ��1`+���p��.���|�0a$�{����(4$ܘ��P�b�;��.ĕ>���HЕ0a5�=���8M�Y�8]�=�`�0b�!�?�	 6�O�:�s�^������� ůׯ���j]���  �"Y�$r �d�rph�P�HZU�)x t�������,�����LR��N��c<�?33�38ep�9d|Y�qD/�  C] G�P /?fff8a>!q}T <�\�T��
8-���\� d]8o2�`�<����1߀$%_���rߐ*��F@ �հ��Xr��DzF��԰Ϣ�t�2�8�1�?�9 ܀ϒ� �϶��ώ����߸��� 4�FߐF�X�j�|�� ������������� 0�B�T�f�x���hz������n���� �߶���������b� ��+=Oa /��)/�/�� //_/�]?#��/?!?+����90E#�y ��/�>�ozS�/�?� (��p�90(uB�t@q �v5p�U�yx*1O{'�` x491�D�N u��!H�044�n�L�O�H>���04�J`?r?�? �?�?�?�?�_�?OO &OTO�_\OnO�O�O�O �O�o�O�O�o_"_4_ F_h_"|_�_g�_�_ �_�_oo�0oBoTo foxo^�o�o���o$|@�/-?��я���2N� ,�>�P�b�s�R���2������ӟ���	� �-�?�Q�X�O�r��� �t���|48�8�,� A'Q�S���J�A�f��t쀁���������Yq>�!ȿc�p��E�յ>L���EϢd�<#�
�a�rpտt���s�����Yq�u�q���­p�@YĠ"�� c�+t<)��4
�ϋr\~�B�q����W�x�@��m߮���s{]�>���1�\�R���It$� ,�$}�>�2�
�^�A�^���*�<捰+�����.�����匱$�=���(4$����޾�;��. �>���H,���5���<�8M�YH���=@�d���5�u���	�� �����������!�3EW��l�D.i  8�� ��U�  �]������������������ :Ø%?333������ة�D/ � C�pG�P ?fff��>}�٤�% ���of��S"�-�� ����)��Z/l/�/�u�h��t/�/�z F�@  5!t�� Dz�!4/�/�/�*���� ��� / /$/�?H/R?O&O�/ �/�o�?�?�?�?�?�? .O�O�O_VOhOzO�O �O�O�O�O_�_�_U_._�\�h_�/@o�/ ? ?$?6?H?No�-o?o �ocouo�o�o�o�ow �o�o�i;M_ q�i5��?Y�k�}��8�L_���s�{ 1���֣@�9�e� %�b����`�!Ԝ�@� �����z���w�Ԅ ��{
h��\�}��������<�N�Z�>�����Z���Ώ��� ��(��L�^�p��� ��R���ʟܟ� �� �6�H�!�l�~����� į~�د���� �2� D�r�h�&ߌ�����¿ Կ����
���.π�W� ���-�?�U�2�,����������2 ����/�A�S�e�w� �������$�.����� DD9ܐ]���ҝ_ �W�߯)gy����H��I[	_�	
����>�q$��b8b��1>Lzax��+��<#�
H�(�p1�eq����������P�	�h@�Qi�r/�� �ĘR��G&�Z-/�¸���B)�QM/�/�/�/ �/
??�˹>!���o?FIt$ Z�?$��>��
h?�7AE�?b?�?�?�6�� +���(E.����4E�$敕DE(4$�PEOK�;��.|E>��yH�E�5���EO8M�Y�E��=a �E����O�;	�?_ �O+_WdOV_k_}_�_��_�_"/���~�W  �����\" � ee 
a�,o>o@Pobo�Byogn��y��u?333��(b�4	h!D/  �C�G�P ?fff�>�5�uy qL����_�r�� �g��/��������V�*�H�ipF@� \�hq�e"ipDz �`}�hZ�,��z{�[�M� �8J\n �F����p����� H����"�4�J�X��� H�Z�{���ğ֟��� ��0�r� �2�����D��į&���J�\�n� ��������D����U� ��ѿ�������=� O���s��ϗϩϻ��� �Ņ�ۏ�������Ȩ�����s)�W�� K�h2�ߕ�l��b�  p������}$��&� ``)0���3�y0��р�Z��B��pf������?&/������>����Զ��*�<�N�`� r��]�������� ��&�8�J�\�n�G ����}��������  �4F/j|�� ���/��0 /Tf??������w?�?�?�52��?�?HOO+M
?CB2>O gOyO�O�O�O�O�O�O �O	_��*^U1u$�i �j�,��i�i�"��ߧ 	?��_�_o�_ft$�09g�_�Y�1egQC!>Yрo=w�l��#�e>L�`�a�<�R9<#�
��"�p�o,bi��/+f`R��!P%T!�eDre �e@��dX�p?� ����v쪉C"/6;B�!�e��0�B�%�f�x�++p>iq�dox
oˏ�SIt$ �-$5F>��b
ď�A�T���8���E`�+��̄�.��y���Da$敕���(4$ܬ�d�v�;���.ؕ>��H��Da5����8'M�Y �L]=�`�Db�!-�S�	J�c�N� ��r�����ǯٯ�������$CCSC�H_GRP17 �2���@��&� \�4>��79   �"m�8rt�rp���� \Z��=x����Ϳ߿@�(���`R�b��cP�?333Le��Md�Y��qD/  Cq G�P ?fffLa>5q�TPՑɉ��8 b��p�x]Log�t�P� 3�E�f�8% _��Mߧ�<�*��F@ ����M�lr��Dz{�������ߩ�g��1�?�9 ܵ�����������!� +�����i�{ߤ{�� �������������� /�A�S�e�w�������@����.��A �����������!� '�b�<N` r��P/��^/� B//&/8/J/�/B�q?`X�2?D?V?`��% n0z#�yT�
?�>�o�S ?O�]��p�n0<u 9B�tTq�vIp�U�y�* fO�'�`�4n1T�AD�Nu�VHe4H��\<'_3X>���e43Z �?�?�?�?�?�?O�_ %O7OIO[O�O+o�O�O �O�O�O�O�o_!_�o E_W_i_{_�_W�_�_ ��_�_ooKoAo� eowo�o�o�o��o�o ��Y|0?b?���.�2��a�s�������	����2������ �,�>�P�b�t����� �ާ�ҁ�t���i m�m�a�v\����@� R��v����t!����"�4�8��Γ�q>��!������z�
��>LS�:�z���<'#�
!q�p
ϩ�p�J���ݢ���q@�u�q)����pA�@� B��"�Ϙ�`tq^ � i
��r���B�*� &ߌ߭߿ߢ����ߨ{��>��fđ���H���It$ a�$��>%�g�
A��A����;��_�q�°+��=��.�������$敕�(4$��)�����;��.�U�>��Ha���5���q�8M�Y}�ɭ=:�����j�����	��������=��/DVhz����$CCSCH_G�RP18 2�����&� \��v/��  m�� �� ��5Ғ�٪�� &8J\��saݢ��� o��%?33�3ɵ"ʴ�A�D/�  C�pG�P /?fffɱ>��� �%)!%����"�- ��ɿ��)�߰/�/�/��u��P/�/$?!�c F@ V5b!���c Dz�w4b/T?&?�*8T�4�&� �2/D/ V/h/z/@O�/�?jO|O �/�/!�?
OO.ODO RO�OB_T_u_�O�O�O �O�O__*_l_o,o�_�_>l��_ ?�oD? V?h?z?�?�?�oo �oO�o�o�o�o �7I�m��� ����5��?����ӏ�8Ȣ_��sL� ���E�A������fe �Z�jb뀹Ŷ�V��� u���9�9�*��-�R� *���
��<���jӘ�����ϒ�����>���ℰ��$�6� H�Z�l�~�W�����Ɵ ؟���� �2�D�V� h�Aό���w�¯ԯ� �����.�@��d�v� ����ȿ��|����� �*��N�`�9����@��ߏq����2 < ������%��=�28�a�s��������� ������
4>$O� oԚ����]���� �_�W�9����n���3��	��_K��>S�z�pqbfb�Ӈ>L���ρ�<#�
��~�p�&ce��%Z���J�NѦ>"_о@a�R�j/ ����R�ϝ&�Z�/=��0�Bѧ�/	?*?@<??`?r?%� >c!���?�It$� �?$/�>��
�?GA�O�?2O�?��6?+���~E.�����E>$�=��E(4$ܦE^O�pK;��.�E>���H�E>5����E8M�Y�EF=@�U>��'_MK	DO ]_H_�_lW�O�_�_�_��_�_	ok�$CC�SCH_GRP1�9 2����:a&� �\.��1�  ��g�2"$�"  �eeV
�a7(�o�o�o��o:R�o�nZ�\�<�J�?333F�b�G�	�!D/  C�k�G�P ?fffF>/!�J��y�q ���\o�j�rFaw n�J?-�?�`�2���G������pF@ `Ӆ�qGuf"�pDzup ��я��a����� ܯ���� ���%����c�u��� u���������ϟ��� ѯ�)�;�M�_�q��� ����鯗���(�����;������ӏ��� 	��!Ϛ ����6� H�Z�l�~ϐ�Jߴ��� X���<�� �2�Dߎ߀<�k�R�,�>�P�Z���h�t��)Ng��� �����Wr� � h�6%3��$N!�&C � �)��`������h�Nj@;���%�fP�_�BO�|/!->��� _�-
���������� ����1�C�U���% �������������	 �?Qcu�Q/ ���/��E ;�/_q����/ ���?/S,*�\��? OO(E2}�[OmOO$�O�M�?�B2�O�O �O__&_8_J_\_n_ �_��~��^�1�$yz <c�gygy[2p�V��?���:oLoyopo�f�$�@�go.i2A�g�C�!>���o�=��t3u>LMp4qt/�R��9<#�
!�"p��b�D?�f�R���!�%�!#u�r� ;u@��<t����?Z$k��X/�c� ��"�/�;B �!$u ���������ݏ+�p>�q`t�o�o�B�cIt$ [�$��F>�ar
;���A�d��5���Y�k��`+������.������a$敕�(�4$�#�۟�;�{�.O�>��H[�޻a5��k�8M�Yw��]=4p���bd1��ʛ	��گů�� �7�)�>�P�b�t�������$CCSCH�_GRP1A 2������&� \�>|p߮9  g2 �Яr�t/��p����Z ��x �2�D�VϷ�mϔ[��R���is��?333�e��di;��D/  C� GÿP ?fff�a> �qd��� �/�8ٿ �����]�o����Ǐ�� ���߯%�_J����:]�F@ P�\����r]�Dz��q�\�N�� ���NA.O I � ,�>�P�b�t�:��ߢ� d�v�����/���� (�>�L�~�<No�� �������� $f &�~8��� �>�P�b�t��� r}�I/���� �/�/1/C/�/g/�/ �/�/�/�/?���?��0�?�?�?��Ȝ�0 �#F�˷�??N;c�? �O`��T�d�0�u�B P��qo��p3e3�$:�O '7Lp$D�1˺�D6^�ud��H�4����\�_�X>����4�ZO O0OBOTOfOxOQo�O �O�O�O _�o__,_ >_P_b_;�_�_q�_ �_�_�_o�(o:o� ^opo�o�o�o�ov��o �o $
�HZ3� ~�|�?�?k�}������2��؟�������7�22�[�m���� ����ǯٯ������ �I�i��ɔʉ���� ��؂�����ٷ�ɿ����h���-Ǚ�P����Y�E��>M1�t��k`��>�L�����{��<#�
�qx�p�� �]8���T����D� H���8�Y���@�� L2d���t�����
}�7��*�By��ŝ� �$�6��Z�l��	Ё>]�������I�t$ ��$)�>���
��
�A��
����,�����9�+��̞x�.�����8�$�敕��(4$�x��X�j�;��.���>��H��8�5{����8M�Y��@�=��8��!G�	>�WB{f���������$�CCSCH_GR�P1B 2����4&�� \(��/+�  �a0,�� ��	БyP�~1؝����4��T���V0��D5?333�@řAĄ���D/ � Ce�G�P ?fff@�>)х�D5 �)}!��V�"d=l� @�['h9D�'?9?Z?,����/A?�?��� F�@ �5�!A%`�� Dzo �4�/�?�?[:ˑ���� ܩ/�/�/ �/�/�O?O�O�O]? o?�oO�O�O�O�O�O �O�_�_�_#_5_G_Y_ k_}_�_�_�_�o�o"o�_�l�5o�?�?�? �?�?OO���o �0BTfx�D� ��R��6���,� >���6Ee�LO&�8�J�TH�ob�n���H �����ς����eQ" ���bb�0�-���H��� =а��١�Z������� b�H5�����J�Y��<�v�	��'�>���Y�'��������� џ���ο�+�=�O� }�υ�������ͯ߯ ������9�K�]�o� ��Kߥ�����ۿ��� �?�5���Y�k�}Ϗ� �χ����ϰ���M�$� V������"�2w<U��g�y�����{��2 �������� 2D Vhz�4x>����� )*�]ma)a)U�jo Pgz�|94Fsj����(,��
����>ʁ����b8�bn��>LG .!xn����<#�
���p���e>����������%�"��5%@�a6$ɂ�/�� T�ebR�6]j�/�҅���B��%?�?�?�? �?�?�?�ۆ >�!Z$��{<OIt$ ZUO$��>�["
5O�GA�O/O�OSOeF޶+����E.����U�$敕U(4$�U�O�K�;��.IU>��yHUU�5��eUO8M�YqU�=.  �U�^�_�K	�O�_ �_�_�W1_#o8oJo\o�no�o�k�$CCS�CH_GRP1C 2����a�&� �\��j���  a�ހ�"~$)2� u �e�
�a�(,>PP�RgU~��Ӏc#��?333�r�|51D/  C���G�P ?fff�>�!����q� ���o|�����w� �?����׏�ՑD���x��W�F@ J�0V��u�"W�Dz�pk��V�H��؊H�(�� �&�8�J�\�n�4� ����^�p�ڏ��� ���"�8�F�x�6�H� i�����į֯������`�� ϟ�x�2̸ �����8�J�\�n��� ����"wω�C߭Ͽ� ���������+�=��� a߳߅ߗߩ߻�ﳕ���ɟ�����ј� ������@9�g{�9�5/ ����Z��rN0^��� �%��J4�!i6� --9 ���!�F ����j�� 0�%^v�����O�/x���>����� �
��*�<�N�`�r� K����������� &8J\5/�� k/�����/" 4?Xj|��� p?���//?B/ T/-Ox/�,����eOwO�O�E2��O�O�O_]�?1R2,_U_g_ y_�_�_�_�_�_�_�_ ����nCAc4�y�z�< ڽ�y�y�2�ͷ�?��@�o�o�o�ovb4�@@'w�o�i�ASw?S�!>G�n	Me�Z��3{u>L�p�q�/ub
IO<#�
�!r2p{�rWŻ?vNb����!>5B1�u2�S0�u@ ���tF�^�	O�$��/@��ںw�12?$KBs1 �u�����0��T�f�;�>W��t�o��^�cIt$ ҟ$#VK>��r
���A�d����&�П�3p+�{��r�.���~��2q$敕��(4�$ܚ�R�d�;��=.ƥ>��Hҥ2q�5���8M�	Y�:m=�p
�2r�1�A�	8�Q�<�u�`� ������ǿٿ������$CCSCH_�GRP1D 2����.�?&� \"N��>%I  �2[� &��t�����s�Jjx� +��ϩϻ���.������Nb�P��s>�?3�33:u��;t~i��D�/  C_0G�P_ ?fff:q>#� d>��wі/HP��� ^�fm:U�b�>�!�3� T�&5o��;��:��F@ ����;�Z���Dzi��������pU��A�O�I ܣ� �������߱����� ��W�i�/i�{����� ���������/ ASew��������/��/ �����������/�r �/�/*/</N/`/r/ �/>?�/�/L?�/0?? ?&?8?�?0�_OF� O2ODON��\@h3 ��B��?�N�|cO _ �K�ˀ�\@*�'RǄ B��7��e���:T_�7 �p�D\AB�/T�^���DXSD6�p�lo!h>���SD!j�O�O �O�O�O�O�O�o_%_ 7_I_w__�_�_�_ �_�_��_o�3oEo Woio�oE��o�o���o �o�o9/�Se w����������G�OPO�����2@q�O�a�s�����u���2��ү����� ,�>�P�b�t�{�r ������ �W[�[� O�dJt�v�.�@�m�dω�߄����"�(&��Ǽ�|�>�1�������h���>L�A�(�h�򲇙<#�	
��p�ϗ��8���˲��|�����կ�Ѐ/�@|0��2 �߆�N�_L��W�������B����z��������>���T��u�6��Itk$ O�$��>�U�	
/���Aā�)���xM�_���+������.�������$�{��(4$������;��.C>���HO��5�=�_8M�Yk���=(Ї��X����	 ������+2�DVhz��$C�CSCH_GRP�1E 2�����&� �\��d?��  [��0��x�#� ��%�Ǻ���/&/@8/J/�a/O.˲��0y]ӻ5?333���"����/�D/  �C܀G�P ?fff��>�����5�) �!����v2�=㽷� �'�9��?�?�?�����>?�?O�Q0F@� DEP1�%��Q0Dz � eDP?BOO�:B�"�� � ?2?D?V? h?._�?�OX_j_�?�? ��O�O
__2_@_r_ 0oBoco�_�_�_�_�_ �_ooZo�oro,|��oO�2ODOVO hOzO�O��q�=� ��������%� 7�ɏ[���������� ���Eܟ�O�������HȐoِ�:�u� 3�/�����}�Tu�"H� Xrِ�դ�D��c�� '�'��ѯ�@��ّ����*��X&��Д���߀�����>���Д�� ��$�6�H� Z�l�Eϐ�����Ư�� ����� �2�D�V�/� z���e߰�¿Կ�� ���.��R�d�vψ� �Ϭ�j��������� ��<�N�'�r��ܛ�͟_�q�����2�<����H����+2& Oas����� ���4�>=�]�) �*}��m�)�)���o�g ���9����&\���!'����M'9��>A�h/�_rTr��u%>L� �!��<o�<#�
��l�pu/"Qu��&H����8�<�%,2M��%@�a�$@�X?��� �b�ߋ6�jq?+����Bm�%�?�?O*OONO`O�� >Q1�$�x��O�It$ �O-$>��"
�O�GA��O�O _�O�F- �+���lU.��y�xU,!$敕�U�(4$ܔUL_^[;���.�U>��H��U,!5���U8'M�Y�U4=� e,"��o;[	2_Ko6o ooZg�_�o�o�o�o�o��o{�$CCSC�H_GRP1F �2���(q�&� \����   ��U� 2�$�2� �umu Drq%8����(b(��~H�J��#8�?3334%�r5$x��1D/  CY�G�P ?fff4!>1y8�y�q���� J�X�`4/O�\�8O �-�N� ���5���<��΀F@ ��́5�T2΀Dzc��͏�����O������ ܝ�����ӏ叫�	� �կ�Q�c���c�u� ��������ﯭ���� �)�;�M�_�q�����@׿�ϗ��￩̸)� ��߯���ӟ���	� ߈"�� ߺ�$�6�H� Z�l�~�8�ߴ�F��� *���� �2�|�*�Y�`@��,�>�H��� V�b�9<w����/v �����E��0��V�$5 !�4<1�610��9�� N�� ��V�<z)��%�v>M�0_j?�<>���M� }�������������� 1Cq/y� �����/�	�/ -?Qc�??�� �?���/3/)/�? M/_/q/�/�/{?�/�/ �O�/A<�J��O�O _U2k�I_[_m__�]	oO�R2�_�_�_�_ oo&o8oJo\onou� l��n�A�4���<Q� U�U�IB^�D�nOp�( :g^�v�4	P�w�
y Q�w�Sv1>�����M����bC�u�>L;�"�b?�b�I<'#�
	1�2p��rp��2O�v�b��v1@�5�1����0)�@v� *���Տ�OH4Y�F?� Q�2y?�KB�1� �t�������˟ݟ�;z�>΁N�yo0�s�It$ I�$�V>%�O�
)�{�At{��#���G�Y��p+��=��.������q�$敕�(4$���ɯ۫;��.�=�>��HI��q5���Y�8M�Ye��m="����rRA����	��ȿ���׷%���,�>�P�b�tσ���$CCSCH_G�RP1G 2������&� \�N^�I  UB���� r��z�����j���� � �2�Dߥ�[�I��b����W���?33�3�u
Ҳt�i)�D/�  C�0G�P /?fff�q>���d ������?�H��p��� �m����鵟����5�o8���	JK�F@ >�J��тK�Dz��_�J�<����8<Q_Y ��,� >�P�b�(���Rd ����	?����, :l*<]��� ��� T//�l&,���~/,� >�P�b�t����/�k/ }/7?�/�/�/�/�/�/ �??1?�?U?�?y?�? �?�?�?���O���O�O�O��Ȋ�@�34� ��oO-^)��c~Ow_N% ��B�R"�@���R>��� ]���!u!�J�_G:� T�A�ʦT$ny�RֻX��D���zl�o�h>����D�j�O__ 0_B_T_f_?�_�_�_ �_�_��_oo,o>o Po)�to�o_��o�o�o �o��(�L^ p���d����  ����6�H�!�l���@�O�OY�k�}���2�� Ưد�����%�2 �I�[�m������ ��ǿٿ������7� W��ق�w������ƒ �����Ϸ����� �V���ׇϙɝ�G�3��>;Ab���pY"N"ߓo�>L����ߏi���<#�
��f�po��K%���B����2�6���&�G���@���:BR� ��ń�Ï���k�%����Bg��Ջ����@$��H�Z����>K�������ϭ���It$� ��$�>���
����A�����������'�+���f.����r&�$�=��(4$܎F�X;��.�>���H�&�5����8M�Y�.�=@���&�ϑ5	, E0iT�������� +�$CC�SCH_GRP1�H 2����"!&� �\��?�  ҒO@��Ԛ��� %g%>�l!�/�/�/��/"�/�.B��D@<��2E?333.Շ"�/�rɦ�D/  C�S�G�P ?fff.�>�s�2Es9k1 �� �D/�2RMZ�.�I7 VI2�O'OHO�ϵ?�/O�O���0F@ `�E�1/5N��0Dz]0 �D�?�O�OIJ������ ܗ?�?�?�?�? �_O_�_�_KO]O�� ]_o_�_�_�_�_�_�o �o�oo#o5oGoYoko }o�o�o��o�|�#�O��O�O�O�O �O_	�������� 0�B�T�f�x�2����� @�ҏ$�����,�v��$US�:_�&�8�BX�P�\���6'쟪� ��p������u?2���r P�����6���+��� �鏚H����Џ�P�6*@#������&8�G�*�d���	��>��� G��w���������ѯ 㯼���+�=�k�� s���������Ϳ��� ���'�9�K�]��9� �ϥ�~���������-� #���G�Y�k�}ߏ�u� ���ߞ���;��D�������2eLCUg$y�i��2�� ��� 2DV hoDfN������)�* ��K}O9O9C�X>wh��jI"/4/a/X/}&��� �'/)�'�p�>���/z��r�r\��%>L501\���{�<#�
���p��/�"�u,��&���p���5�2��#5@pq$4���?z�B�Sr�@�FKz�?��s��B ��5OnO�O�O�O�O�O��t0>�1H4s/i/�*_#It$ C_$��>�I2
#_uWA� $u__�_A_SV� +�����U.�����U�!$敕�U(�4$�e�_�[;�{�.7e>��HCeޣ!5��Se8M�Y_e�=0{e�"L�o�[	�_�o�o�o �go&8J\n�}{�$CCSCH�_GRP1I 2�����q&� \��|X���  O� ̐�2l4Bt0�u�u� �q�8��,�>��bU��C�����Q3��?333�%��$�#A�D/  C��GÿP ?fff�!> �1�������}�� j�ϝ��/Ƈә�O�� ��ş��2�����E�F@ 8�D����2E�DzڀY�D�6���ƚ6	 � �&�8�J�\�"����� L�^�ȟڟ�گ��� �&�4�f�$�6�Wώ� ����Ŀֿ����N� ��ߍ�f� ܸ��� x�&�8�J�\�n����� �"e�w�1�߭߿��� ���߯��+��O�� s���������0��������Ȅ��� ��.I�wi�'#?�x� qHռ�<@L���5� 8D�1WF�0%I�� �40��z�s5L�����_�?t��>�������� *<N`9/� �����/� &8J#?n�Y?� �����?/"/�? F/X/j/|/�/�/^O�/ �/�/�/?�?0?B?_ f?�<����S_e_w_�U�2��_�_�_�_m�Ob2oCoUogoyo �o�o�o�o�o�o�� ~1QQD|�|�qL��̉ ̉�B�ϻ��O癟����vPD�P��P�y�QA�-c�1>5��\��MS�H��Ci�>�L�����?cr�I<#�
�1`Bpi��E�8�O�<r���1,E 0A�� �A@��@���� 4�L��O�4�½?���e�B�?[BaA���� ����B�T�K�>E�ń����~sI�t$ ��$f>�Ƃ
���A}t򯚯����Ц!�+��̞`�.���l� �$�敕|�(4$�x��@�R�;��.���>��H�� �5{��е8M�Yܵ(}=���� ��A	�/�	&�?�*�c�Nǜ�����ϵ����������$�CCSCH_GR�P1J 2�����&�� \^��Y  �BI��� ���y�a�8zf���߀�ߩ߻������<r��>�΃,�?333�(���)�ly��D/ � CM@G�P ?fff(�>�mt,� m�e�?�H>���L�T} (�C�P�,��!�B�E��o��)����J��F�@ ����)�H���DzW��������C��Q�_�Y ܑ��� ��������E� W��?Wi{��� ����/A Sew��y/�/
/��,�/��/���� ��������?|��/�/ �??*?<?N?`?r?,O �?�?:O�?O�?OO &OpOM_4_ _2_<�/JPVC��0� �O�^��js�O�_�%9� ���"JP�b��0�Ԗ %��u���JBo�G���T JQ0�d�n����2hAT�$�^��lx>���ATzq_�_�_�_ �_�_�_�oo%o7o eo�moo�o�o�o�o ���o�o֏!3EW y3���x���� �'��۟A�S�e�w� ��o��������5�_ >_Я���
�2_�=��O�a�s���c���2 ����ҿ�����,� >�P�b�i�`��ή�Δ �����E-I�I�=�R/ 8'b�d��.�[�R�w�͔����������
��j�>�A��t��"8�"V���>L/��xV���u�<#�
��ݒp�߅��%&��ֹ���j����������@j!�B��t� <�M":���E*�m���Bޑ��h����� ~�������n�>��B��m�c�$��It$ Z=$��>�C�
oA��o�;Mޞ�+����.�������$敕�(4$����;��.1>��yH=��5��MO8M�YY��=� u��F���	�� ���/ /2/D/�V/h/w+�$CCS�CH_GRP1K 2����!�&� �\��RO��  I��@��f��n��% �%���!��??&?8?P�O?=>����@K��E?333���"��|���D/  Cʐ�G�P ?fff��>���ĩE�9�1� w��/dB�M�ͥ��7�I ���O�O�O��y�,O�Ox _��?@F@ 2U0>A�5��?@Dz�0ST�>O0__�J0��� �O O2ODOVOo zO�_FoXo�O�O���_ �_�_
o o.o`o0 Q�o�o�o�o�o�o�o�H���`�� ��Or� _2_D_V_h_ z_����_�q�+����� ��ˏݏ��%��� I���m������ퟛU�ʯ�_�������X� ~Ǡӓ(��'c�!�� ��r�k�B��26�F�Ǡ �咲2���Q����� ���	�.��ǡ�*�� �m�F6�������xǹό�>����� ��� ��$�6�H�Z� 3�~�������⿄�� ��� �2�D��h�z� S�ϰ������ϰ�
� ���@�R�d�vߤߚ� X������������*� <�`�쉯��M_q�2�L������2=O as������ �D�N .+K�v9v:k� �}�9�9����w���I@�/�/�/�/�&J�z @7{/�)�;7'��>/�V?��M�B���c5>L�0�1��]"��O<#�
z�Z�pc?�2?���66"�����&�*�5B;�5@ �q�4.�FO�����r��@yF�z_O���B[� �5O�O__�O<_N_��0>?A�4�/�/�_^x#It$ �_$K>��2
�_�WAw$��_�_o�_�V0+�{��Ze.���fe�1$敕ve(4�$܂e:oLk;��=.�e>��H�e1�5���e8M�	Y�e"-=�0�e2��)k	 o9$]Hw �o������$[