��   ?Q�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N   &S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I I9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  ��5�!IRTU�AL�/�!;LDU�IMT  ���� ���4MAX�DRI� ��5
�4.1 �%� � d%�Open han�d 1����% t?�? �"  1�3�0Close�o?�?�?	O�9�7Relax�?�?GOmO�9�6j82oOPO�OtO�3�?�O�O&_�O �6 +O__�_;_�4��FBlowi�ng�_x[  LO�W�_�_��(C�A(@%�
HG GRIP�PER�_{X
GR7EIF� HG;o��	:73�1f�_�o�_�o�[�3d%Oe�ffnen�o�k�fenf.�b\!cSchli�ess�o�jCLOSEgfmTS�AHpaЅo��o��o�l �+��O�����4� ��X�j���񏠏�ď ֏K���[���0�B��� f�۟��������G� ���}�,���P�b��� �ԯ���ίC��g� �(�b���^�ӿ���� 	ϸ�-�ܿ�(�u�$� ��H�Z���~���ߴ� ��;���_�� ߕ�D� ����zߌ���%��� ��3�m�X��@�R��� v�������3���W� ����<���`�r��� ��������Sc �8J�n��� �O��4 �Xj���/� �K/�o//0/j/�/ f/�/�/�/?�/5?�/ �/0?}?,?�?P?b?�? �?�?O�?�?CO�?gO O(O�OLO�O�O�O�O 	_�O-_�O�O;_u_`_ �_H_Z_�_~_�_�_�_ �_;o�__oo o�oDo �ohozo�o�o%�o �o[
k�@R� v���!���W� ����<���`�r��� ����̏ޏS��w� &�8�r���n�㟒��� �ȟ=����8���4� ��X�j�߯����į ֯K���o��0���T� ��ۿ�������5�� ��C�}�hϡ�P�b��� ���Ϫϼ���C���g� �(ߝ�L���p߂߼� 	��-�����c��s� ��H�Z���~����� )���&�_�� ���D� ��h�z�����%�� ��[
.@z� v���!�E� @�<�`r� ��/��S//w/ &/8/�/\/�/�/�/�/ ?�/=?�/�/K?�?p? �?X?j?�?�?O�?�? �?KO�?oOO0O�OTO �OxO�O�O_�O5_�O �Ok__{_�_P_b_�_ �_�_�_�_1o�_.ogo o(o�oLo�opo�o�o 	�o-�o�oc� 6H��~��� )��M���H���D� ��h�z����%�ԏ �[�
��.�@���d� ��럚���!�ПE��� �S���x���`�r�� �����̯�S��w� &�8���\�ѿ����̿ �ȿ=����s�"σ� ��X�j��ώ�߲����9���6�o��0�
S�end Even�ts�S�SEND�EVNT��Q�8އ� %	��Da�ta�߶�DATA������%��S�ysVar;��S�YSVw���O�%�Get�x�G�ET+���9W����Request �Menu���REQMENU?��(� ��^ߟ�Z���~�,��� ������e� 8J�n���� +�O��4� �j|��/�� #/]/H/�/0/B/�/f/ �/�/�/�/#?�/G?�/ ?}?,?�?P?b?�?�? �?O�?�?CO�?SOyO (O:O�O^O�O�O�O	_ �O_?_�O _u_$_�_ H_Z_�_�_�_o�_�_ ;o�__oo oZo�oVo �ozo�o�o%�o�o  m�@R�v ����3��W�� ���<���Ïr����� ���̏ޏ+�e�P��� 8�J���n�㟒���ޟ +�ڟO������4��� X�j���񯠯�į֯ K���[���0�B���f� ۿ��������G��� �}�,ϡ�P�bϯ��� ��߼���C���g�߀(�b߯�^��߂ߔ���$MACRO_M�AXX�������Ж�SO�PENBL ���2��ݐ���_���"�PDIM3SK�2�<�w��SU���TPDS?BEX  K��U)�2�����-�