��   P�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����PM_CFG�_T   � �$NU( HNL�  $IOD�_KEEP?ER�R_SEV?DE_V_FLG?CG	�CT
SCAN_M�ULT?CH1_wENB>CH2��SPARE1�2�3�e�   G ��i�2����  &STA�T- \ $�BD$?UPDA�TE_FW?PM�TK_DBGLV�>PMUIQEX}PE_VERS? �$CURp ��$$CLASS ? �������b��b�tION��  ��5�IRTUA�L��'/ �b� � � � //0/B/T/ f/x/ 
 ���/�/�/ �/�/�// ?2?D?V? h?z?�/�?�?�?�?�?0�?���6����:@