��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk"& 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&�B4��_sC3���r��"�A_p�d`U��@VA}DCMVROU
b��1PERIO�sF31P���2D-��32%T��1_D��2H�ĺ3��T����K�95K��K�7CL����0�ADJ����_U�drYRAUX�@�	/ 4�@C�P?a$� A�&�n@ q�UX_AXS� �JF�� 
 h�D�rӠ�C d��C�t�C�F�@�H�G�1P�FOXp4XAXI=SU� Tj��D�͡Na�E��AP@M@ �	BQ܀HR
$�IDX\PRV�QSa�G�RT�L $�F�E_Uנ���TTOOL�R�p;�A��p�y1DOf`� \��0R_PK�G�RQ BQ SNR�PBQS�P=[Q 2	hQ2�P�S�P2�Q�Q�ba	�1�ad�$VFLfw0IM�,�LT�r �:a��Tc�6Tb�����$DYG��C$d0JgGUg	�d�4�d��cMPSWP ��$ @��  �;���a   I@�`��`VERSION��h�@�5~�aIRTUAL�o��avS?�h&�  �aL|J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��a|+u|P11 29{�\�`�@�� �֓Ә��  {?�a @�`<����A�  ��� ��#����3��-�?��Q�?�g�U���� � D  Bp � =��Ϳ�?333?�a�̠�̤�@��ߥA ��/ � & G�P ?�fffˡ>�� ߥ�������0�ܙD� ��̤ˡ��k�C�Z� [��`�0�����ӿٲ��B�ђǟI�ÿ���;���F@ `K���������Dz���l�W�I��ٺ��ܑ�P`��w���ēV��'�9�K�]�o�5ߓ� ��_�q�ۿ������ �#�9�G�y�7�I�j� �߳�����������@a��!���y�3���� ϋ�9�K�]�oρϓ� ����x���D������ �����,>�b�������� ����ɤ����ȗ�Đؓ��� 2/d���L����^/\�Ϣ�]�ĐW��"�`�"��'B���������/"  $đƚ��$1>B,4_��(�����1?��?�?�8>����ā�//@/�? T/f/?O�/�/�/�/�/ �/�O??,?>?P?b? ;_�?__�?�?�?�?�? OO(O�_o^OpO�O �O�O�O�O�O�O __ $_�oH_Z_3~_�W� �fx���2������	���o2�2 -�V�h�z������� ԏ��������Dqdd �����l��ߩߩ�b�� ���o����ğ���cd�p(������qT�
@� a>Ho�
}��8[��c|�>LŠ��x�_v���<#�
�Qsbp|��X��o�C��� a?e?a��3�T`��@ �G_�
 �T���_����x�2bo%{Bta�������1� �U�g�k�`>X�ؤ�����ϑ�It$ Z��$$�>�٢
���A��߭�'������4�+���s�.����Ճa$敕��(4$ܛ�S�e��;��.��>��yH�Ճa5����O8M�Y��;�=�� �3��a�B�	9�R� =�v�a�ߡ�����������m����  �b\'����� �`k�S�K�X�,�w���@����/�����C��Qy�??333;��s�<��saD/  �C``G�P ?fff/a>$���?_	 W�_��0��_g�;� 5c?�4'e��u�j� F@� ��[�� Dz I ���w5���y ܃��� ��/���/�/7I �_I/[/m//�/�/�/ �?�?�?�/?!?3?E? W?i?{?�?kO}O�?�?�L�Oq�O��� ����O���O�O�_ 
__._@_R_d_o�_ �_,o�_o�_�_oo bo%`&/ $.(��?��>�"��o ����}��o��E+̰ �B��+��ȴC��8� ����{j4�~gĠ{t���"�������$�3t�7�q�����>���3t�cu��� �������)�W� ��_�q����������� ݏ�ȯ�%�7�I�k� %����j���ǟٟ� ��Ϳ3�E�W�i�{� a�������կ�L�o0��������2Q/�A�HS�e�v�Uώ�2�� ������������0� B�T�[Ru������ ���7M;	;	/�DO*G T�V� �M�D�i���Op�����Ѱ����A>�a��f��B�BH���>L! H�<��g�<#�
�ϲ�p��w�E�v������A��7������@\A�b�f��D ?B,��7J���_���Bб���Z{�p��N���>�4_�xU�/��It$ //-$��>�5
/a'A��a/	/�/-/?&���+����%.��y��%��$敕�%�(4$��%�/�+;���.#5>��H�/5��5��?58'M�YK5��= g5��8�x?�+	�/�?�? �?�7?�?O$O6OHO�ZO�o�GnlG  ;¸`�X�� �E�E��A��O�O�O�	_�2 _^����`<=�e?333���B������D/  C���G�P ?fff��>���e�Y�Q �iȌOVb�m����W �i�]ooo�o��k��_�wo�o�`F@ `uawU�`Dz�P $to�o�j"���� ��_�_oo'o �KoU�)��o�o� ������1�� �"�Y�k�}������� ŏ׏�ǟٟX�1����k��oC��o' 9KQ���0�B���f� x���������z���� ���l�>�P�b�t����lu�ς\�nπϊx�O�������4��� ��C�<���R(� ���c�$�C� � ��׺��ڷ  �Ę�~J@k���_V�؏��/��?�Q�]�>��� ��]���������� +��O�a�s߅߳�U� ������������9� K�$o������ ������#�5�G�u� k�)����������� ���1ǼZό�/0/B/X%2�l�/�/�/$�/�-��"2�/?  ?2?D?V?h?z?�?�? �?�d�n�>�GYGZ <���Y�Y��������ijO|O�O�O�F�K �GLO^Ib!W�#�> �'_����4U>L}PdQ�.B��<#�
K+p�4_�B�t�FB�����SU�RkU@��lT��o�δ����ζ��0o��eB ,TUPo�o�o�o�o��P>a�T�O�O�rICIt$ �$��&>��R
k�wA�HD�e���v�@+����+�.����7��A$敕G�(�4$�S���;�{�.�>��H����A5����8M�Y���==dPÅ�B�ԏ�{	�
���.� �g�Y�n����������%o�=��ȗ  B��R�T_b�P#� �J��X/�A�S�e�P�|�j�B�	��S��?333�E+��D|7IcaD/  C�G�P ?fff�A>�Q8D����O =X蟲��M�O�� �o��˿���?Y�ӿx-�Kl�F@ _�0k�ӥbl�Dz��Āk�]�/��~!^/P) �;�M�_�q���I� ����s߅���K� �%�7�M�[ߍ�K�]� ~�����������!�3�u�#�5����Sl� ��)ϟ�M�_�qσϕ� �ϭ�GR����X���� ����
�@R� v��������/�ϸ����� ��� viڗ�N.k_ =C��/o�㢄`s�� �U�"�d�Q�f�PcEci 3�/6|P3$�ښ�$ E>�Us��(��)ox�<�?�8>���� �:/-/?/Q/c/u/�/ `O�/�/�/�/?�O? )?;?M?_?q?J_�?�? �_�?�?�?O#O�_7O IO"omOO�O�O�O�O �o�O�O_!_3_oW_ i_B�_{���z���u2	�����.�F�2A�j�|� ������ď֏���� �
�-�Xqxd�����l �����b�����@Ɵ؟���!�wd�p@<������qh�T�_a>\��}z�o� s��>L٠�� o��yO<#�
�Q�bp���/�l��o.�c����_aSeWa��G�h`ǥ@ �Ȥ[s��T���_@�V�ꌿFbo9{B�a �����3�E�(�i�{�.k�>l������^��It$ ��$8�K>��
���A������;�����H�+�{�̇�.������G�$敕��(4�$ܯ�g�y�;��=.��>��H��G��5����8M�	Y�O�=���G��a0�V�	M�f�Q��u� �ߵ������� �����'��$�   �bp;������g� _�l�@���������C�(����c��e��S?333O���P����ñD/  Ct`G�P ?fffO�>8���Ss	k�_!x D�s{�O�IwS� 'H;e#��/�<�j� F@ ��/o�� Dz] �����I�q��y ܗ�����/ /�/�/K]�_]/o/ �/�/�/�/�/�?�?�? ?#?5?G?Y?k?}?�?@�?O�OO�?g|�#O ��O�����/ 	_���O�O�__0_B_ T_f_x_2o�_�_@o�_ $o�_oo,ovo$%t`:/&8B(�O Pp\cҹ6��o�~ǯ�� �o��E?��BPp?� �ܴW���L������j H��gؠ�tPq6�#������8�GtK߅���<	��>���Gt� w�������� ��+�=�k��s��� ������͏����ܯ '�9�K�]��9����� ~�ɟ۟���-�#�� G�Y�k�}���u���ů ���lD�������2eC�U�g�yߊ�	iϢ�2�������� ��� �2�D�V�h�o f���Դ������KM O	O	C�XO>Gh�j"� 4�a�X�}�ӴИ���������p�>��a��z��B�B\����>L5 \���{�<'#�
��p����p�E,ϊ�����p�@�����İ#@pA $�b�z�B�SB@� KJ���s���B� n�������t >�Hs�i�*/�It$ C/$��>%�I
#/u'A �u/�/�/A/S&��+��=��%.����%���$敕�%(4$��5�/�+;��.�75>��HC5��5���S58M�Y_5��= {5��L��?�+	�/�?�?�?�7?�O&O8OJO\OnO}K��$CCSCH_G�RP12 2�����A&� \��Xo��  O��`� lt �E�E���A� __,_>_�2U_C^�����`Q�e?33�3��R����#D/�  CаG�P /?fff��>��� �e�Y�Q�}��Ojb�m ����W�i��o�o�o����2o�o�E`F@ 8uDa�U�E`Dz�PYtDo6�j86��� �o&o 8oJo\o"��o�L�^� �o�o�����&� 4�f�$�6�W������� ď֏����N������f����x�& 8J\n�����e� w�1�������ѯ��� ���+���O���s��� �����u�Ϸ�ϣ��ϿxȄ���ٳ. ��i�'�#��x�q�H� �R<L������8� W� �����4  ����J���sLV�؂���/�t���>����Ē����� *�<�N�`�9��ߖߨ� ���ߊ�����&�8� J�#n��Y����� �����"��F�X� j�|�����^������ ���0B/f�@����S/e/w/�%2�l �/�/�/�/=�22?C?U?g?y?�?�? �?�?�?�?�d�nN1! Q|Y|Zqȝ�Y�Y� ՟����i�O�O�O�O�FP� W�O�I�!AW-3�>5�\_�pS�H��iU>L�P�Q�cB�<#�
�`pi_RE��V<B���,0�U bA�U@푡T4�Lo ��В�fȚeo��Ba�U�o�o@BT�P>Ea��T�O�O�~CIt$� �$6>��R
��wA}D������v!P+���`�.����l� Q$�=�|�(4$܈�@��R�;��.��>���H�� Q5���Ѕ8M�Y܅(M=@�P�� R�	�/�	&� ?�*�c�N����������ǟٟ�Zo Mؾ��  �I�b�T �b�PX�@�8JE�hd��v����������<B��>��S,�?333�(U`�)TlI�aD/ � CMG�P ?fff(Q>amD,� L�D�����L�TM (_"�P�,� �!���?���bπ��F�@ �Š��Hb��Dz6��Ġ���d�"ʳ!�/�) �p����� ����~�ܿ�Ϩߺ�$� 6π6�H�Z�l߂ߐ� �߀�������� � 2�D�V�h��X�j���������^����ϔ� �ϸ�������|R���� ���	-?Q u������ O��M/���/����) 5�i� ��.�_nC��/��� �`��) e�"�d0a�f %`�E�ih!?k�Ph$ )!��$z>�U��8 $�$�^o�<�?�8>��� $�:P/b/t/�/ �/�/�/�O�/�/?? D?�OL?^?p?�?�?�? _�?�?�_ OO$O6O XOolO~OWo�O�O�O �O_�O�o _2_D_V_ h_No�_�_w�_l� /����u2>���.�@�R�c�B{�2 v�����ÏՏ���� �/�A�H�?�b��q�d ةت�l$�(�(�r1� �AC����:�1�V��d�pq�ݟ��q��
��Ia>���S}��8��5sť>L���x5o��Ty<#�
�Q�bpůd���c�����Ia�e�a�|��`��@I������S d,�o۶$���{bLon{B�a��G�h�z� ]Ϟϰ�ckM�>��!��L�B��ړIt$ Z�$m�>�"�
��N�AٔN���p��,��}�+��̼�.������|�$敕��(4$��՜߮��;��.�>��yH�|�5��,�O8M�Y8儝=�� T�|�%qe��	�ߛ� �����������#��5�G���\�4Y�  (r�p�E�� M���������u�����@����x�������y*��?333����ș��D/  �C�`G�P ?fff��>m�ɔ��	 ��_Vxy�C����� ~���J\}peX���d��j� F@� ��d��� Dz � $���~���y ���� �/8B/??�� �_�/�/�/�/�/�/? �?�?OF?X?j?|?�? �?�?�?O�O�OEOO�L�XO�0_��/ /&/8/>_آ_/_�_ S_e_w_�_�_�_go�_ �_uooYo+o=oOoao �oY%�o/I[mw(�<O�p�c�k�! �~��Γ0)� Ut� R�pt�P�Č�0Ɓ� �����j}��g��t�q�k�X�֎L�m�|t��ߺ�,�>�J�>���|tJ������ ���<�N�`�r��� B�����̏ޏ���ۯ &�8��\�n������� n�ȟڟ�����"�4� b�X��|�������į ��������p�Gy��/�E�2�xߊ�H�߮߿�����2�� ����1�C�U�g�y� ��������	�4	 4
)̀M�	�	xOsG �ϟW�i��������8���9�K�O����� Q>�a��R R��!>Lj Q��<��<#�
8�p!���EaϿ����� Q��@���X@�AY�b��w� �Bu�7�Jײ����B�A=�����/��� >�}��x��_/6�It$ x/-$��>�~
X/�'A5��/R/�/v/�&���+���5.��y�$5��$敕45�(4$�@5�/
;;���.l5>��H�x5��5���58'M�Y�5��=Q �5����?�+	�/�?�? OGT?FO[OmOO�O�O��n�G  ��p��L�  U�E���A�_._@_�R_�2i_W^����`<��e?333��R���$�XD/  C��G�P ?fff��>�-��ei�Q <����O�b}����W y��o�o�o̵��Fo��o8�Y`F@ `LuXa�U Y`Dz�P mtXoJ�jk�K�=� �(o:oLo^opo 6��o�`�r��o�o8� � ��$�:�H�z�8� J�k�����Ə؏��� � �b��"���z�4������:L^p ����4y���E��� ��ӯ���	�ÿ-�?� ѿc�����������π�u���Ϸ����xȘ����c�G}�;� X&�υ�\��Rq`� �����m��� P� P ���#�i  ����J@��2�`V�����/�����>��� �Ħ���,�>�P�b� t�M��ߪ߼����ߞ� ��(�:�L�^�7�� ��m���������� $�6�Z�l�~����� ��r������  DV//z�����g/y/�/�%2�l�/�/�/$
?=�322.?W? i?{?�?�?�?�?�?�? �? t�nNE!e�Y�Z �ܝ�Y�Y��ϗ���i�O�O�O�OVd�� )W�O�I�!UWA3L>I�p_-g�\��}U>L�P�Q�wB�)<#�
�tp�}_RY��VPB��L@D�U4bU�U@��TH�`o/�䒀��fܚyo3&+B u�U�o�o 2Vh`>Ya�T_�O���CIt$ �$�%6>��R
��A��D��(���v5P+����t�.������4Q$敕��(�4$ܜ�T�f�;�{�.ȅ>��Hԅ�4Q5���8M�Y��<M=�P�4R��C�	:�S�>�w� b�������ɟ۟����noM��  �]�(b�T�b`l� T�LJY�-hx�������P0�ů��PB�R��S@�?333<Ut�=T|�I�aD/  Ca�G�P ?fff<Q>%a�D@�`�X�� (1���`�hM<_6�d� @��5�(O���xvϔ��F@ ��0���\b��DzJ��Ā����x�6��!�/�) ܄�������̿�� ��ϼ���8�JϔJ� \�n߀ߖߤ��ߔ�� �����"�4�F�X�j�|��l�~������� �r����ϨϺ����� �����R����� /ASe��- ���c��a/'�//%//�� ��= I�i#���.�_ ~C��/��,��`��=  ,e2�dDa�f9`�E�i |5?�P|$=!#�4 �>e��%84$8�rox�<�?H>���4$ Jd/v/�/�/�/�/�/ �O�/??*?X?�O`? r?�?�?�?�?�_�?�? �_O&O8OJOlO&o�O �Oko�O�O�O�O__ �o4_F_X_j_|_bo�_ �_��_(l�1/����u2R�0�B�T�f�w�V��2����ŏ ׏�����1�C�U� \�S�v��q�d���l 8�<�<�0rE�+�UW�@�!�N�E�j��d�p@���������]a>�̯g}���Is٥>L"�	�IoӒhyO<#�
�Q�bpٯ�x���w������]a�e�a�����`�@ ]�����g/d@�-o@�8�տ�b`o�{B�a ����[�|ώ�qϲ���wka�>��5�`�V��^�It$ 0�$��K>�6�
�b�A��b�
߄�.�@֑�+�{����.�����ސ�$敕��(4�$��հ���;��=.$�>��H0吡�5��@�8M�	YL嘝=	�h吢9qy��	�߯����� ����%�7�I�[�j���$CCSCH_�GRP13 2������?&� \�~E>�y  <r� ��Y��a��������� ����+��B0ʬ���>��?3�33����ܙ�D�/  C�`G�P_ ?fff��>�� ᔜ�	��_jx��W �ĝ������� ��el����j2F@ %%1���2Dz� F$1#/�p�#���y � %7I?mw/9? K?���_�/�/�/�/ ?!?S?O#ODO{?�? �?�?�?�?�?�?;O�O�OzOSO\��O�e_ /%/7/I/[/m/s_� R_d_o�_�_�_�_�_ �_�ooo�o<o�o`o ro�o�o�o�%��/~���(�qO�p�c ɠ�V��ޓe^� 5U�)�9R�p����%� ��Dƕ����j���g !��t�q�����`�9���t��οa�s��>����t��� ��)�;�M�&�q��� ����Տw�ݏ��� %�7��[�m�F����� ��ǟ韣�����3� E�W�i�����Kϱ�ï կ���߿�/��S����|�@�R�d�z�2@��߿����������2�0�B�T�f�x� ������������ �>�i	i
^̵M�	�	 ���O�G�������������=�m�n���(��.�ڱ>"qI���@R5R��V>L�� �ƿP���<#�	
m�M�pV��2U����)���ڱ��u.��@�A�!r 9�Ϭ��B��l�JR�ݿ��BN�vr���/�//A/��� >�2������/k�Itk$ �/$��>��	
�/�'Aj��/�/?x�/�& +���M5�.���Y5$�{��i5(4$�u5�-??;;��.�5>���H�55�=��58M�Y�5��=� �5���?;	 ?,OOPO;G�?{O�O �O�O�O�OG���n�G  ��6p ��� EU-U%�2Q Q_c_u_�_	B�_�^)���+p�u?33�3MRY��D/�  C:�G�P /?fff>�Z� u9i1aq���
_�b9} A�g=y/�o�o����{o�oOmʎ`F@ �u�a�U5�`Dz#`�t�oQz8�р�r� �]ooo �o�o�ok��o����� #m�#�5�G�Y�o� }���m����׏��� ��1�C�U���E�W�֟��i���K��o �����ϯi�� ��z������,�>� ��b�t�Ϙ�꿼�ο ��<��u:� ���������͟�"Ø �G��pލW��Ϻߑ� b�����Ң ����U��XǞ  U���J��g���V�؂�?K������>������=�O�a� s߅ߗߩ߂������� �1���9�K�]�o�� ��l��������� #�E��Y�k�D���� ���������1 CU;y�d/�@��
ߜ/�/�/�%2+| 	??-???P=//h22c?�?�?�?�?�?�? �?
OO.O5t,~ONz! ��Y�Z��ii	" ��./0y�O�O'__CV�� ^W�O�I�!�Wv3��>~��_@-p����"#�U>L�P��Q"�BA)<#�
��p�_QR���PV�B����uy�Uib��U@6��T}o @/��f��oh9[+B��U�o4U@gJ��P:`>�a�d9_/_��CIt$� 	�$Z6>�b
�;�A�D;��]����jP+��̩�.������iQ$�=�Ņ(4$�х��ޛ�;��.��>���H	�iQ5����8M�Y%�qM=@�PA�iR!R�x�	o� ��s������ן�����"�4��oIM!�F�  "��]b2d �b:`�����J��bh�����ѯ�e���讅B���cu�?333�qU��rT�I�aD/ � C�G�P ?fffqQ>Za�Du� �����C(f�0͝M q_k���u7�I�j�]�EO׿Qϫ���F�@ ���Q��b�Dz�����ϭ�k��!�/�) ܹ�˿ݿ ����%�/����m� ��ߑߣߵ����� �������3�E�W�i� {���������2�����E������� ����%�+�R
 �@Rdv��T ��b�F*< N�FՖ/\�6/H/Z/d��)�r ~�iX� /�.�_�C/?��a� p��r ae=2�dyav n`�E�i�j?��P�$ r!X�E4�>9e�Z8i$�m��oL+O7H>���i$7J�/�/�/�/ �/�/?�O)?;?M?_? �?/_�?�?�?�?�?�? �_O%O�_IO[OmOO �O[o�O�O�o�O�O_ !_O_E_i_{_�_�_ �_�o�_�_�o]l4/ f/�
��2�2��e��w��������Ă2 �������0�B�T� f�x����ĈΫ��q�d !�!�|m�q�q�erz� `����D�V���z����d%���&�8�<��
҃��>���}��8��~s�>LW�>�x~o��y<#�
%arp�����N��������e�a-�Ų�`E�@��F��� ddu�bo$�m�
��b�o�{Bq.�*ϐϱ��� �����Ϭk��>�j�𕯋�L�#�It$ Ze�$��>�k�
E���A"���?߹�c�u��Ơ+����.�����š$敕!�(4$�-������;��.Y�>��yHe�š5��u�O8M�Y��͝=>� ��Ţnq����	���� �����A�3�H�Z�l��~�������}��  qr�����9� ������ݚ��	@-?��VD���ys��?333ͥ�Τ�E�D/  �C�`G�P ?fff͡>�����	 �)o�x������ͯ ���ϓ���e���3�/%zFF@� 9%E��FDz � Z$E7/	/�X�8�*� �'9K ]#?��/M?_?�� %o�/�/�/?'?5?g? %O7OXO�?�?�?�?�? �?�?OOO�O_�OgO!\��O/y_'/9/K/ ]/o/�/�_!�f_x_2o �_�_�_�_�_�_�oo ,o�oPo�oto�o�o�o �o�%��/����(ȅO�p�cPɴ�j (�E��yr�IU�^� MR�p����Z�ձy�ʰ =�=�zƏwV���q��������M���t����u�����>����t�����+�=� O�a�:���������� �����'�9�K�$� o���Z�����ɟ۟�� ���#���G�Y�k�}� ����_�ůׯ���� �1�C��g�����T�f�xߎ�2�����H������� �2� D�V�h�z������ �������2�R�}	 }
r��M�	�	���O�G �������������Q���������B.�9�>6q]��TRIR��j>L� �ڿ<d���<#�
��apj	FU��=���9�-�1��!B��@�A�5rM���� �B����Jf ���Bb����///C/U/�� >F���x���/�It$ �/-$�>��
�/�'A~��/�/?�/�&" �+���a5.��y�m5!$敕}5�(4$܉5A?S;;���.�5>��H��5!5���58'M�Y�5)�=� �5!��
O0;	'?@O+O dOOG�?�O�O�O�O�O��O[��n�G  ��Jp���  YUAU9�FQe_w_�_��_B�_�^=��?p<�-u?333)aR�*m��D/  C�N�G�P ?fff)>n�-uMiEa ����_�bM}U�)#g Qy-/�o"���o�	c�ʢ`F@ `�u�a	eI�`Dz7` �t�o�e#z�є߆� �qo�o�o�o�o ��o�����%7�� 7�I�[�m�����Ï�� ��������!�3�E� W�i���Y�k��ß}����_կ���� ���}¯ԯ���� 
��.�@�R��v��� Ϭ���п����Pπ�uN���� �����*�6ìW�τ� �k����ߥ�b��� *��Ҷ1�&�� �i�"�lǲ i�*�Z@��{���V�!�%?�_������>��� !���Q�c�u߇ߙ߫� �ߖ�������E��� M�_�q������ ����%�7�Y� m��X�������� ���!3EWiO ��x/���߰/�/�/�%2?|?/?A?$S?d=C/|22w?�? �?�?�?�?�?OO0O BOIt@~cN�!��Y�Z �%�)i)i"2��B/�Dy�O_;_2_WV��� rW�O�I�!�W�3J>���_T-����6#�U>L`�Q6�B�U)<#�
��p��_eR��/dV�B��J���U}b��U@J��T�©oT/-���f%��o|Mo+B ��U�oHi{^��dN`>�a"dM_C_���CIt$ �$�n6>�#b
�O�A��DO��q��-�~P+���̽�.����Ʌ}Q$敕م(�4$�兝���;�{�.�>��H��}Q5��-�8M�Y9��M=�PU�}R&!f���	�������� ����� ��$�6�H��W��$CCSCH�_GRP14 2����y�&� \m.|2�p)  )" ��qbFd�bN`֥���J ávh�����y�/����B���+c��?333�Uޢ�T�I�a�D/  C�GÿP ?fff�Q> na�D��ʹ±�W(�� D©ͱM�_���ɉl� ~ϟ�qYOφ�����F@ �����b�Dz��3�����Ϡ�1�/�) � � ��$�6���Z�d� &�8�ϴ�������� �� ��@����1�h� z����������(� ����g�@����z��� R ��$�6�H�Z�` �R?Qu��� �����){ M_q��{ժ/��0k/}/�/���^��  �y��C/>�_�CR/ K?"��p&� uer2 t�a1v�`�E�i��? �`�$�!��z4�>Me&��8�$���oNL`OlH>����$lJ�/ �/�/??(?:?_^? p?�?�?�?d_�?�?�?  OO$O�_HOZO3o~O �O�O�O�O�o�O�O�o  _2_D_V_�_z_8�_ �_�_�_�_�o
oo� @o�li/�/-�?�Q�g��2�̚�����Џ����2��/�A�S� e�w����������Ľ� ���+tV�V�K|���� ���r�������y�������Ԧ*tZ��[�Pm�q����a>!�6��}-"�sC�>�L��s��o=��y<#�
Za:rpC��8������au 
qb���pz�@��{� "&���d��oYƢ�?��b�o�{B;qc�_� ���������.��k˰�>���ʯ����X�I�t$ ��$�>���
z���AW���t���ߘߪ���+��̞:�.���F���$�敕V�(4$�xb��,�;��.���>��H����5{����8M�Y���=s������q��	�	 ���=�(�v�h� }���������4�ڝ�>��  �r#  �ôn�˰2� �>Pbt��y��� ��%?3�33�:�F�z�D�/  C'pG�P_ ?fff�>� G�%&^o�x��� &-.���*)��� ��e֟h�</Zz{F@ n%z�"�{Dz�$zl/>/p���m�_� �J \n��X?��/�? �?�/Zo?"?4?F? \?j?�?ZOlO�O�?�? �?�?OO0OBO�O2_D_�O�OV\��O8/�_ \/n/�/�/�/�/�_V� �_�_go�_�_�_oo +o�oOoao�o�o�o�o �o�o�o)�%'��/����(ȺO�s �����]�z�H���� ~U����R��΂�� 
�����r�r�Bz��Ew ��B����քT�ʵ���t��8Ϫ���Ș>����tȚ*�<� N�`�r�����o���̏ ޏ�����&�8�J�\� n���Y�������ڟ� ���2��F�X�1�|� �������֯����� �0�B�(�f�x�Qߜ������ߛ߭���2@,����,�=��U�2P�y������ ������	��"$.<� gчĲ	�
���M ��_�G�)����0����K����(��wc�#�>kq��-݉R~Rӟ>L�� �ϙ�.�<#�	
����p�>{U��=r���#�b�f��Vw��@#Q�jr �-���R��J�U�&�H�B����!/�B/T/7/x/�/=�'>�{�&�/��Itk$ �/$G�>��	
�/(7A��(?�/J?x�/6W +��̖5�.����5V$�{���5(4$ܾ5�v?�;;��.�5>���H�5V5�=�E8M�YE^��=� .EV��?Oe;	 \?uO`O�O�G�?�O�O �O�O_!_�6�~3W  �pJ �'�UvUn�{QO �_�_�_�_RB�_�^r���tpbu?33�3^�R_���D/�  C��G�P /?fff^>G�� bu�iza��0�S_r�} ��^Xg�yb/$6W�J�2��o>����`F@ �u�a>e~�`Dzl`�t�o��Xz8���߻� ܦo�o �o�o�o���ޏ�� Zl��l�~������� Ə����ȟ� �2�D� V�h�z�����������������2��
�� ��� ������ 	�ÿ-�?�Q�c�u��� Aϫ���O��3��� )�;υ�3���I�#�5�G�Q���_�k�� EW�Ϲ����
��ڥ Nb�ޢ_�N*��f 
&[�����W���  ��_�EZ2��&�VG�V�Z?���$�>���V�$��ߘߪ� �����������(�:� L�z�������� �� ���6�H�Z� l���H��������� ��<2�Vhz ������/�J@!�S��/�/	?52t| R?d?v?�?�=x/�22�?�?�?�?OO/O AOSOeOwO~tu~�N�! �ij,Z�^i^iR" g�M�w/yy1_C_p_g_�V�0�W_%Y)1�W�3>���_�-p�ڢk#�U>LD`�+ak�B�)<#�
�p�_�Rץ;/�V�B����e�b�2e@�3d���o �/Qb�OvZ��o���+B�e}�@������`>�a�Wd�_x_9�SIt$� R�$�6>�Xb
2���AT��,���P��b��P+����.�������Q$�=��(4$��ҏ��;��.F�>���HR��Q5���b�8M�Yn��M=@+`���R[!����	�� џ������.� �5�G��Y�k�}��o�MjΏ�  ^"���b{d &r�`�ҥ�Jס�h�����,���C�1��B����`c��?333�U�T�I2qD/ � C�G�P ?fff�Q>�a�D�� ޹ֱ�(��y����M �_���ɾ�ϒϳϦ��O Ϛ���*3�F�@ &�2����b3�DzȰG�2�$��ϴ�E1%?9 ���&� 8�J��n�x�:�L�� �����������"� T��$�E�|���� ��������<�����{�T������f�&� 8�J�\�n�tbSe ������� �=�as� �����/��/�/�/���r�� �=y�� W/>2o�Cf/_?6�� Kp:� �e�2Gt�afv �`*U*y��?�C`�$ �!���4N�e:��8�$����obLtO�H>����$�J�/�/?? *?<?N?'_r?�?�?�? �?x_�?�?OO&O8O o\OnOGo�O�O�O�O �O�o�O_�o4_F_X_ j_�_�_L�_�_�_�_ �_�oo0o	�To�l}/ �/A�S�e�{�2�̮����ҏ�����2 �1�C�U�g�y����� ����ӟ�������?t j�j�_|�������r�� ����ɍ���̯ï�>tn��o�����/�
��a>#!J��}A86�sW�>L����x�oQ��y<#�
naNrpW���3���*����auqv��/p��@��"":�� �d��omƶ�S�r�o �BOqw�s������ ��0�B��k߰>3����ޯԯ��l�It$ Z��$��>���
����Ak��߈��߾���+���N�.����Z��$敕j�(4$�v�.�@��;��.��>��yH���5����O8M�Y���=�� ����q���	�-� �Q�<���|������������H�����  �r7 �״�� ߰F.&�3�Rd@v�
��*��, y��%?333��N�Z���D/  �C;pG�P ?fff�>��[�%: 2ro�x�:-B�� >)���/u��|�P/nz�F@� �%��6Dz $�$��/R/*����s� �^p�� �l?��/�?�?/$/ no$?6?H?Z?p?~?�? nO�O�O�?�?�?O O 2ODOVO�OF_X_�O�Oj\��OL/�_p/�/�/ �/�/�/�_j��_�_{o �_�_	oo-o?o�oco uo�o�o�o�o�o�o =�%;�?���	8��O�#s����� q���`�����U�� �R��₣����� ����Vz�Yw��V������h�޵������LϾ�Пܘ>����ܚ>�P�b�t��� ������Ώ����2� ԯ:�L�^�p�����m� ��ʟ��� ��$�F�  �Z�l�Eϐ�����Ư ��ꯨ�� �2�D�V� <�z���e߰�����߯�����2,,
��H.�@�Q�0�i�2d� ������������� �/�6$-.P�{ћ��	 �
��]
�_W /�1)����(D����_�����ыw�7�>q�AݝR�R#ӳ>L� �#�<��B�<#�
ʱ�p�R�U��Q����7�v�z��j���@7Q�~r�A�	� R��Z�i�:�\�B����5/V/h/K/�/�/Q�;>�:x0�/��It$ 
?-$[�>�
�/<7A��<?�/^??6k �+��̪5.��y��5j$敕�5�(4$��5�?�;;���.�5>��H�
Ej5��E8'M�Y&Er�=� BEj�SOy;	p?�OtO �O�G�?�O�O�O_#_�5_D[�$CCSC�H_GRP15 �2���fQ�&� \�Z�]�   ғp^3�;�U�U ���Qc�_�_�_ofB(o
n����pvu?333r�Rs����D/  C��G�P ?fffr>[��vu�i�aοD� �_1r�}��r�g�yv/ Yk�^�F��os�<��pF@ �uqse�pDz�` �����z������ ��o�o�o#�G Q��%���ʿ���� ŏ׏���-����� U�g�y���������ӟ@�ïկT�-�笸g� �?����#�5�G� M��,�>���b�t��� ������v����� h�:�L�^�pϺ�h���`~�X�j�|߆��K� �Р��zW0������ ?�8���b ���b _��z&o����� ����� �Ԕ�zZg���:f|��n?�;�<M�Y�>�����Y� ����������'�  K�]�o���Q���� ��������5�G�  k�}�������}���� �1Cqg%/ �������	 �/-V߈�?,?>?T52�|�?�?�?�?�=	�/�22�?
OO.O @OROdOvO�O�O�O�t �~�N�!$CiCj8,�� �i�i�"�����/�yf_ x_�_�_�V$G0�W�H_ZY^1g�3�>���#o�-���#0e�>Ly``a�*R�)<'#�
G'"p0o�Rp�p/�VR���@��Oe�b ge@�� hd���/����Fv ��,���+B(!Pe L����	����`>q�d�_�_n�ES�It$ ��$�6>%��b
g���ADT���a�ۏ�����P+��=�'�.���3��Q�$敕C�(4$��O���;��.�{�>��H���Q5�����8M�Y���M=``���R�!П��	���*��c� U�j�|�������!�M|��ħ  �" ��b�d[r�`���J ��h+�=�O�a��x��f�R���c��?333�U'��T3Ygq�D/  C GÿP ?fff�Q> �a4T����K�(� ���]�_����� ������OU���)�G*h�F@ [�g�ϵrh�Dz��|�g�Y��+���z1Z?L9 � 7�I�[�m��E�ϭ� o������G���!� 3�I�W��G�Y�z��� ����������/�q� 1����C���%� �I�[�m�ߑߣߩ Cb��T���� �<N�r� ����/��?��0�/�/�/��ȧ��  �ry֧�/J>go1S�/ �?k߲�po� �e�2 |t�a�v�`_U_y/*�? 2'x`/4�!֪�4AN�eo��8�$�%�L�O�H>����$�J? )?;?M?_?q?�?\_�? �?�?�?O�_O%O7O IO[OmOFo�O�O|o�O �O�O�O_�o3_E_ i_{_�_�_�_�_��_ �_oo/oSoeo>� �o�l�/�/v��������2������*�	�B�2=�f�x����� ����ҟ������ )�T�tt�����|��� ��r�����
�¯ԯ����st��8���P����d�P�q>X!���vk�s��>�Lհ���o���<#�
�a�rp��+�h8�*�_���qOu Sq��C�dpõ@Ĵ W"o���d���o������Br5�B�q���� �/�A�$�e�w�*{��>h���	��ߡ�I�t$ ��$4�>��
���A�����7�����D�+��̞��.�����C�$�敕��(4$�x��c�u�;��.���>��H��C�5{����8M�Y��K�=���C��q,�R�	I�b�M���q���� ��������}�#��>   �rl  7�ķ��{c[�h <ȇ���?����_��a �O%?3�33K��L�����D�/  CppG�P_ ?fffK�>4� ��O%og�o�@
" o-w�K�Es)O�/#/ D/7u��+/�/�z�F@ �%�+k��DzY�$��/�/pE*ց���� ܓ �����?�	?�? �?G/Y/�oY?k?}?�? �?�?�?�O�O�OOO 1OCOUOgOyO�O�O{_�__�O�\�_�/�_ �/�/�/�/�/�/o�� �_�_�oo,o>oPobo to.�o�o<�o �o (r 5p�6?�"�4�>8�_L�Xs ��2���ÿ����� �U;���RL�;���� S���H����ɋzD��w ԰��L�2
�����4�C�G�����>���C��s��� ������͏ߏ���� '�9�g�	�o������� ��ɟ�����ؿ#�5� G�Y�{�5Ϗ���z�ů ׯ���)����C�U� g�y���qϯ�����忀7��@��������2@a,?�Q�c�u��e���2����������
� �.�@�R�d�k$b.�� �����	�
��G]KK ?�T_:Wd�f)0]Ty���Д 	(����l�>�q��v��R�RX��>L�1X���w�<#�	
����p���U(������l��ů����@lQ �r �v�>�OR<��GZ���oϑ�B��/j/��/�/�/�/�/��p>��Doe&?��Itk$ ??$��>�E	
?q7A��q??�?x=?O6� +����5�.����5�$�{���5(4$�E��?�;;��.3E>���H?E�5�=�OE8M�Y[E���=wE�HшO�;	 �?�O�O�O�GO_"_ 4_F_X_j_��W~|W  K��p� h"p�U�U���Q� �_�_oo�B0on�����pM�u?33�3��R���!D/�  C��G�P /?fff�>��� �u�i�a�y؜_fr�} ����g�y�/m����{����� pF@ �q�e� pDz�`4����z82��� ��o %7��[e�'�9� ������Ǐُ�� �A����2�i�{��� ����ß՟�)�ׯ�h�A����{��S�� �%�7�I�[�a��@� R��v���������п ����Ϙ�*�|�N�`� rτ���|��ߒ�l�~��ߚ��_��д�*) �WD����S�L�#� �b8 '��Зs�4$� S&�)�ʠ���0 �ԨюZ{���o'f�肟��?�O�a�m�>�����m������� ��)�;�_�q�� ����e�������� %��I�[�4����� ����������!3 EW�{9/��� ����/A�@jߜ�.?@?R?h52�| �?�?�?�?�=�/�22�?O0OBOTOfOxO �O�O�O�O�t�~�N1 ,$WiWjL,���i�i�" �����/�yz_�_�_�_�V+$[0�W\_nYr1gC�>�7o�-p.�#��#De>L�`�ta�>R�)<#�
[;"pDo�R ��/�VR���%!ce�b {e@ȡ|d�' �/����Zv��@���+B<!de`��@���/���`> q�d�_�_��YSIt$� ��$�6>��b
{�͇AXT͏u������P+���;�.����G��Q$�=�W�(4$�c���-�;��.��>���H���Q5�����8M�Y��]=@t`ӕ�R�!�
�	� ��>�)�w�i�~��������Ư5�M��ا  �"$��b�d or�`3��Z ��h?��Q�c�u�����z�R����c�?333�e;�dGY{qD/ � C( G�P ?fffa>�aHT� '��_�(����'�/] o��+�����������Oi���=�[*|�F�@ o�{��#r|�Dz���{�m�?��ʎ1n?`9 �K�]�o� �ϓ�Y���߃���� �[�#�5�G�]�k� ��[�m����������� ��1�C���3E����W���9߯]�o� �ߓߥ߷߽Wb�� h���,� Pb������ �*/��(?���/�/�/��Ȼ�0#�y� �/^>{oES�/�?� �p�0�e�2�tq�v  psUsyC*�?F'�`C4 1��4UN�e���8�$���9�L�O�H>����$�J+?=?O?a? s?�?�?p_�?�?�?�? O�_'O9OKO]OoO�O Zo�O�O�o�O�O�O_ 3_�oG_Y_2}_�_�_ �_�_�_��_oo1o Co)goyoR��o�l�/ �/������ą2����	��-�>��V�2 Q�z�������ԟ� ��
��#��=�h��t �����|�����r ����֯���1��t��L���ʩ΁x�
d�$q>l!��.��8���>L�бx��/�<#�
�a�rp��?�|�>�s���$qcugq��W�xp׵@$شk"��.� �d�o������Vr'I�B�q����"�C�U� 8�yߋ�>{(�>|����'���ߵ�It$ Z��$H�>���
��)�A��)���K�����X�+��̗�.������W�$敕��(4$ܿ�w���;��.��>��yH��W�5���O8M�Y�_�=а /�W� �@�f�	]�v� a����������������"1�$CCS�CH_GRP16 2���S�&� �\G�/J�  �� K� ���(�� �o��Pȼ���PS�	�s��u �c%?333_��`�|����D/  C�p�G�P ?fff_�>H���c%���o 1�u"�-��_�z�) c�F/X/y/Ku3��`/x�/�z�F@ �%0�`��Dz�4���/�/z*�ʏ�� �����/�? 4/>? OO|/�/�o�? �?�?�?�?�?O�O�O _BOTOfOxO�O�O�O��O_�_�_A__�\� T_�/,o�/�/�/?"? 4?:o��o+o�oOoao so�o�o�oc�o�oq U'9K]�U5���k?E�W�i�s8� 8_���s��g�ێ׿ ��,�%��Up�� b�� O�L���g��\�ϥ�� �zy��w�����g
T� Ҟ'� i�x�[��x(�:�F�>���x� F�����̏ޏ���� �8�J�\�n���>��� ��ȟڟ���׿"�4� �X�j�|�����j�į ֯������0�^�T� �x������������ �����l�C�u���+�A�2�,t����������2����	� �-�?�Q�c�u����� �$�.�����00%� |]��t҉_oW�ߛ)@Se����4�@�5G	K������>�q��b�R��>LfM����O<#�
4��p��U]߻�����������<���T@ �QU�r /��sĄRq�@3&|Z/�¤���B� =9/�/�/�/�/�/?�˥>�y��[?^2It$ t?$��K>�z
T?�7A1��?N?�?r?�6� +�{��E.��� E��$敕0E(4�$�<E�?K;��=.hE>��HtE��5���E8M�	Y�E��=M�E�}��O�;	�?�O�O_W POB_W_i_{_�_�_/����~�W   ���p��H"�e�U ���Q�o*o<oNo�B(eoSn����p��u?333�b� 	�T!D/  C�G�P ?fff�>�!�u y�a8Ϯ� �_�r ���g��/ ����Ű�B��<4�UpF@ H�Tq�e�UpDz�`i�T�F���zg�G�9� �$6HZl2�� ��\�n���4���� � �6�D�v�4�F�g� ����ԟ���
��@^�����v�0���� ���6�H�Z�l�~��� ��0u���Aϫ���Ͽ ��Ͽ�)�;���_� �σϕϧϹ�߱��`Ǐ�߳���ψȔ� ����_)�Wy�7�T �߁�X��bm \���� ��i$��&�LL)� ���e����Z��.��\f�����?/��<����>����Ԣ� ��(�:�L�^�p�I �������� �� $�6�H�Z�3~���i ��������� 2 /Vhz���n/ ���
/@R +?v�����c?u?�?�52�|�?�?�?OM	�//B2*OSOeOwO �O�O�O�O�O�O�O�t �~^A1a$�i�j�,ح �i�i�"�˧�/�y�_ �_�_�_
f`$�0%g��_�Y�1Qg=C�>�E�lo=c�X��#ye�>L�`�a�sR9<'#�
�p"pyobpU��/fLR���@<%@!�e0rQ �e@�� �dD�\?����v تu/" /";Bq!�e ���.��R�d�+p>Uq�d o�_���S�It$ Џ$!F>%��b
���A�T�એ$�Ώ��1`+��=�p�.���|�0a�$敕��(4$�ܘ�P�b�;��.�ĕ>��HЕ0a5�����8M�Y�8]=�`�0b�!�?�	6�O�:�s�^��� ����ůׯ���j]|���  �" Y�$r�d�rph�P�HZ U�)xt�������,������LR�N��c<�?3338ep�9d|Y�q�D/  C] GÿP ?fff8a> !q}T<�\�T��
8-� ��\�d]8o2�`�<��� �1�$%_���rߐ*��F@ �հ��Xr��DzF��԰Ϣ��t�2��1�?�9 � �ϒϤ϶��ώ����� ����4�FߐF�X�j� |������������ ��0�B�T�f�x��� hz������n� ��ߤ߶�������� �b���+= Oa/��)/�/ ��//_/�]?#�0�/?!?+����90 E#�y��/�>�ozS�/ �?�(��p�90(uB �t@q�v5p�U�yx*1O {'�`x491�D�N u��!H044�n�L�O�H>���04�J`? r?�?�?�?�?�?�_�? OO&OTO�_\OnO�O �O�O�O�o�O�O�o_ "_4_F_h_"|_�_g �_�_�_�_oo�0o BoTofoxo^�o�o�� �o$|�/-?��я����2N�,�>�P�b�s�R���2������ӟ� ��	��-�?�Q�X�O� r����t���|48� 8�,�A'Q�S���J�A�f��t쀁��P�������Yq>�!�ȿc���E�յ>�L��EϢd�<#�
�a�rpտt��8�s�����Yq�u �q���­p�@Y� �"��c�+t<)��4
�ϋr\~�B�q���� W�xߊ�m߮���s{]��>��1�\�R���I�t$ ,�$}�>�2�
�^�A�^�����*�<捰+��̞��.����匱$�敕��(4$�x����;��. ��>��H,���5{��<�8M�YH���=�d���5�u���	������������ !3EW��l�D.>i  8��  ��U� �]������ �������ʨ��� :Ø%?3�33�����ة�D�/  C�pG�P_ ?fff��>}� ٤�%���of��S" �-������)��Z/l/ �/�uh��t/�/�z F@  5!t�� Dz�!4/�/�/p�*���� �� � //$/�?H/R?O &O�/�/�o�?�?�?�? �?�?.O�O�O_VOhO zO�O�O�O�O�O_�_�_U_._�\�h_�/@o �/ ??$?6?H?No� -o?o�ocouo�o�o�o �ow�o�o�i; M_q�i5��?Y�k�}��8�L_���s �{1���֣@�9� e�%�b����`�!� ��@֑����z���w �Ԅ��{
h��\�}�������<�N�Z�>�����Z���Ώ �����(��L�^� p�����R���ʟܟ�  ���6�H�!�l�~� ����į~�د����  �2�D�r�h�&ߌ��� ��¿Կ����
���.π��W����-�?�U�2@�,�����������2����/�A�S� e�w��������$�.�� ���DD9ܐ]�� �ҝ_�W�߯)gy����H��I[	(_�	����>�q$��bb��1>L�za��+��<#�	
H�(�p1�eq����������P�	�h@�Qi�r /�߇ĘR��G&�Z-/�¸���B)�QM/�/��/�/�/
??�˹>�!���o?FItk$ �?$��>��	
h?�7AE�?b?�?x�?�6� +���(E�.���4E�$�{��DE(4$�PE�OK;��.|E>���H�E�5�=��E8M�Y�E���=a�E����O�;	 �?_�O+_WdOV_k_ }_�_�_�_"/���~�W  ���� �\"� ee 
a� ,o>oPobo�Byogn�����u?33�3�(b�4	h!D/�  C�G�P /?fff�>�5 �uyqL����_�r� ��g��/��������V�*�H�ipF@ \�hq�e"ipDz�`}�hZ�,��z8{�[�M� �8J \n�F����p��� ��H����"�4�J� X���H�Z�{���ğ֟ �����0�r� �2�����D��į&���J� \�n���������D�� ��UϿ�ѿ����� ��=�O���s��ϗϩ� �����Ņ�ۏ�������Ȩ�����s) �W��K�h2�ߕ�l� �b� p������}$� �&�``)0���3�y 0����Z��B��pf�����?&/������>����Զ��*�<� N�`�r��]����� �����&�8�J�\� n�G����}������ �� �4F/j| �����/�� 0/Tf??��@����w?�?�?�52� �?�?OO+M
?CB2>OgOyO�O�O�O�O �O�O�O	_��*^U1 u$�i�j�,��i�i�" ��ߧ	?��_�_o�_ft$�09g�_�Y�1egQC!>Yрo=pw�l��#�e>L�`�a��R9<#�
��"p�o,bi��/+f`R��!P%T!�eDre �e@��dX�p ?�����v쪉C"/6;B�!�e��0�@B�%�f�x�++p>iq��do
oˏ�SIt$� �$5F>��b
ď�A�T���8�⏼�E`+��̄�.������Da$�=���(4$ܬ�d��v�;��.ؕ>���H�Da5�����8M�Y �L]=@�`�Db�!-�S�	J� c�N���r�����ǯٯ�������$CC�SCH_GRP1�7 2����@�&� �\4>��79  �"m�8rt�rp ����\Z��=x����Ϳ�߿@����`R�b�<�cP�?333Le���Md�Y�qD/  C�q G�P ?fffLa>5q�TPՑɉ� �8b��p�x]Log� t�P�3�E�f�8% _���Mߧߤ*��F@ `����M�lr��Dz{� �����ߩ�g��1�?�9 ܵ��������� ��!�+�����i�{ߤ {����������� ����/�A�S�e�w��� ��������.��A���������� �!�'�b�< N`r��P/�� ^/�B//&/8/J/�/�B�q?X�2?D?V?`��%n0z#�yT�
?�> �o�S?O�]��p� n0<u9B�tTq�vIp�U �y�*fO�'�`�4n1T�@AD�Nu�VHe4H���\'_3X>��� e43Z�?�?�?�?�?�? O�_%O7OIO[O�O+o �O�O�O�O�O�O�o_ !_�oE_W_i_{_�_W �_�_��_�_ooKo Ao�eowo�o�o�o� �o�o��Y|0?b?���.�2��a�s���$��������2��� ����,�>�P�b�t� ���Ԅާ�ҁ�t�� �im�m�a�v\�����@�R��v����t�!���"�4�8��Γ�q>�!������z�
�>LS�:�z����<#�
!q�p�
ϩ��J���ݢ���q�u�q)����pA�@�B��"�Ϙ�`tq�^ �i
��r���B �*�&ߌ߭߿ߢ����ߨ{��>��fđ����H��It$ a�$���>�g�
A��A����;��_�q�°+�����.�������$敕�(�4$�)�����;�{�.U�>��Ha����5��q�8M�Y}�ɭ=:�����j�����	������ ��=�/DVhz����$CCSCH�_GRP18 2�����&� \��|v/��  m� � ��5Ғ�٪ ��&8J\��s�aݢ�� o��%?333ɵ"ʴ�A��D/  C�pGÿP ?fffɱ> ����%)!%��� �"�-��ɿ��)�߰/ �/�/�u��P/�/$?!�c F@ V5b!���c Dz�w4b/T?�&?�*T�4�&� � 2/D/V/h/z/@O�/�? jO|O�/�/!�?
OO .ODORO�OB_T_u_�O �O�O�O�O__*_l_ o,o�_�_>l��_ ? �oD?V?h?z?�?�?�o o�oO�o�o�o�o �7I�m� ������5��?0����ӏ�8Ȣ_� �sL����E�A���� ��fe�Z�jb뀹Ŷ� V���u���9�9�*�� -�R�*���
��<���jӘ����ϒ�����>���ℰ�� $�6�H�Z�l�~�W��� ��Ɵ؟���� �2� D�V�h�Aό���w�¯ ԯ������.�@�� d�v�����ȿ��|�� ����*��N�`�9� ���̭�ߏq����2 <������%��=�28�a�s����� ����������
4> $O�oԚ����]� ����_�W�9����n���3�P�	��_K��>S��z�qbfb�Ӈ>�L���ρ�<#�
��~�p�&ce8��%Z���J� NѦ>"_о@a� R�j/����R�ϝ&�Z�/=��0�Bѧ�/ 	?*?<??`?r?%� �>c!��?�I�t$ �?$/�>��
�?GA�O�?�2O�?�6?+��̞~E.����E>$�敕�E(4$�x�E^OpK;��.�E�>��H�E>5{���E8M�Y�EF=�U>��'_MK	DO]_H_�_lW�O�_��_�_�_�_	ok�$�CCSCH_GR�P19 2����:a&�� \.��1�  ��g�2"$ �" �eeV
�a7(�o��o�o�o:R�o�nZ��\��J�?333�F�bG�	�!D/ � Ck�G�P ?fffF>/!�J� �y�q���\o�j�r Fawn�J?-�?�`�2���G������pF�@ Ӆ�qGuf"�pDzup��я��a������ ܯ�� �����%����c� u���u���������ϟ ���ѯ�)�;�M�_� q�������鯗���(�����;������ӏ ���	��!Ϛ �� ��6�H�Z�l�~ϐ�J� ����X���<�� �2� Dߎ�<�k�R�,�>�P�Z���h�t��)Ng �������Wr � �h�6%3��$N!�& C ��)��`������ h�Nj;���%�fP�_��BO|/!->���_�-
������ ��������1�C�U� ��%������������ �	�?Qcu �Q/���/�� E;�/_q�� ��/���?/S,*� \��? OO(E2}�[O�mOO�O�M�?�B2 �O�O�O__&_8_J_ \_n_�_��~��^�1�$ yz<c�gygy[2p� V��?��:oLoyopo�f�$@�go.i2A�g
�C�!>���o�=�8�t3u>LMp4qxt/�R�9<#�
!�"p�b�D?�f�R���!�%�!#u�r� ;u@��<t����? Z$k�X/�c� ��"�/�;B�!$u ������� ��ݏ+�p>�q`t��o�oB�cIt$ Z[�$�F>�ar
;���Ad��5���Y�k�޼`+�����.������a$敕�(4$�#�۟��;��.O�>��yH[��a5��k�O8M�Yw��]=4p ���bd1��ʛ	��گ ů���7�)�>�P�b��t������$CCS�CH_GRP1A 2������&� �\�>p߮9  g2�Яr�t/��p� ���Z��x �2�D�V�P��m�[��R���is��?333�e��d|i;�D/  C� �G�P ?fff�a>�qd��� �/ �8ٿ�����]�o���� Ǐ�߼��߯%�_J���x�:]�F@ P�0\����r]�Dz��q�\�N� ���NA.O I �,�>�P�b�t�:� �ߢ�d�v�����/�� ��(�>�L�~�<N o���������� �$f&�~8� ��>�P�b�t�� ��r}�I/�� ���/�/1/C/�/ g/�/�/�/�/�/?����?��?�?�?��� ��0�#F�˷�??N; c�?�O`��T�d�0 �u�BP��qo��p3e3� $:�O'7Lp$D�1˺�D 6^�ud��H�4���x�\�_�X>����4 �ZOO0OBOTOfOxO Qo�O�O�O�O _�o_ _,_>_P_b_;�_�_ q�_�_�_�_o�(o :o�^opo�o�o�o�o v��o�o $
�H Z3�~�|�?�?k�}�����2��؟�������7�22�[�m� �������ǯٯ��� ����I�i��ɔʉ� �����؂������@��ɿ����h���@-Ǚ�����Y�E��>M1t��k`��>L�����{��O<#�
�qx�p��� �]���T�����D�H���8�Y���@ ��L2d���t��@���
}�7��*�By� �ŝ��$�6��Z�l��	�>]��������^��It$ ��$)�K>���
��
�A���
���,�����9�+�{��x�.������8�$敕��(4�$ܠ�X�j�;��=.��>��H��8��5����8M�	Y��@�=��8��!G�	>�WB{f ���������$CCSCH_�GRP1B 2����4?&� \(��/>+�  �a0 ,�Ԭ�	БyP�~ 1؝���4���T��V0��D5?3�33@řAĄ���D�/  Ce�G�P_ ?fff@�>)� ��D5�)}!��V�" d=l�@�['h9D�'?9? Z?,���/A?�?��� F@ �5�!A%`�� Dzo �4�/�?�?p[:ˑ���� ܩ/ �/�/�/�/�O?O�O �O]?o?�oO�O�O�O �O�O�O�_�_�_#_5_ G_Y_k_}_�_�_�_�o�o"o�_�l�5o�? �?�?�?�?OO�� �o�0BTfx �D���R��6�� �,�>���6Ee�LO&�8�J�TH�ob�n� ��H�����ς��� �eQ"���bb�0�-��� H���=а��١�Z��� ����b�H5�����J�Y�<�v�	��'�>���Y�'����� ����џ���ο�+� =�O�}�υ������� ͯ߯������9�K� ]�o���Kߥ�����ۿ ����?�5���Y�k� }Ϗϡχ����ϰ��πM�$�V������"�2@w<U�g�y�����{���2��������  2DVhz�4x>� ����)*�]ma)a) U�joPgz�|94Fsj����((,������>ʁ�����b�bn��>L�G .!n����<#�	
���p���e>�����������%�"��5%@�a6$ɂ �/��T�ebR�6]j�/�҅ߧ�B��%?�?��?�?�?�?�?�ۆ >��!Z$�{<OItk$ UO$��>�["	
5O�GA�O/O�OxSOeF�+����E�.���U�$�{��U(4$�U��O�K;��.IU>���HUU�5�=�eU8M�YqU��=. �U�^�_�K	 �O�_�_�_�W1_#o8o�Jo\ono�o�k�$C�CSCH_GRP�1C 2�����a&� �\��j���  a�ހ�"~$)2 � u�e�
�a�(,@>P�RgU~��Ӏyc#��?333��r�51D/  �C��G�P ?fff�>�!��� �qߏ��o|���� �w��?����׏�Ց�D�����W�F@� J�V��u�"W�Dz �pk�V�H��؊H�(�� �&�8�J�\� n�4�����^�p�ڏ� �����"�8�F�x� 6�H�i�����į֯� ����`�� ϟ�x�2̸�����8�J�\� n�������"wω�C� �Ͽ����������+� =���a߳߅ߗߩ߻� ﳕ��ɟ�����јȖ�����@9�g{� 9�5/����Z��rN0 ^���%��J4�!i6�  --9���!�F ����j��0�%^v�����O�/���>�����
��*�<�N� `�r�K���������� �&8J\5/ ��k/���� �/"4?Xj|� ��p?���// ?B/T/-Ox/�,����eOwO�O�E2��O�OH�O_]�?1R2,_ U_g_y_�_�_�_�_�_ �_�_����nCAc4�y �z�<ڽ�y�y�2�ͷ �?���o�o�o�ovb4�@'w�o�i�ASw?S�!>G�n	Me�Z��3{u>L�p�q�/<ub
I<#�
�!r2�p{rWŻ?vNb���!>5B1�u2�S0�u@���tF�^�	O�$ ��/��ںw�12?$KBs1�u�����0��T�f�;�>W��tx�o���cIt$ ҟ-$#V>��r
���A�d���&�П�3p�+���r�.��y�~�2q$敕���(4$ܚ�R�d�;���.ƥ>��H�ҥ2q5���8'M�Y�:m=�p
�2r�1�A�	8�Q�<� u�`�������ǿٿ������$CCSC�H_GRP1D �2���.��&� \�"N��%I   �2[�&��t�����s� Jjx�+��ϩϻ���.�(����Nb�P��s>�?333:u��;t~i���D/  C_0G�P ?fff:q>#�d>��wі/H P���^�fm:U�b�>� !�3�T�&5o��;��<�:��F@ ����;�Z���Dzi���������U��A�O�I ܣߵ������߱�� �����W�i�/i�{� ������������� /ASew��@������/ ��/����������� /�r�/�/*/</N/ `/r/�/>?�/�/L?�/ 0???&?8?�?0�_O`F� O2ODON�� \@h3��B��?�N�|c O _�K�ˀ�\@*� 'RǄB��7��e���: T_�7�p�D\AB�/T�^���DXSD6�p�l<o!h>���SD!j �O�O�O�O�O�O�O�o _%_7_I_w__�_ �_�_�_�_��_o� 3oEoWoio�oE��o�o ���o�o�o9/� Sew������ ���G�OPO�����2q�O�a�s�����	u���2��ү��� ��,�>�P�b�t�{� r������ �W [�[�O�dJt�v�.� @�m�dω�߄��Ǡ�"�&��Ǽ�|�>��1�φ���h����>LA�(�h�򲇙<'#�
��p�ϗ�p�8���˲��|�@����կ�Ѐ/�@| 0��2�߆�N�_L�� W�߮����B��� �z���������>��T��u�6�ïIt$ O�$��>%�U�
/���Aā��)���M�_���+��=���.��������$敕(4$������;��.�C>��HO��5���_8M�Yk��=(Ї��X����	������+�2DVhz���$CCSCH_G�RP1E 2�����&� \��d?��  [��0�� x�#��%�Ǻ��� /&/8/J/�a/O.˲���0]ӻ5?33�3��"����/�D/�  C܀G�P /?fff��>���� �5�)�!����v2�= 㽷��'�9��?�?�?�����>?�?O�Q0F@ DEP1�%��Q0Dz� eDP?BOO�:8B�"�� � ?2? D?V?h?._�?�OX_j_ �?�?��O�O
__2_ @_r_0oBoco�_�_�_ �_�_�_ooZo�oro,|��oO�2O DOVOhOzO�O��q �=������� ��%�7�ɏ[������ �������Eܟ�O�������HȐoِ�:� �u�3�/�����}�Tu �"H�Xrِ�դ�D�� c��'�'��ѯ�@� �ّ���*��X&���Д���߀�����>���Д�� ��$� 6�H�Z�l�Eϐ����� Ư������� �2�D� V�/�z���e߰�¿Կ �����.��R�d� vψ϶Ϭ�j������� ����<�N�'�r���@��͟_�q�����2�< ��������+2&Oas��� �����4�>=� ]�)�*}��m�)�)�� �o�g���9����&\���!'����M'9��>A�h/�p_rTr��u%>L� �!��o�<#�
��l�pu/"Qu��&H����8�<�%,2M�%@�a�$@�X? ����b�ߋ6�jq?+����Bm�%�?�?O@*OONO`O�� >Q1��$���O�It$� �O$>��"
�O�GA��O�O _�O��F- +���lU.����xU,!$�=��U(4$ܔUL_�^[;��.�U>���H�U,!5����U8M�Y�U4=@� e,"��o;[	2_ Ko6oooZg�_�o�o�o��o�o�o{�$CC�SCH_GRP1�F 2����(q&� �\���  ��U� 2�$�2�  �umuDrq%8�����(b��~H�J�<�#8�?3334%�r�5$x�1D/  C�Y�G�P ?fff4!>1y8�y�q� ���J�X�`4/O� \�8O�-�N� ����5�����΀F@ `��́5�T2΀Dzc� �͏����O������ ܝ�����ӏ� ��	��կ�Q�c��� c�u���������ﯭ� ����)�;�M�_�q� ����׿�ϗ��￩��)ϋ�߯���ӟ� ��	�߈"�� ߺ�$� 6�H�Z�l�~�8�ߴ� F���*���� �2�|�*�Y�@��,�>�H���V�b�9<w��� �/v�����E��0�� V�$5!�4<1�610� �9��N�� ��V�<z@)��%�v>M�0_�j?�>��� M�}����������� ���1Cq/ y������/� 	�/-?Qc�?? ���?���/3/ )/�?M/_/q/�/�/{? �/�/�O�/A<�J��O�O _U2k�I_[_m_$_�]oO�R2�_�_ �_�_oo&o8oJo\o nou�l��n�A�4�� �<Q�U�U�IB^�D�nO�p�(:g^�v�4�	P�w
y Q�w�Sv1>����M����bC�u>L;�"�b?�b��I<#�
	1�2p���r��2O�v�b��v1�5�1����0)�@v�*���Տ�OH4YF?�Q�2y?�KB �1��t�������˟ݟ�;z�>΁N�yo�0�sIt$ I�$��V>�O�
)�{�A�t{�#���G�Y��p+�����.�������q$敕�(�4$��ɯ۫;�{�.=�>��HI�ީq5��Y�8M�Ye��m="����rRA����	��ȿ��� ׷%��,�>�P�b�t�����$CCSCH�_GRP1G 2������&� \�N|^�I  UB ����r��z�����j ����� �2�Dߥ�[ߔI��b���W���?333�u
Ҳt�i)��D/  C�0GÿP ?fff�q> ���d������?�H�� p����m����鵟�� ����5�o8���	JK�F@ >�J��тK�Dz��_�J�<�����<Q_Y � �,�>�P�b�(��� Rd����	?���� ,:l*<]� ����� T //�l&,��� ~/,�>�P�b�t����/ �k/}/7?�/�/�/�/ �/�/�??1?�?U?�? y?�?�?�?�?���O��0�O�O�O��Ȋ�@ �34���oO-^)��c~O w_N%��B�R"�@���R >���]���!u!�J�_ G:�T�A�ʦT$ny�RֻX�D���zl�o�h>����D�j�O __0_B_T_f_?�_ �_�_�_�_��_oo ,o>oPo)�to�o_��o �o�o�o��(� L^p���d�� �� ����6�H�!� l����O�OY�k�}����2��Ưد�����%�2 �I�[�m�� ������ǿٿ����� �7�W��ق�w���� ��ƒ�����Ϸ����� �V���ׇ�P�ɝ�G�3��>;A�b���Y"N"ߓo�>�L�П�ߏi���<#�
��f�po��K%8���B����2� 6���&�G���@��� :BR���ń�Ï���k�%����Bg��Ջ� ���$��H�Z���Ё>K������ϭ���I�t$ ��$�>���
����A�����������'�+��̞f.���r&�$�敕�(4$�x�FX;��.��>��H�&�5{���8M�Y�.�=���&�ϑ5	,E0iT�������� +�$�CCSCH_GR�P1H 2����"!&�� \��?�  ҒO@��� ����%g%>�l!�/��/�/�/"�/�.B���D@��2E?333�.Շ"/�rɦ�D/ � CS�G�P ?fff.�>�s�2E s9k1�� �D/�2RMZ� .�I7VI2�O'OHO��ϵ?/O�O���0F�@ �E�1/5N��0Dz]0�D�?�O�OIJ������ ܗ?�?�? �?�?�_O_�_�_KO ]O��]_o_�_�_�_�_ �_�o�o�oo#o5oGo Yoko}o�o�o��o�|�#�O��O�O �O�O�O_	����� ���0�B�T�f�x�2� ����@�ҏ$����� ,�v�$US�:_�&�8�BX�P�\���6' 쟪���p������u?2 ���rP�����6��� +��Ş鏚H����Џ� P�6*#������&8�G��*d���	��>���G��w������� ��ѯ㯼���+�=� k��s���������Ϳ ������'�9�K�]� �9�ϥ�~������� ��-�#���G�Y�k�}� ��u���ߞ���;�� D�������2eLC�Ugy�i��2 ����� 2 DVhoDfN����� �)�*��K}O9O9C�X >wh�jI"/4/a/X/}&�� �'/)�'
�p�>���/z��r8�r\��%>L501x\��{�<#�
���p�/�"�u,��&���p���5�2��#5@pq$4���?z� B�Sr@�FKz�?��s���B��5OnO�O�O �O�O�O��t0>�1H4�s/i/*_#It$ ZC_$�>�I2
#_uWA $u__�_A_SVޤ +����U.�����U�!$敕�U(4$�e�_�[�;��.7e>��yHCe�!5��SeO8M�Y_e�=0 {e�"L�o�[	�_�o �o�o�go&8J�\n}{�$CCS�CH_GRP1I 2����q�&� �\��X���  O�̐�2l4Bt0�u �u��q�8��,�>�P�bU�C�����Q3��?333�%��$|�#AD/  C���G�P ?fff�!>�1������� }��j�ϝ��/Ƈә �O����ş��2���x��E�F@ 8�0D����2E�DzڀY��D�6��ƚ6	 ��&�8�J�\�"� ����L�^�ȟڟ�گ ����&�4�f�$�6� Wώ�����Ŀֿ�����N���ߍ�f� ܸ ���x�&�8�J�\�n� �����"e�w�1�߭� �������߯��+�� O��s������������������� ������.I�wi�'#? �x�qHռ�<@L��� �5�8D�1WF�0%I ���40��z� s5L�����_�?xt��>����� ���*<N` 9/������/� &8J#?n� Y?������?/ "/�?F/X/j/|/�/�/ ^O�/�/�/�/?�?0? B?_f?�<����S_e_w_�U2��_�_�_�_m�Ob2oCoUo goyo�o�o�o�o�o�o ��~1QQD|�|�qL ��̉̉�B�ϻ��O�@�����vPD�P@���y�QA�-c�1>5�\��MS�H��Ci�>L�����?cr�IO<#�
�1`Bpi���EթO�<r����1,E0A�� �A@��@ ����4�L��O�4�½?@���e�B�?[BaA ��������B�T�K�>E�ń����^~sIt$ ��$fK>�Ƃ
���A}t�򯚯���Ц!�+�{��`�.���l�� �$敕|�(4�$܈�@�R�;��=.��>��H�� ��5��е8M�	Yܵ(}=���� ��A	�/�	&�?�*�c�N� ���ϣϵ�����������$CCSCH_�GRP1J 2�����?&� \^��>Y  �BI� �鄔��y�a�8zf� ��ߗߩ߻�������<r�>�΃,�?3�33(���)�ly��D�/  CM@G�P_ ?fff(�>� mt,�m�e�?�H>��� L�T}(�C�P�,��!� B�E�o��)����J��F@ ����)�H���DzW��������pC��Q�_�Y ܑ� ���������� �E�W��?Wi{� ������ /ASew��y/�/
/��,�/��/ ������������?|� �/�/�??*?<?N?`? r?,O�?�?:O�?O�? OO&OpOM_4_ _2_<�/JPVC ��0��O�^��js�O�_ �%9⹐�"JP�b�� 0�Ԗ%��u���JBo�G ���TJQ0�d�n����2hAT$�^��lx>���ATzq_�_ �_�_�_�_�_�oo %o7oeo�moo�o�o �o�o���o�o֏!3 EWy3���x�� ���'��۟A�S� e�w���o�������㏀5�_>_Я���
�2@_�=�O�a�s���c���2����ҿ���� �,�>�P�b�i�`��� ��Δ�����E-I�I� =�R/8'b�d��.�[�R�w�͔�������(��ת�j�>�A���t��"�"V���>L�/��V���u�<#�	
��ݒp�߅��%&��ֹ���j������⾐�@j!�B ��t�<�M":���E*����m���Bޑ��h������~�������n�>���B�m�c�$��Itk$ =$��>�C�	
oA��o�x;M��+�����.������$�{���(4$����;��.1>���H=��5�=�M8M�YY�́=�u��F���	 �����/ /�2/D/V/h/w+�$C�CSCH_GRP�1K 2�����!&� �\��RO��  I��@��f�� n��%�%���!��??@&?8?�O?=>����@yK�E?333����"�����D/  �CʐG�P ?fff��>���ĩE�9 �1�w��/dB�M�ͥ� �7�I���O�O�O��y��,O�O _��?@F@� 2U>A�5��?@Dz �0ST>O0__�J0��� �O O2ODO VOozO�_FoXo�O�O ���_�_�_
o o.o`o 0Q�o�o�o�o�o �o�oH���`����Or� _2_D_ V_h_z_����_�q�+� ������ˏݏ�� %���I���m������ ퟛUʯ�_�������X�~Ǡӓ(��'c� !����r�k�B��26� F�Ǡ�咲2���Q��� �����	�.��ǡ��*���m�F6�������ǹό�>�������� ��$�6� H�Z�3�~�������� ������ �2�D�� h�z�S�ϰ������� ��
����@�R�d�v� �ߚ�X���������� ��*�<�`�쉯��M_q�2�L��H����2 =Oas���� ���D�N .+K�v9 v:k��}�9�9����w ���I�/�/�/�/�&J�z 7{/�)�;7'��>/�V?��M�B���c5>L�0�1��<]"��<#�
z�Z�pc?2?���66"����&�*�5B;��5@�q�4.�FO���� �r��yF�z_O���B[�5O�O__�O<_N_��0>?A�4�/x�/�_x#It$ �_-$>��2
�_�WAw$�_�_o�_�V0�+���Ze.��y�fe1$敕ve�(4$܂e:oLk;���.�e>��H��e15���e8'M�Y�e"-=�0�e2��)k	 o9$ ]Hw�o����� �$[