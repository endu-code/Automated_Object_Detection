��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk" 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&�B4��_sC3���rs�"�A_p�d`U��@VA}DCMVROU
b��1PERIO�sF31P���2D-��32%T��1_D��2H�ĺ3��T����K�95K��K�7CL����0�ADJ����_Uzdr���AUX�@��	 4�@C�P?a$� A�&�n@� qUX_AXS��XP  LD�� ?
 h�D�r Ӡ�Cd��C�t�C�F�@��H�G1P�FOYq3XA�XISU� T@j��D͡�q�E��AP@M@ 	BQ܀HR�
$IDX\PRV�QS�a�GRT�L w$F�E_Uנz���TTOOL�R��p;�Aѡp�y1DO�f` \��0R_gPKG�RQ BQO NR�PBQ5S�P[Q H��Rf�P2�S�P2�Q��Qba	�1�ad�$VF�Lw0IM�,�LT �r�:a��Tc�6Tb��>��$DYG��C)$d0JgGUg	�d�4�d�cMPSWP  ��$ @��  �����a�@&�@ �&�`VERSIO�N�h  ��5�aIRTU�AL�o�avS?��h&�   �aL|J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T��f�x��a+u|P11 ;29{\�@p��� ֓Ә���  ?�a �@�@����A�  �����#����3��-�?�Q�?�g�U�����  D  �Bp  =���~��?333?�a��̠�̤@��ߥA /  & GÿP ?fffˡ>��ߥ������� 0�ܙD���̤ˡ�� k�C�Z�[��`�0������ӿٲ��B�ђ�ǟI�ÿ��;���F@ K���������Dz��l�W�I��ٺD��ܑ�P`��w���ēV��'�9�K�]� o�5ߓ���_�q�ۿ� �������#�9�G�y� 7�I�j�߳������� ����a��!���y�3����ϋ�9�K�]� oρϓϙ���x���D �����������, >�b������� ����ɤ����ȗ�Đؓ ���2/d���L����^/\�Ϣ�]�ĐW�(�"�@�"��'B����������/"   $đƚ�$1>B,4_��(����1?��?�?�8>����ā�/ /@/�?T/f/?O�/�/ �/�/�/�/�O??,? >?P?b?;_�?__�?�? �?�?�?OO(O�_o ^OpO�O�O�O�O�O�O �O __$_�oH_Z_3 ~_�W��fx��Ł2�����	���o2�2-�V�h�z��� ����ԏ������� �Dqdd�����l��ߩ ߩ�b�����o����ğ���cd�p(���P���qT�@� a>H�o�
}��[��c|�>�LŠ���_v���<#�
�Qsbp|��X�8�o�C��� a?e ?a��3�T`��@ � G_�
�T���_����x�2bo%{Bta���� ���1��U�g�k�`�>X�ؤ����ϑ�I�t$ ��$$�>�٢
���A��߭��'�����4�+��̞s�.���Ճa$�敕��(4$�x��S�e�;��.���>��H�Ճa5{����8M�Y��;�=���3��a�B�	9�R�=�v�a�ߡ� ����������m���>�  �b\ '������`k�S�K�X� ,�w�������/������C��Q�??3�33;�s�<��saD�/  C``G�P_ ?fff/a>$� ��?_	W�_��0�� _g�;�5c?� 4'e��u�j� F@ ��[�� DzI ���wp5���y ܃ �����/���/ �/7I�_I/[/m// �/�/�/�?�?�?�/? !?3?E?W?i?{?�?kO}O�?�?�L�Oq�O �������O�� �O�O�_
__._@_R_ d_o�_�_,o�_o�_ �_oobo%`&/ $.(��?��>� ��"��o����}��o� �E+̰�B��+��ȴ C��8�����{j4�~g Ġ{t��"�������$�3t7�q�����>���3t�cu ��������� �)�W���_�q����� ������ݏ�ȯ�%� 7�I�k�%����j��� ǟٟ���Ϳ3�E� W�i�{�a�������կ��L�o0��������2@Q/�A�S�e�v�U���2�߲��������� ��0�B�T�[Ru� ���������7M;	;	 /�DO*GT�V� �M�D�i���Op�����(Ѱ����A>�a���f��B�BH���>L�! H���g�<#�	
�ϲp��w�E�v������A��7������@\A�b �f��D?B,��7J���_���Bб���Z�{�p��N���>��4_�U�/��Itk$ //$��>�5	
/a'A��a/	/�/x-/?&��+����%�.����%��$�{���%(4$��%��/�+;��.#5>���H/5��5�=�?58M�YK5��= g5��8�x?�+	 �/�?�?�?�7?�?O $O6OHOZO�o�GnlG  ;¸`� X���E�E��A� �O�O�O	_�2 _^�����`=�e?33�3���B�����D/�  C��G�P /?fff��>��� �e�Y�Q�iȌOVb�m ����W�i�]ooo�o���k��_wo�o�`F@ uawU�`Dz�P$to�o�j8"���� ��_�_ oo'o�KoU�)� �o�oﯥ���� �1���"�Y�k�}� ������ŏ׏�ǟٟX�1��̸k��oC��o '9KQ���0� B���f�x��������� z�������l�>�P� b�t���lu�ς\�n��ϊx�O����� ��4�����C�<�� �R(����c�$� C� ���׺��ڷ   �Ę�~Jk���_V�؂���/�?�Q�]�>�����]������ ����+��O�a�s� �߳�U���������� ���9�K�$o��� ����������#� 5�G�u�k�)������ ��������1Ǽ@Zό�/0/B/X%2�l �/�/�/�/�-��"2�/? ?2?D?V?h? z?�?�?�?�d�n�>� GYGZ<���Y�Y� ������ijO|O�O�O�FK �GLO^Ib!W�#�> �'_�p���4U>L}P�dQ�.B�<#�
K+p4_�B�t�FB�����SU�RkU@��lT��o �δ���ζ��0o��eB,TUPo�o�o@�o�o��P>a��T�O�OrICIt$� �$�&>��R
k�wAHD�e����v�@+���+�.����7��A$�=�G�(4$�S����;��.�>���H���A5�����8M�Y���==@dPÅ�B�ԏ�{	� 
���.��g�Y�n����������%o�=��ȗ  B��R�T _b�P#��J��X/��A�S�e��|�j�B��	��S��?333��E+��D7IcaD/ � CG�P ?fff�A>�Q8D�� ��O=X蟲��M �O���o��˿����?Y�ӿ-�Kl�F�@ _�k�ӥbl�Dz���k�]�/��~!^/P) �;�M�_� q���Iߧ���s߅�� �K��%�7�M�[� ��K�]�~�������� ���!�3�u�#�5�����Sl���)ϟ�M�_� qσϕϧϭ�GR���� X��������
� @R�v���� ���/�ϸ����ȫ�� viڗ �N.k_=C��/o�� �`s���U�"�d�Q�f �PcEci3�/6|P3$ �ښ�$E>�Us��(���)o�<�?�8>�����:/-/?/Q/ c/u/�/`O�/�/�/�/ ?�O?)?;?M?_?q? J_�?�?�_�?�?�?O #O�_7OIO"omOO�O �O�O�O�o�O�O_!_ 3_oW_i_B�_{�� �z���u2	������.�F�2 A�j�|�������ď֏ �����
�-�Xqxd �����l�����b�� ���Ɵ؟���!�wd�p<������qh�
T�_a>\��}z�8o� s��>L٠��x o��y<#�
�Q�bp��/�l��o.�c���_aSeWa��G�h`ǥ@�Ȥ[s� �T���_�V�ꌿFbo9{B�a�����3�E� (�i�{�.k�>l������ϥ�It$ Z��$8�>��
���A�����;������H�+��̇�.������G�$敕��(4$ܯ�g�y��;��.��>��yH��G�5����O8M�Y�O�=�� �G��a0�V�	M�f� Q��u��ߵ�������� ����'��$�  �bp;���� ��g�_�l�@�����@����C�����c��ey��S?333O����P���ñD/  �Ct`G�P ?fffO�>8���Ss	 k�_!xD�s{�O� IwS�'H;e#��/��j� F@� ��/o�� Dz ] ����I�q��y ܗ��� ��//�/�/K] �_]/o/�/�/�/�/�/ �?�?�??#?5?G?Y? k?}?�?�?O�OO�?g|�#O��O��� ��/	_���O�O�_ _0_B_T_f_x_2o�_ �_@o�_$o�_oo,o vo$%t:/&8B(�OPp\cҹ6��o �~ǯ���o��E?� �BPp?��ܴW���L� �����jH��gؠ�tPq�6�#������8�Gt�K߅���	��>���Gt�w���� ������+�=�k� �s���������͏�� ��ܯ'�9�K�]�� 9�����~�ɟ۟��� -�#��G�Y�k�}��� u���ů���lD�������2eC�U�Hg�yߊ�iϢ�2�� ��������� �2�D� V�h�of���Դ�� ����KMO	O	C�XO>G h�j"�4�a�X�}�ӴИ��������p�>�a��z��B�B\���>L5 \�<��{�<#�
�㲁p�����E,ϊ�����p������İ#@pA$�b�z�B� SB@�KJ���s���B�n�������t >�Hs�xi�*/�It$ C/-$��>�I
#/u'A �u//�/A/S&���+����%.��y��%��$敕�%�(4$�5�/�+;���.75>��H�C5��5��S58'M�Y_5��= {5��L��?�+	�/�?�? �?�7?O&O8OJO\O�nO}K�$CCSC�H_GRP12 �2����A�&� \���Xo��   O��`�lt �E�E ���A�__,_>_�2(U_C^����`Q�e?333��R����#D/  CаG�P ?fff��>���e�Y�Q�}� �Ojb�m����W�i� �o�o�o���2o�o<�E`F@ 8uDa�U�E`Dz�PYtDo�6�j6��� �o&o8oJo\o"��o �L�^��o�o��� ��&�4�f�$�6�W� ������ď֏����@N������f���� x�&8J\n� ����e�w�1������� ѯ������+���O� ��s��������u��`��ϣϵϿxȄ� ��ٳ.��i�'�#�� x�q�H��R<L���� ��8�W� �� ���4 ����J���sLV�����/�t�<���>����Ē� ����*�<�N�`�9� �ߖߨߺ��ߊ���� �&�8�J�#n��Y ����������"� �F�X�j�|�����^ ���������0B /f�����S/e/w/�%2�l�/�/�/�/=	�22?C?U?g? y?�?�?�?�?�?�?�d �nN1!Q|Y|Zqȝ �Y�Y�՟����i�O �O�O�O�FP� W��O�I�!AW-3�>�5�\_�S�H��iU�>L�P�Q�cB�<'#�
�`pi_RpE��V<B���@,0�U bA�U@� �T4�Lo��В�f Țeo��Ba�U �o�oBT�P>Ea�T�O�O�~C�It$ �$6>%��R
��wA}D������v!P+��=�`�.���l� Q�$敕|�(4$�܈�@�R�;��.���>��H�� Q5���Ѕ8M�Y܅(M=�P�� R�	�/�	&�?�*�c�N��� ������ǟٟ�Zo M|ؾ��  � I�b�T�b�PX�@�8J E�hd�v�����������<B�>��S,�?333(U`�)TlI�a�D/  CMGÿP ?fff(Q> amD,�L�D���� �L�TM(_"�P�,�  �!��?���bπ��F@ �Š��Hb��Dz6��Ġ����d�"ʳ!�/�) � p���������~�ܿ�� �ߺ�$�6π6�H�Z� l߂ߐ��߀����� ��� �2�D�V�h�� X�j���������^� ���ϔϦϸ������� |R�������	- ?Qu��� ���O��M/�0��/����)  5�i���.�_nC� �/����`��) e�" �d0a�f%`�E�ih!? k�Ph$)!��$z>�U��8 $$�^o�<�?�8>��� $�:P/ b/t/�/�/�/�/�O�/ �/??D?�OL?^?p? �?�?�?_�?�?�_ O O$O6OXOolO~OWo �O�O�O�O_�O�o _ 2_D_V_h_No�_�_w �_l�/����u�2>��.�@�R�c�B{�2v�����ÏՏ �����/�A�H�?� b��q�dةت�l$�(� (�r1��AC����:�1�V��d�pq�ݟP��q����Ia>����S}���5sť>�L���5o��Ty<#�
�Q�bpůd���8c�����Ia�e �a�|��`��@I��� ���Sd,�o۶$���{bLon{B�a�� G�h�z�]Ϟϰ�ckM��>��!�L�B��ړI�t$ �$m�>�"�
��N�AٔN����p��,�}�+��̞��.�����|�$�敕��(4$�x�՜߮�;��.��>��H�|�5{��,�8M�Y8���=��T�|�%qe��	�ߛ�������� ���#�5�G���\�4>Y�  (r� p�E��M��������� u���������x���ʘ���*��?3�33����ș��D�/  C�`G�P_ ?fff��>m� ɔ��	��_Vxy�C �����~���J\ }peX��d��j� F@ ��d��� Dz� $���p~���y �� ���/8B/? ?���_�/�/�/�/ �/�/?�?�?OF?X? j?|?�?�?�?�?O�O�OEOO�L�XO�0_ ��//&/8/>_آ _/_�_S_e_w_�_�_ �_go�_�_uooYo+o =oOoao�oY%�o/I[mw(�<O�p�c �k�!�~��Γ0)�  Ut�R�pt�P�� ��0Ɓ������j}��g ��t�qk�X�֎L�m�|t�ߺ�,�>�J�>���|tJ��� ������<�N� `�r���B�����̏ޏ ���ۯ&�8��\�n� ������n�ȟڟ���� �"�4�b�X��|��� ����į���������p�Gy��/�E�2@�xߊߜ߮߿�����2������1�C� U�g�y������ ��	�4	4
)̀M�	�	 xOsG�ϟW�i��������8���9�K�(O����� Q>�a��R R��!>L�j Q����<#�	
8��p!���Ea������� Q��@���X@�AY�b ��w��Bu�7�Jײ����B�A=������/��� >��}����_/6�Itk$ x/$��>�~	
X/�'A5��/R/�/xv/�&��+���5�.���$5��$�{��45(4$�@5��/
;;��.l5>���Hx5��5�=��58M�Y�5��=Q �5����?�+	 �/�?�?OGT?FO[O mOO�O�O��n�G  ��p� �L� U�E���A� _._@_R_�2i_W^�����`��e?33�3��R��$�XD/�  C�G�P /?fff��>�-� �ei�Q<����O�b} ����Wy��o�o�o�̵��Fo�o8�Y`F@ LuXa�U Y`Dz�PmtXoJ�j8k�K�=� �(o:o Lo^opo6��o�`�r� �o�o8�� ��$�:� H�z�8�J�k�����Ə ؏���� �b��"���z�4������: L^p����4y� ��E�����ӯ���	� ÿ-�?�ѿc������� ����ϵu���Ϸ����xȘ����c �G}�;�X&�υ�\� �Rq`������m� �� P�P ���#�i   ����J��2�`V�؂���/����>����Ħ���,� >�P�b�t�M��ߪ߼� ���ߞ���(�:�L� ^�7���m������ ����$�6�Z�l� ~�������r������  DV//z�@����g/y/�/�%2�l �/�/�/
?=�322.?W?i?{?�?�?�? �?�?�?�? t�nNE! e�Y�Z�ܝ�Y�Y� �ϗ��i�O�O�O�OVd� )W�O�I�!UWA3L>I�p_-pg�\��}U>L�P�Q�wB)<#�
�tp}_RY��VPB��L@D�U4bU�U@��TH�`o /����fܚyo3&+Bu�U�o�o @2Vh`>Ya��T_�O��CIt$� �$%6>��R
��A�D��(����v5P+���t�.������4Q$�=���(4$ܜ�T��f�;��.ȅ>���Hԅ4Q5����8M�Y��<M=@�P�4R��C�	:� S�>�w�b�������ɟ�۟���noM��  �]�(b�T �b`l�T�LJY�-hx��������0�ů��PB��R��S@�?333�<Ut�=T�I�aD/ � CaG�P ?fff<Q>%a�D@� `�X��(1���`�hM <_6�d�@��5�(�O���vϔ��F�@ �Ŵ��\b��DzJ��Ĵ���x�6��!�/�) ܄����� ��̿����ϼ���8� JϔJ�\�n߀ߖߤ� �ߔ�������"�4� F�X�j�|��l�~��������r����Ϩ� �����������R���� �/ASe ��-��� c�a/'�//%//����= I�i#� ��.�_~C��/��,� �`��= ,e2�dDa�f 9`�E�i|5?�P|$ =!#�4�>e��%84$�8�ro�<�?H>���4$Jd/v/�/�/ �/�/�/�O�/??*? X?�O`?r?�?�?�?�? �_�?�?�_O&O8OJO lO&o�O�Oko�O�O�O �O__�o4_F_X_j_ |_bo�_�_��_(l� 1/����u2R�0��B�T�f�w�V��2 ����ŏ׏����� 1�C�U�\�S�v��q�d ���l8�<�<�0rE� +�UW��!�N�E�j��d�p�������
��]a>�̯g}��8��Is٥>L"�	�xIoӒhy<#�
�Q�bpٯx���w�����]a�e�a�����`�@]�����g /d@�-o�8�տ�b`o�{B�a����[�|ώ� qϲ���wka�>��5��`�V���It$ Z0�$��>�6�
�b�A�b�
߄�.�@�ޑ�+�����.�����Ր�$敕��(4$��հ����;��.$�>��yH0吡5��@�O8M�YL嘝=	� h吢9qy��	�߯� ���������%�7��I�[�j��$CCS�CH_GRP13 2������&� �\�~E�y  <r���Y��a��� ��������+P��B0����>��?333����|ܙ�D/  C�`�G�P ?fff��>��ᔜ�	��_ jx��W�ĝ���� �����el��x��j2F@ %%01���2Dz� F$�1#/��#���y �%7I? mw/9?K?���_�/ �/�/�/?!?S?O#O DO{?�?�?�?�?�?�?��?;O�O�OzOSO\� �O�e_/%/7/I/[/ m/s_�R_d_o�_�_ �_�_�_�_�ooo�o <o�o`oro�o�o�o�%���/~���(� qO�p�cɠ�V�� ޓe^�5U�)�9R�p ����%Ġ�Dƕ��� �j���g!��t�q���� �`�9���t��οxa�s��>����t �����)�;�M� &�q�������Տw�ݏ ���%�7��[�m� F�������ǟ韣��� ��3�E�W�i����� Kϱ�ïկ���߿� /��S���|�@�R�d�z�2��߿����������2�0�B� T�f�x�������� �����>�i	i
^� �M�	�	���O�G���@����������=�m�@n�����.�ڱ>"qI��@R5R��V>L� �ƿP���O<#�
m�M�pV���2U����)����ڱ��u.��@ �A�!r9�Ϭ��B��@l�JR�ݿ��BN� vr��/�//A/��� >2������/^k�It$ �/$��K>��
�/�'Aj���/�/?�/�& +�{��M5.���Y5�$敕i5(4�$�u5-??;;��=.�5>��H�5�5���58M�	Y�5�=� �5���?;	?,OOPO;G �?{O�O�O�O�O�OG����n�G   ��6p��� EU-U %�2QQ_c_u_�_	B(�_�^)��+p�u?333MRY���D/  C:�G�P ?fff>�Z�u9i1aq��� 
_�b9}A�g=y/ �o�o���{o�oO<mʎ`F@ �u�a�U5�`Dz#`�t�o�Qz�р�r� �]ooo�o�o�ok��o �����#m�#�5� G�Y�o�}���m���� ׏�����1�C�U�@��E�W�֟��i��� K��o����� ϯi����z����� �,�>���b�t�Ϙ� 꿼�ο��<��u:�` ���������͟ �"Ø�G��pލW� �Ϻߑ�b���� �Ң����U� �XǞ U���J��g���V���?K��<����>������ =�O�a�s߅ߗߩ߂� �������1���9�K� ]�o���l���� �����#�E��Y�k� D������������� 1CU;y� d/���
ߜ/�/�/�%2+|	??-???P=	//h22c?�?�?�? �?�?�?�?
OO.O5t ,~ONz!��Y�Z�� ii	"��./0y�O �O'__CV�� ^W��O�I�!�Wv3��>�~��_@-����"#�U�>L�P�Q"�BA)<'#�
��p�_QRp���PV�B����@uy�Uib��U@6� �T}o@/��f ��oh9[+B��U �o4UgJ��P:`>�ad9_/_��C�It$ 	�$Z6>%�b
�;�A�D;���]���jP+��=̩�.�����iQ�$敕Ņ(4$��х����;��.���>��H	�iQ5����8M�Y%�qM=�PA�iR!R�x�	o���s������ ן����"�4��oIM|!�F�  " ��]b2d�b:`�����J ��bh����ѯ�e����讅B���cu�?333qU��rT�I�a�D/  C�GÿP ?fffqQ> Za�Duŕ����C(f� 0͝Mq_k���u7� I�j�]EO׿Qϫ���F@ ���Q��b�Dz��������k��!�/�) � ��˿ݿ����%�/� ���m���ߑߣ� �������������3� E�W�i�{������ ����2�����E��� ��������%�+ �R
�@Rdv ��T��b�F *<N�FՖ/\�06/H/Z/d��)�r  ~�iX�/�.�_�C/ ?��a�p��r ae=2 �dyavn`�E�i�j? ��P�$r!X�E4�>9e�Z8i$m��oL+O7H>���i$7J�/ �/�/�/�/�/?�O)? ;?M?_?�?/_�?�?�? �?�?�?�_O%O�_IO [OmOO�O[o�O�O�o �O�O_!_O_E_i_ {_�_�_�_�o�_�_� o]l4/f/�
��2��2��e�w��������Ă2������� 0�B�T�f�x����Ĉ� ���q�d!�!�|m�q� q�erz�`����D�V���z����d%���&�P8�<��҃��>����}����~s�>�LW�>�~o��y<#�
%arp�����8N��������e �a-�Ų�`E�@��F� ��ddu�bo$�m�
��b�o�{Bq.�*� �ϱ��Ϧ����Ϭk���>�j�����L�#�I�t$ e�$��>�k�
Eߗ�A"���?���c�u�Ơ+��̞�.����š$�敕!�(4$�x-�����;��.Y��>��He�š5{��u�8M�Y��͝=>���Ţnq����	���������A�3� H�Z�l�~�������}>��  qr� ����9�����ݚ�� ��	-?��VD����s��?3�33ͥΤ�E�D�/  C�`G�P_ ?fff͡>�� ���	�)o�x��� ���ͯ���ϓ� ��e��3�/%zFF@ 9%E��FDz� Z$E7/	/p�X�8�*� � '9K]#?��/M? _?��%o�/�/�/? '?5?g?%O7OXO�?�? �?�?�?�?�?OOO�O_�OgO!\��O/y_ '/9/K/]/o/�/�_!� f_x_2o�_�_�_�_�_ �_�oo,o�oPo�oto �o�o�o�o�%��/����(ȅO�p�c Pɴ�j(�E��yr� IU�^�MR�p����Z� ձy�ʰ=�=�zƏw V���q�������M���t���u�����>����t���� �+�=�O�a�:����� ����鏋����'� 9�K�$�o���Z����� ɟ۟�����#���G� Y�k�}�����_�ůׯ �����1�C��g������T�f�xߎ�2@������������ �2�D�V�h�z�� ������������ 2�R�}	}
r��M�	�	 ���O�G�������������Q�������(��B.�9�>6q]���TRIR��j>L� �ڿd���<#�	
��a�pj	FU��=���9�-�1��!B��@�A�5r M�����B����Jf ���Bb�����///C/U/�� >�F������/�Itk$ �/$�>��	
�/�'A~��/�/?x�/�&" +���a5�.���m5!$�{��}5(4$܉5�A?S;;��.�5>���H�5!5�=��58M�Y�5)��=� �5!��
O0;	 '?@O+OdOOG�?�O�O �O�O�O�O[��n�G  ��Jp ��� YUAU9�FQ e_w_�_�_B�_�^=���?p�-u?33�3)aR*m��D/�  CN�G�P /?fff)>n� -uMiEa����_�bM} U�)#gQy-/�o"����o	c�ʢ`F@ �u�a	eI�`Dz7`�t�o�e#z8�є߆� �qo�o �o�o�o��o����� %7��7�I�[�m��� ��Ï���������� !�3�E�W�i���Y�k��ß}����_կ� ������}¯ ԯ����
��.�@�R� �v���Ϭ���п� ���P��uN���� �����*�6ì W�τޡk����ߥ� b���*��Ҷ1 �&���i�"�lǲ  i�*�Z��{���V�!�%?_������>���!���Q�c�u� �ߙ߽߫ߖ������ �E���M�_�q��� ��������%� 7�Y�m��X���� �������!3E WiO��x/�@��߰/�/�/�%2?| ?/?A?S?d=C/|22w?�?�?�?�?�?�? OO0OBOIt@~cN�! ��Y�Z�%�)i)i" 2��B/Dy�O_;_2_WV�� rW�O�I�!�W�3J>���_T-p����6#�U>L`��Q6�BU)<#�
��p�_eR��/dV�B��J���U}b��U@J��T�©o T/-��f%��o|Mo+B��U�oHi@{^��dN`>�a�"dM_C_��CIt$� �$n6>�#b
�O�A�DO��q���-�~P+��̽�.����Ʌ}Q$�=�م(4$�兝�ޯ�;��.�>���H�}Q5���-�8M�Y9��M=@�PU�}R&!f���	�� ����������� ���$�6�H�W��$CC�SCH_GRP1�4 2����y�&� �\m.2�p)  )"��qbFd�bN` ֥���Jávh������y�/���B���<+c��?333�Uޢ��T�I�aD/  C��G�P ?fff�Q>na�D��ʹ± �W(��D©ͱM�_�� �ɉl�~ϟ�qYO��������F@ `�����b�Dz�� 3����Ϡ�1�/�) �� ��$�6� ��Z�d�&�8�ϴ�� �������� ��@��� �1�h�z������ ����(�����g�@����z���R ��$�6� H�Z�`�R?Qu ������� �){M_q���{ժ/��k/}/�/���^�� �y��C/> �_�CR/K?"��p& � uer2t�a1v�`�E �i��?�`�$�!��@z4�>Me&��8�$���oNL`OlH>��� �$lJ�/�/�/??(? :?_^?p?�?�?�?d_ �?�?�? OO$O�_HO ZO3o~O�O�O�O�O�o �O�O�o _2_D_V_�_ z_8�_�_�_�_�_�o 
oo�@o�li/�/-�?�Q�g�2�̚�����$Џ����2�� /�A�S�e�w������� ���Ľ����+tV�V� K|�������r��������y�������Ԧ*t�Z��[�m�q����a>!6��}-"�sC�>L��s��o=���y<#�
Za:rp�C��������au
qb���pz�@��{�"&���d��oYƢ�?��b�o�{B ;qc�_����������.��k˰>���ʯ�����X�It$ ��$��>���
z���A�W���t��ߘߪ���+����:�.����F���$敕V�(�4$�b��,�;�{�.��>��H�����5����8M�Y���=s������q��	�	 ���=� (�v�h�}����������4�ڝ���  �r# �ôn�˰2 ��>PbtP��y�� ��%?333�:�|F�z�D/  C'p�G�P ?fff�>�G�%&^o �x���&-.���*) �����e֟h�x</Zz{F@ n%0z�"�{Dz�$�zl/>/���m�_� �J\n��X? ��/�?�?�/Zo? "?4?F?\?j?�?ZOlO �O�?�?�?�?OO0O�BO�O2_D_�O�OV\� �O8/�_\/n/�/�/�/ �/�_V��_�_go�_�_ �_oo+o�oOoao�o �o�o�o�o�o�o)�%�'��/����(� �O�s�����]�z� H����~U����R� �΂��
�����r�r� Bz��Ew��B����ք T�ʵ���t��8�x����Ș>����t Ț*�<�N�`�r����� o���̏ޏ�����&� 8�J�\�n���Y����� ��ڟ����2��F� X�1�|��������֯ ������0�B�(�f� x�Qߜ�����ߛ�����2,����,�=��U�2P�y�� �����������	�� "$.<�gчĲ	�
�� �M��_�G�)@����0����@K������wc�#�>kq�-݉R~Rӟ>L� �ϙ�.�O<#�
����p��>{U��=r����#�b�f��Vw��@ #Q�jr�-���R�@��J�U�&�H�B�� ��!/B/T/7/x/�/=�'>{�&�/^��It$ �/$G�K>��
�/(7A���(?�/J?�/6W +�{�̖5.����5�V$敕�5(4�$ܾ5v?�;;��=.�5>��H�5V�5��E8M�	YE^�=� .EV��?Oe;	\?uO`O�O�G �?�O�O�O�O_!_��6�~3W   �pJ�'�UvU n�{QO�_�_�_�_RB(�_�^r��tpbu?333^�R_����D/  C��G�P ?fff^>G��bu�iza��0� S_r�}��^Xg�yb/ $6WJ�2��o>�<���`F@ �u�a>e~�`Dzl`�t�o���Xz���߻� ܦo�o�o�o�o�� �ޏ��Zl��l�~� ������Ə����ȟ�  �2�D�V�h�z�����@������������2� �
����� �� ����	�ÿ-�?�Q� c�u���Aϫ���O�� 3���)�;υ�3���`I�#�5�G�Q��� _�k��EW�Ϲ���� 
��ڥNb�ޢ_�N *��f
&[����� W��� ��_�EZ2��&�VG�V�Z?��<�$�>���V�$� �ߘߪ߼��������� �(�:�L�z���� ������� ��� 6�H�Z�l���H���� �������<2� Vhz����� �/�J!�S��/�/	?52t|R?d?v?�?�=	x/�22�?�?�?�? OO/OAOSOeOwO~t u~�N�!�ij,Z� ^i^iR"g�M�w/yy1_ C_p_g_�V�0�W�_%Y)1�W�3>����_�-�ڢk#�U�>LD`+ak�B�)<'#�
�p�_�Rpץ;/�V�B��@��e�b�2e@� 3d���o�/Qb�Ov Z��o���+B�e }�������`>�aWd�_x_9�S�It$ R�$�6>%�Xb
2���AT���,���P�b��P+��=��.������Q�$敕�(4$���ҏ�;��.�F�>��HR��Q5���b�8M�Yn��M=+`���R[!����	��џ������.�  �5�G�Y�k�}��o�M|jΏ�  ^" ���b{d&r�`�ҥ�J ס�h����,���C��1��B���`c��?333�U�T�I2q�D/  C�GÿP ?fff�Q> �a�D��޹ֱ�(�� y����M�_���ɾ�� �ϳϦ�O Ϛ���*3�F@ &�2����b3�DzȰG�2�$���ϴ�E1%?9 � ��&�8�J��n�x� :�L���������� ���"�T��$�E�|� ������������<� ����{�T������ f�&�8�J�\�n�t bSe���� ����=� as������/��0/�/�/���r��  �=y��W/>2o�Cf/ _?6��Kp:� �e�2 Gt�afv�`*U*y��? �C`�$�!���4N�e:��8�$���obLtO�H>����$�J�/ �/??*?<?N?'_r? �?�?�?�?x_�?�?O O&O8Oo\OnOGo�O �O�O�O�O�o�O_�o 4_F_X_j_�_�_L�_ �_�_�_�_�oo0o	� To�l}/�/A�S�e�{��2�̮���ҏ�����2�1�C�U�g� y���������ӟ���� ���?tj�j�_|���� ���r������ɍ���̯ï�>tn��o�P����/���a>#!�J��}A6�sW�>�L�����oQ��y<#�
naNrpW���38���*����au qv��/p��@�� "":���d��omƶ�S�r�o �BOqw�s� �������0�B��k߰�>3���ޯԯ��l�I�t$ ��$��>���
����Ak��߈���߾��+��̞N�.���Z��$�敕j�(4$�xv�.�@�;��.���>��H���5{����8M�Y���=������q���	�-��Q�<���|� ����������H���>��  �r7  �״��߰F.&�3 �Rdv�
���*��, ��%?3�33�N�Z���D�/  C;pG�P_ ?fff�>�� [�%:2ro�x� :-B��>)��� /u�|�P/nz�F@ �%��6��Dz$�$��/R/p*����s� �^ p���l?��/�? �?/$/no$?6?H?Z? p?~?�?nO�O�O�?�? �?O O2ODOVO�OF_X_�O�Oj\��OL/�_ p/�/�/�/�/�/�_j� �_�_{o�_�_	oo-o ?o�ocouo�o�o�o �o�o�o=�%;�?���	8��O�#s �����q���`���� �U���R��₣� ��������Vz�Yw ��V�����h�޵�����LϾ�Пܘ>����ܚ>�P� b�t���������Ώ�� ��2�ԯ:�L�^�p� ����m���ʟ��� � �$�F� �Z�l�Eϐ� ����Ư��ꯨ�� � 2�D�V�<�z���e߰������߯�����2@,,
��.�@�Q�0�i�2d�������� ������/�6$-.P� {ћ��	�
��] 
�_W/�1)����(D����_����(�ыw�7�>q��AݝR�R#ӳ>L�� �#ϭ�B�<#�	
ʱ��p�R�U��Q����7�v�z��j���@7Q�~r �A�	�R��Z�i�:�\�B����5/�V/h/K/�/�/Q�;>��:0�/��Itk$ 
?$[�>�	
�/<7A��<?�/^?x?6k +��̪5�.����5j$�{���5(4$��5��?�;;��.�5>���H
Ej5�=�E8M�Y&Er��=� BEj�SOy;	 p?�OtO�O�G�?�O�O��O_#_5_D[�$C�CSCH_GRP�15 2����fQ&� �\Z�]�  ғp^3� ;�U�U���Qc�_�_@�_ofBo
n����pyvu?333r��Rs���D/  �C��G�P ?fffr>[��vu�i �aοD؈_1r�}��r �g�yv/Yk�^�F���os���pF@� �uqse�pDz �` ����z������ ��o�o�o #�GQ��%��� ʿ����ŏ׏���-� ����U�g�y����� ����ӟ�ïկT�-�笸g��?���� #�5�G�M��,�>��� b�t���������v�� ���h�:�L�^�p� ��h���~�X�j�|߆��K��Р��zW0� �����?�8���b  ���b_��z&o ����ʌ���� �ԔрzZg���:f|���n?�;�M�Y�>�����Y���������� �'� K�]�o��� Q������������ 5�G� k�}������� }�����1C qg%/����� ��	�/-V߈�?,?>?T52�|�?�?H�?�?�=�/�22�? 
OO.O@OROdOvO�O �O�O�t�~�N�!$Ci Cj8,���i�i�"���� �/�yf_x_�_�_�V$G0�WH_ZY^1g�3�>��#o�-���#0e>Ly``a�<*R�)<#�
G'"�p0o�R�p/�VR�����Oe�b ge@��hd���/� ���Fv��,���+B(!PeL����	����`>q�d�_x�_n�ESIt$ ��-$�6>��b
g���ADT��a�ۏ�����P�+���'�.��y�3��Q$敕C��(4$�O���;���.{�>��H����Q5����8'M�Y���M=``���R�!П��	��� *��c�U�j�|�����ಯ!�M��ħ  �"��b�d[r�` ���J��h+�=�O��a��x�f�R��<�c��?333�U'���T3YgqD/  C� G�P ?fff�Q>�a4T���� K�(䯮��]�_� ����������OU����)�G*h�F@ `[�g�ϵrh�Dz�� |�g�Y�+���z1Z?L9 �7�I�[�m�� E�ϭ�o������G ���!�3�I�W��G� Y�z������������ �/�q�1����C���%ߛI�[�m�� �ߣߩCb��T� ����<N �r�����/���?�ߴ/�/�/��ȧ�� �ry֧�/J> go1S�/�?k߲�po � �e�2|t�a�v�`_U _y/*�?2'x`/4�!֪@�4AN�eo��8�$��%�L�O�H>��� �$�J?)?;?M?_?q? �?\_�?�?�?�?O�_ O%O7OIO[OmOFo�O �O|o�O�O�O�O_�o 3_E_i_{_�_�_�_ �_��_�_oo/o Soeo>��o�l�/�/v�������2�����$�*�	�B�2=�f� x���������ҟ��� ���)�T�tt���� �|�����r������
�¯ԯ����st���8�������d�P�q>X!��vk�s��>Lհ���o����<#�
�a�rp���+�h�*�_���qOuSq��C�dpõ@ĴW"o���d���o������Br5�B �q�����/�A�$�e�w�*{�>h���	���ߡ�It$ ��$�4�>��
���A�����7�����D�+���̃�.������C�$敕��(�4$ܫ�c�u�;�{�.��>��H���C�5����8M�Y��K�=���C��q,�R�	I�b�M��� q�������������}�#��   �rl 7�ķ��{ c[�h<ȇ���P?���_��a �O%?333K��L�|����D/  Cpp�G�P ?fffK�>4���O%og�o �@
"o-w�K�Es) O�/#/D/7u��+/x�/�z�F@ �%0�+k��DzY�$���/�/E*ց���� ܓ�����? �	?�?�?G/Y/�oY? k?}?�?�?�?�?�O�O �OOO1OCOUOgOyO��O�O{_�__�O�\� _�/�_�/�/�/�/�/ �/o���_�_�oo,o >oPoboto.�o�o< �o �o(r 5�p�6?�"�4�>8� _L�Xs��2���ÿ ������U;���RL� ;����S���H����� �zD��w԰��L�2
� ����4�C�G��x���>���C� �s���������͏ߏ ����'�9�g�	�o� ��������ɟ����� ؿ#�5�G�Y�{�5Ϗ� ��z�ůׯ���)�� ��C�U�g�y���qϯ� �����7��@��������2a,?�Q�c�u���eߞ�2������ ����
��.�@�R�d� k$b.�������	�
�� G]KK?�T_:Wd�f)@0]Ty����@� 	����l�>�q�v��R�RX��>L1X���w�O<#�
����p����U(߆�����l��ů����@ lQ �r�v�>�OR<�@�GZ���oϑ�B�� /j/�/�/�/�/�/��p>�Doe&?^��It$ ??$��K>�E
?q7A���q??�?=?O6� +�{���5.����5ޟ$敕�5(4�$�E�?�;;��=.3E>��H?E��5��OE8M�	Y[E��=wE�H��O�;	�?�O�O�O�G O_"_4_F_X_j_���W~|W   K��p�h"p�U�U ���Q��_�_oo�B(0on����pM�u?333��R����!D/  C��G�P ?fff�>����u�i�a�y� �_fr�}����g�y�/ m���{���<�� pF@ �q�e� pDz�`4�����z2��� ��o%7��[ e�'�9�������Ǐ ُ���A����2� i�{�������ß՟�@)�ׯ�h�A����{� �S���%�7�I�[� a��@�R��v����� ����п����Ϙ�*� |�N�`�rτ���|���`��l�~ߐߚ��_� �д�*)�WD���� S�L�#��b8 '��З s�4$�S&�)�� ����0�ԨюZ{���o'f����?�O�<a�m�>�����m� ��������)�;� _�q�����e���� ����%��I�[�4 �������������� �!3EW�{9/ ������ �/A�jߜ�.?@?R?h52�|�?�?�?�?�=	�/�22�?O0OBO TOfOxO�O�O�O�O�t �~�N1,$WiWjL,�� �i�i�"�����/�yz_ �_�_�_�V+$[0�W�\_nYr1gC�>��7o�-.�#��#De�>L�`ta�>R�)<'#�
[;"pDo�Rp ��/�VR���@%!ce�b {e@ȡ |d�'�/����Zv ��@���+B<!de `�����/���`> q�d�_�_��YS�It$ ��$�6>%��b
{�͇AXT͏�u�����P+��=�;�.���G��Q�$敕W�(4$��c��-�;��.���>��H���Q5�����8M�Y��]=t`ӕ�R�!�
�	���>�)�w� i�~�������Ư5�M|��ا  �" $��b�dor�`3��Z  ��h?�Q�c�u������z�R���c�?333e;�dGY{q�D/  C( GÿP ?fffa> �aHT�'��_�(�� ��'�/]o��+���� ������Oi���=�[*|�F@ o�{��#r|�Dz���{�m��?��ʎ1n?`9 � K�]�oρϓ�Y���� ������[�#�5� G�]�k��[�m����� ��������1�C��� 3E����W���9� �]�o߁ߓߥ߷߽ Wb��h��� ,�Pb��� ����*/��(?��0�/�/�/��Ȼ�0 #�yꧠ/^>{oES�/ �?�p�0�e�2 �tq�v psUsyC*�? F'�`C41��4UN�e���8�$��9�L�O�H>����$�J+? =?O?a?s?�?�?p_�? �?�?�?O�_'O9OKO ]OoO�OZo�O�O�o�O �O�O_3_�oG_Y_2 }_�_�_�_�_�_��_ oo1oCo)goyoR� �o�l�/�/������ą�2���	��-�>��V�2Q�z������� ԟ���
��#�� =�h��t�����|��� ��r����֯���1��t��L���Pʩ΁x�d�$q>l!���.�����>�L�б��/�<#�
�a�rp��?�|8�>�s���$qcu gq��W�xp׵@$ش k"��.��d�o������Vr'I�B�q���� "�C�U�8�yߋ�>{(��>|���'���ߵ�I�t$ ��$H�>���
��)�A��)����K����X�+��̞��.�����W�$�敕��(4$�x��w��;��.���>��H��W�5{���8M�Y�_�=а/�W� �@�f�	]�v�a����������������"1�$�CCSCH_GR�P16 2����S&�� \G�/J�  �� K� � ��(���o��Pȼ����S�	�s���u �c%?333�_��`�����D/ � C�pG�P ?fff_�>H���c% ���o1�u"�-�� _�z�)c�F/X/y/Ku�3��`/�/�z�F�@ �%�`��Dz�4��/�/z*�ʏ�� ���� �/�?4/>? OO|/ �/�o�?�?�?�?�?�? O�O�O_BOTOfOxO �O�O�O�O_�_�_A__�\�T_�/,o�/�/ �/?"?4?:o��o+o �oOoaoso�o�o�oc �o�oqU'9K ]�U5��k?E�W�i�s8�8_���s��g �ێ׿��,�%��Up �� b��O�L���g�� \�ϥ���zy��w��� ��g
T�Ҟ'� i�x��[��(�:�F�>���x�F�����̏ޏ �����8�J�\�n� ��>�����ȟڟ��� ׿"�4��X�j�|��� ��j�į֯������ 0�^�T��x������� ����������l�C� u���+�A�2�,t��������2 ����	��-�?�Q�c� u������$�.����� 00%�|]��t҉_ oW�ߛ)Se����4��5G	K��
����>�q��b8�R��>LfMx����<#�
4��p��U]߻����������<���T@�QU�r /�� sĄRq�3&|Z/�¤���B�=9/�/�/�/ �/�/?�˥>�y��[?2It$ Zt?$��>�z
T?�7A1�?N?�?r?�6�� +���E.���� E�$敕0E(4$�<E�?K�;��.hE>��yHtE�5���EO8M�Y�E��=M �E�}ѽO�;	�?�O �O_WPOB_W_i_{_��_�_/���~�W  ���p��H" �e�U���Q�o*o@<oNo�BeoSn����py��u?333��b� 	T!D/  �C�G�P ?fff�>�!�u y �a8Ϯ��_�r �� �g��/����Ű��B��4�UpF@� H�Tq�e�UpDz �`i�TF���zg�G�9� �$6HZ l2����\�n��� 4����� �6�D�v� 4�F�g�����ԟ� ��
��^�����v�0�������6�H�Z� l�~�����0u���A� ����Ͽ��Ͽ�)� ;���_ϱσϕϧϹ� ߱��Ǐ�߳���ψȔ�����_)�Wy� 7�T�߁�X��bm  \������i$��&� LL)����e��р�Z��.��\f������?/������>����Ԣ���(�:�L� ^�p�I�������� � ��$�6�H�Z�3 ~���i�������� � 2/Vhz� ��n/���
 /@R+?v�����c?u?�?�52�|�?�?H�?OM�//B2*O SOeOwO�O�O�O�O�O �O�O�t�~^A1a$�i �j�,ح�i�i�"�˧ �/�y�_�_�_�_
f`$�0%g�_�Y�1Qg=C�>E�lo=c�X��#ye>L�`�a�<sR9<#�
�p"�pyobU��/fLR���<%@!�e0rQ �e@���dD�\?� ���vتu/" /";Bq!�e���.��R�d�+p>Uq�d ox�_���SIt$ Џ-$!F>��b
���A�T���$�Ώ��1`�+���p�.��y�|�0a$敕���(4$ܘ�P�b�;���.ĕ>��H�Е0a5����8'M�Y�8]=�`�0b�!�?�	6�O�:� s�^�������ůׯ����j]���  �"Y�$r�d�rp h�P�HZU�)xt��������,�����LR�N�<�c<�?3338ep��9d|Y�qD/  C�] G�P ?fff8a>!q}T<�\�T� �
8-���\�d]8o2� `�<����1�$%_����rߐ*��F@ `�հ��Xr��DzF� �԰Ϣ�t�2��1�?�9 ܀ϒϤ϶��� �����߸���4�Fߐ F�X�j�|������ ��������0�B�T� f�x���hz������n���ߤ߶��� ������b��� +=Oa/�� )/�/��//_/��]?#��/?!?+����90E#�y��/�> �ozS�/�?�(��p� 90(uB�t@q�v5p�U �yx*1O{'�`x491�@D�N u��!H044��n�L�O�H>��� 04�J`?r?�?�?�?�? �?�_�?OO&OTO�_ \OnO�O�O�O�O�o�O �O�o_"_4_F_h_" |_�_g�_�_�_�_o o�0oBoTofoxo^ �o�o���o$|�/-?��я���2N�,�>�P�$b�s�R���2���� ��ӟ���	��-�?� Q�X�O�r����t�� �|48�8�,�A'Q��S���J�A�f��t�쀁���������Yq>�!ȿc���E�յ>L��EϢ�d�<#�
�a�rp�տt���s�����Yq�u�q���­p�@YĠ"��c�+t<�)��4
�ϋr\~�B �q����W�xߊ�m߮���s{]�>��1�\�R����It$ ,�$�}�>�2�
�^�A��^���*�<捰+������.�����匱$敕��(�4$�����;�{�. �>��H,�ތ�5��<�8M�YH���=�d���5�u���	������� �����!3EW���l�D.i  8�� ��U� �]�� ���������P������ :��%?333�����|ة�D/  C�p�G�P ?fff��>}�٤�%���o f��S"�-������) ��Z/l/�/�uh��t/x�/�z F@  50!t�� Dz�!4�/�/�/�*���� ��� //$/�? H/R?O&O�/�/�o�? �?�?�?�?�?.O�O�O _VOhOzO�O�O�O�O��O_�_�_U_._�\� h_�/@o�/ ??$?6? H?No�-o?o�ocouo �o�o�o�ow�o�o� i;M_q�i5���?Y�k�}��8� L_���s�{1��� ֣@�9�e�%�b�� ��`�!Ԝ�@֑��� �z���w�Ԅ��{
h� �\�}�������x<�N�Z�>����� Z���Ώ�����(� �L�^�p�����R��� ʟܟ� ���6�H� !�l�~�����į~�د ���� �2�D�r�h� &ߌ�����¿Կ���� 
���.π�W����-�?�U�2�,�����������2���� /�A�S�e�w������� �$�.�����DD9� �]���ҝ_�W�߯)@gy����H�@�I[	_�	����>�q$��bb��1>Lza��+��O<#�
H�(�p1��eq�����������P�	�h@ �Qi�r/�߇ĘR��@G&�Z-/�¸���B)� QM/�/�/�/�/
??�˹>!���o?^FIt$ �?$��K>��
h?�7AE��?b?�?�?�6� +�{��(E.���4E��$敕DE(4�$�PEOK;��=.|E>��H�E��5���E8M�	Y�E��=a�E����O�;	�?_�O+_W dOV_k_}_�_�_�_"/����~�W   �����\"� ee  
a�,o>oPobo�B(yogn����u?333�(b�4	�h!D/  C�G�P ?fff�>�5�uyqL��� �_�r���g��/ �������V�*�<H�ipF@ \�hq�e"ipDz�`}�h�Z�,��z{�[�M� �8J\n�F�� ��p�����H���� "�4�J�X���H�Z�{� ��ğ֟�����0�@r� �2�����D��į &���J�\�n������� ��D����UϿ�ѿ� ������=�O���s� �ϗϩϻ����Ņ�`ۏ�������Ȩ� ����s)�W��K�h2 �ߕ�l��b� p���� ��}$��&�``)0� ��3�y0����Z��B��pf�����?&/��<����>����Զ� �*�<�N�`�r��] ����������&� 8�J�\�n�G����} �������� �4F /j|�����/ ��0/Tf ??������w?�?�?�52��?�?OO+M	
?CB2>OgOyO�O �O�O�O�O�O�O	_� �*^U1u$�i�j�,� �i�i�"��ߧ	?��_ �_o�_ft$�09g��_�Y�1egQC!>�Yрo=w�l��#�e�>L�`�a��R9<'#�
��"p�o,bpi��/+f`R��!@P%T!�eDre �e@� �dX�p?�����v 쪉C"/6;B�!�e ��0�B�%�f�x�++p>iq�do
oˏ�S�It$ �$5F>%��b
ď�A�T�ྏ8���E`+��=̄�.�����Da�$敕��(4$�ܬ�d�v�;��.�ؕ>��H�Da5�����8M�Y �L]=�`�Db�!-�S�	J�c�N���r������ǯٯ�������$CCSCH_G�RP17 2����@�&� \4>��79  �"m�8r t�rp����\Z��=x ����Ϳ߿@����`R��b��cP�?33�3Le��Md�Y�qD/�  Cq G�P /?fffLa>5q�T PՑɉ��8b��p� x]Log�t�P�3�E�f߀8% _��Mߧߤ*��F@ ����M�lr��Dz{������ߩ�g�8�1�?�9 ܵ��� ��������!�+����� i�{ߤ{������ ���������/�A�S� e�w�����������.��A���� �������!�'�b �<N`r�� P/��^/�B//&/ 8/J/�/B�q?X�2?D?V?`��%n0z#�y T�
?�>�o�S?O� ]��p�n0<u9B�tTq �vIp�U�y�*fO�'�` �4n1T�AD�Nu�VH�e4H��\'_3X>���e43Z�?�?�? �?�?�?O�_%O7OIO [O�O+o�O�O�O�O�O �O�o_!_�oE_W_i_ {_�_W�_�_��_�_ ooKoAo�eowo�o �o�o��o�o��Y|@0?b?���.�2�� a�s�����������2�������,�>� P�b�t����Ԅާ�ҁ �t���im�m�a� v\����@�R��v����t!���"�4�8��Γ�q>�!����p��z�
�>LS��:�z���<#�
!q�p
ϩ��J���ݢ���q�u�q)����pA�@�B��"�� ��`tq^ �i
��r���B�*�&ߌ߭�@�ߢ����ߨ{��>���fđ���H��It$� a�$��>�g�
A��A���;��_�q�°+����.�������$�=��(4$�)������;��.U�>���Ha���5���q�8M�Y}�ɭ=@:�����j�����	�� ������=�/DV�hz���$CC�SCH_GRP1�8 2�����&� �\��v/��  m�� ��5Ғ� ٪��&8J�\��saݢ�� <o��%?333ɵ"�ʴ�A�D/  C��pG�P ?fffɱ>����%)! %����"�-��ɿ� �)�߰/�/�/�u��P/��/$?!�c F@ `V5b!���c Dz� w4b/T?&?�*T�4�&� �2/D/V/h/z/ @O�/�?jO|O�/�/! �?
OO.ODORO�OB_ T_u_�O�O�O�O�O_ _*_l_o,o�_�_>l��_ ?�oD?V?h?z? �?�?�oo�oO�o �o�o�o�7I �m��������5��?����ӏ�8Ȣ_��sL����E� A������fe�Z�jb 뀹Ŷ�V���u���9� 9�*��-�R�*���
@��<���jӘ�����ϒ�����>��� ℰ��$�6�H�Z�l� ~�W�����Ɵ؟��� � �2�D�V�h�Aό� ��w�¯ԯ������ .�@��d�v�����ȿ ��|������*�� N�`�9���̭�ߏq�����2 <�����$�%��=�28�a� s��������������� 
4>$O�oԚ� ���]�����_�W�9����n����3��	��_K��>S�z�qbfb���>L���ρ��<#�
��~�p��&ce��%Z���J�NѦ>"_о@a�R�j/����R��ϝ&�Z�/=��0�B ѧ�/	?*?<??`?r?%� >c!���?�It$ �?$�/�>��
�?GA��O�?2O�?�6?+����~E.�����E>$敕�E(�4$ܦE^OpK;�{�.�E>��H�E�>5���E8M�Y�EF=�U>��'_MK	DO]_H_�_ lW�O�_�_�_�_�_	o�k�$CCSCH�_GRP19 2����:a&� \.�|�1�  �� g�2"$�" �eeV
 �a7(�o�o�o�o:R�o��nZ�\��J�?333F�bG�	�!�D/  Ck�GÿP ?fffF> /!�J��y�q���\o �j�rFawn�J?-� ?�`�2��G������pF@ Ӆ�qGuf"�pDzup��я࣏a����� � ��������%� ���c�u���u����� ����ϟ���ѯ�)� ;�M�_�q�������� ����(�����;��� ���ӏ���	��!� � ����6�H�Z�l� ~ϐ�Jߴ���X���<� � �2�Dߎ�<�k�R�0,�>�P�Z���h� t��)Ng����� ��Wr� �h�6%3� �$N!�&C ��)��`� �����h�Nj;���%�fP�_�BO|/!->���_�-
�� ������������� 1�C�U���%������ �������	�? Qcu�Q/���/ ��E;�/_ q����/���? /S,*�\��? OO(E�2}�[OmOO�O�M�?�B2�O�O�O__ &_8_J_\_n_�_��~� �^�1�$yz<c�gy gy[2p�V��?��:oLoyopo�f�$@�goP.i2A�g�C�!>����o�=��t3u>�LMp4qt/�R�9<#�
!�"p�b�8D?�f�R���!�% �!#u�r� ;u@��<t ����?Z$k�X/�c� ��"�/�;B�!$u � ��������ݏ+�p�>�q`t�o�oB�cI�t$ [�$�F>�ar
;���Ad��5��Y�k��`+��̞��.�����a$�敕�(4$�x#�۟�;��.O��>��H[��a5{��k�8M�Yw��]=4p���bd1��ʛ	��گů���7�)��>�P�b�t������$�CCSCH_GR�P1A 2������&�� \�>p߮9  g2�Яr�t /��p����Z��x π2�D�VϷ�m�[��R����is��?333��e��di;�D/ � C� G�P ?fff�a>�qd�� � �/�8ٿ�����] �o����Ǐ�߼��߯%��_J����:]�F�@ P�\����r]�Dz��q�\�N� ���NA.O I �,�>�P� b�t�:��ߢ�d�v��� ��/����(�>�L� ~�<No�������� �� $f&�~8���>�P� b�t���r}� I/�����/�/ 1/C/�/g/�/�/�/�/ �/?���?��?�?�?��Ȝ�0�#F�˷ �??N;c�?�O`�� T�d�0�u�BP��qo� �p3e3�$:�O'7Lp$D �1˺�D6^�ud��H�4�����\�_�X>����4�ZOO0OBO TOfOxOQo�O�O�O�O  _�o__,_>_P_b_ ;�_�_q�_�_�_�_ o�(o:o�^opo�o �o�o�ov��o�o  $
�HZ3�~�|�? �?k�}�����2��؟��������7�2 2�[�m��������ǯ ٯ�������I�i� �ɔʉ������؂� ����ٷ�ɿ����h���-Ǚ�����Y�
E��>M1t��k8`��>L����x�{��<#�
�qx�p�� �]���T����D�H���8�Y���@��L2d�� �t�����
}�7��*�By��ŝ��$�6� �Z�l��	�>]��������It$ Z��$)�>���
��
�A��
���,������9�+���x�.������8�$敕��(4$ܠ�X�j��;��.��>��yH��8�5����O8M�Y��@�=�� 8��!G�	>�W B{f���������$CCS�CH_GRP1B 2���4�&� �\(��/+�  �a0,�Ԭ�	Б yP�~1؝���P4��T��V0��D5?333@řA�|����D/  Ce��G�P ?fff@�>)х�D5�)}!� �V�"d=l�@�['h9 D�'?9?Z?,���/A?x�?��� F@ �50�!A%`�� Dzo �4��/�?�?[:ˑ���� ܩ/�/�/�/�/�O ?O�O�O]?o?�oO �O�O�O�O�O�O�_�_ �_#_5_G_Y_k_}_�_��_�_�o�o"o�_�l� 5o�?�?�?�?�?O O���o�0B Tfx�D���R� �6���,�>���6E�e�LO&�8�J�TH� ob�n���H������ �����eQ"���bb� 0�-���H���=а��� ��Z�������b�H5� ����J�Y�<�v�x	��'�>���Y� '���������џ��� ο�+�=�O�}�υ� ������ͯ߯���� ��9�K�]�o���Kߥ� ����ۿ����?�5� ��Y�k�}Ϗϡχ��� �ϰ���M�$�V������"�2w<U�g�y�����{��2������ �� 2DVhz �4x>�����)*� ]ma)a)U�joPgz�|9@4Fsj����@�(,������>ʁ����b�bn��>LG .!n����O<#�
���p����e>�����������%�"��5%@ �a6$ɂ�/��T�ebR�@6]j�/�҅ߧ�B�� %?�?�?�?�?�?�?�ۆ >�!Z$�{<O^It$ UO$��K>�["
5O�GA��O/O�OSOeF�+�{���E.���U޵$敕U(4�$�U�O�K;��=.IU>��HUU��5��eU8M�	YqU�=. �U�^��_�K	�O�_�_�_�W 1_#o8oJo\ono�o�k��$CCSCH_�GRP1C 2�����a?&� \��j�>��  a�ހ �"~$)2� u�e�
�a �(,>P�RgU~���Ӏc#��?3�33�r�51D�/  C��G�P_ ?fff�>�! ����qߏ��o|� ����w��?���� ׏�ՑD�����W�F@ J�V��u�"W�Dz�pk�V�H��p؊H�(�� �&� 8�J�\�n�4�����^� p�ڏ������"� 8�F�x�6�H�i����� į֯�����`�� ϟ�x�2̸����� 8�J�\�n�������" wω�C߭Ͽ������� ���+�=���a߳߅� �ߩ߻�ﳕ��ɟ������јȖ����� @9�g{�9�5/���� Z��rN0^���%��J4 �!i6� --9���!� F ����j��0�%^v�����O�/���>�����
�� *�<�N�`�r�K���� �������&8 J\5/��k/�� ���/"4?X j|���p?�� �//?B/T/-Ox/��,����eOwO�O�E2@��O�O�O_]�?1R2,_U_g_y_�_�_ �_�_�_�_�_����n CAc4�y�z�<ڽ�y�y �2�ͷ�?���o�o�o�ovb4�@'w�o�i(�ASw?S�!>G�n�	Me�Z��3{u>L��p�q�/ub
I<#�	
�!r2p{rWŻ?vNb���!>5B1�u2�S0�u@���tF� ^�	O�$��/��ںw�12?$KBs1�u������0��T�f�;�>�W��t�o���cItk$ ҟ$#V>��r	
���A�d���&�xП�3p+���r��.���~�2q$�{����(4$ܚ��R�d�;��.ƥ>���Hҥ2q5�=��8M�Y�:m�=�p
�2r�1�A�	 8�Q�<�u�`��������ǿٿ�����$C�CSCH_GRP�1D 2����.�&� �\"N��%I  �2[�&��t�� ���s�Jjx�+��ϩ�@����.�����Nb�P�y�s>�?333:u��;t~i��D/  �C_0G�P ?fff:q>#�d>�� wі/HP���^�fm: U�b�>�!�3�T�&5o���;��:��F@� ����;�Z���Dz i��������U��A�O�I ܣߵ����� �߱�������W�i� �/i�{����������� ���/ASe w��������/��/������ �����/�r�/�/ */</N/`/r/�/>?�/ �/L?�/0???&?8? �?0�_OF� O2ODON��\@h3��B��? �N�|cO _�K�ˀ �\@*�'RǄB��7� �e���:T_�7�p�D\A�B�/T�^���DXSD�6�p�lo!h>���SD!j�O�O�O�O�O �O�O�o_%_7_I_w_ _�_�_�_�_�_� �_o�3oEoWoio�o E��o�o���o�o�o 9/�Sew�� �������G�OPO�����2q�O�a�Hs�����u���2�� ү�����,�>�P� b�t�{�r����� � �W[�[�O�dJ t�v�.�@�m�dω�߄����"�&��Ǽ�|�>�1�φ���h���>LA�(�h�<򲇙<#�
�p�ϗ��8���˲��|�����կ�Ѐ/�@|0��2�߆�N� _L��W�߮����B����z���������>��T��xu�6��It$ O�-$��>�U�
/���Aā�)���M�_����+�����.��y�����$敕�(4$�����;���.C>��H�O��5��_8'M�Yk��=(Ї��X����	���� ��+2DVh�z��$CCSC�H_GRP1E �2�����&� \���d?��   [��0��x�#��%� Ǻ���/&/8/J/�(a/O.˲��0]ӻ5?333��"�����/�D/  C܀G�P ?fff��>�����5�)�!��� �v2�=㽷��'�9�� �?�?�?����>?�?O<�Q0F@ DEP1�%��Q0Dz� eDP?�BOO�:B�"�� � ?2?D?V?h?._�? �OX_j_�?�?��O�O 
__2_@_r_0oBoco �_�_�_�_�_�_oo@Zo�oro,|��o O�2ODOVOhOzO�O ��q�=���� �����%�7�ɏ[� ������������Eܟ`�O�������HȐo ِ�:�u�3�/��� ��}�Tu�"H�Xrِ�� ��D��c��'�'�� ѯ�@��ّ���*��X&��Д���߀�<����>���Д��  ��$�6�H�Z�l�E� ������Ư�������  �2�D�V�/�z���e� ��¿Կ�����.� �R�d�vψ϶Ϭ�j� ����������<�N� '�r��ܛ�͟_�q�����2�<������	��+2&Oas ��������4 �>=�]�)�*}��m �)�)���o�g���9� ���&\���!'�����M'9��>�A�h/�_rTr��u%�>L� �!��o�<'#�
��l�pu/"pQu��&H����@8�<�%,2M�%@�a �$@�X?����b�ߋ6 �jq?+����Bm�% �?�?O*OONO`O�� >Q1�$���O��It$ �O$>%��"
�O�GA��O�O _�O�F- +��=�lU.���xU,!�$敕�U(4$�ܔUL_^[;��.��U>��H�U,!5����U8M�Y�U4=� e,"��o;[	2_Ko6oooZg�_��o�o�o�o�o�o{��$CCSCH_G�RP1F 2����(q&� \���  ��U� 2 �$�2� �umuDrq%8 ����(b��~H��J��#8�?33�34%�r5$x�1D/�  CY�G�P /?fff4!>1y 8�y�q����J�X� `4/O�\�8O�-�N�� ���5�����΀F@ ��́5�T2΀Dzc��͏����O�8����� ܝ��� ��ӏ叫�	��կ� Q�c���c�u������� ��ﯭ�����)�;� M�_�q�����׿�ϗ��￩̸)ϋ�߯� ��ӟ���	�߈"��  ߺ�$�6�H�Z�l�~� 8�ߴ�F���*����  �2�|�*�Y�@��,�>�H���V�b�9 <w����/v����� E��0��V�$5!�4<1 �610��9��N��  ��V�<z)��%�v>�M�0_j?�>���M�}����� ���������1 Cq/y���� ��/�	�/-?Q c�??���?�� �/3/)/�?M/_/q/ �/�/{?�/�/�O�/A<@�J��O�O _U2k� I_[_m__�]oO�R2�_�_�_�_oo&o 8oJo\onou�l��n�A �4���<Q�U�U�IB ^�D�nOp�(:g^�v�4	P�w
y Q�w�Sv1>����Mp����bC�u>L;��"�b?�b�I<#�
	1�2p��r��2O�v�b��v1�5�1����0)�@v�*���Տ �OH4Y�F?�Q�2y?�KB�1��t���@����˟ݟ�;z�>΁�N�yo0�sIt$� I�$�V>�O�
)�{�At{�#���G��Y��p+����.�������q$�=��(4$��ɯ�۫;��.=�>���HI��q5���Y�8M�Ye��m=@"����rRA����	�� ȿ���׷%��,�>��P�b�tσ��$CC�SCH_GRP1�G 2������&� �\�N^�I  UB����r��z� ����j����� �2ߠDߥ�[�I��b���<W���?333�u
���t�i)�D/  C��0G�P ?fff�q>���d������ ?�H��p����m��� �鵟�����5�o8����	JK�F@ `>�J��тK�Dz�� _�J�<����<Q_Y ��,�>�P�b� (���Rd����	? ����,:l* <]������  T//�l&,���~/,�>�P�b� t����/�k/}/7?�/ �/�/�/�/�/�??1? �?U?�?y?�?�?�?�?����O���O�O�O��Ȋ�@�34���oO-^ )��c~Ow_N%��B�R" �@���R>���]���!u !�J�_G:�T�A��@�T$ny�RֻX�D����zl�o�h>��� �D�j�O__0_B_T_ f_?�_�_�_�_�_� �_oo,o>oPo)�to �o_��o�o�o�o�� (�L^p�� �d���� ���� 6�H�!�l����O�OY�k�}���2��Ưد�$����%�2 �I� [�m��������ǿٿ ������7�W��ق� w������ƒ��럀��Ϸ����� �V����ׇϙɝ�G�3��>;Ab���Y"N"ߓo�>L�П�ߏi��<#�
��f�p�o��K%���B����2�6���&�G���@���:BR���ń��Ï���k�%����B g��Ջ����$��H�Z����>K������ϼ����It$ ��$��>���
����A�����������'�+����f.����r&�$敕�(�4$܎FX;�{�.�>��H��&�5���8M�Y�.�=���&�ϑ5	,E0i T�������� +�$CCSCH�_GRP1H 2����"!&� \�|�?�  Ғ O@��Ԛ���%g%>� l!�/�/�/�/"�/��.B��D@��2E?333.Շ"/�rɦ��D/  CS�GÿP ?fff.�> �s�2Es9k1�� �D/ �2RMZ�.�I7VI2�O 'OHO�ϵ?/O�O���0F@ �E�1/5N��0Dz]0�D�?�O��OIJ������ � �?�?�?�?�?�_O_ �_�_KO]O��]_o_�_ �_�_�_�_�o�o�oo #o5oGoYoko}o�o�o ��o�|�#�O ��O�O�O�O�O_	� �������0�B�T� f�x�2�����@�ҏ$� ����,�v�$US�:_0�&�8�BX�P� \���6'쟪���p��� ���u?2���rP��� ��6���+��Ş鏚H� ���Џ�P�6*#������&8�G�*d���	��>���G��w� ��������ѯ㯼�� �+�=�k��s����� ����Ϳ������'� 9�K�]��9�ϥ�~� ��������-�#���G� Y�k�}ߏ�u���ߞ� ��;��D��������2eLCUgy�i��2�����  2DVhoDfN ������)�*��K}O9 O9C�X>wh�jI"/4/a/X/}&�� �'/P)�'�p�>����/z��r�r\��%>�L501\��{�<#�
���p�/�"�u8,��&���p�� ��5�2��#5@pq$4 ���?z�B�Sr@�FKz�?��s��B��5O nO�O�O�O�O�O��t0�>�1H4s/i/*_#I�t$ C_$�>�I2
#_uWA $u__�_A_SV� +��̞�U.����U�!$�敕�U(4$�xe�_�[;��.7e�>��HCe�!5{��Se8M�Y_e�=0{e�"L�o�[	�_�o�o�o�go�&8J\n}{�$�CCSCH_GR�P1I 2�����q&�� \��X���  O�̐�2l4 Bt0�u�u��q�8���,�>��bU�C������Q3��?333�%��$�#AD/ � C��G�P ?fff�!>�1��� ����}��j�ϝ� �/Ƈә�O����ş���2�����E�F�@ 8�D����2E�DzڀY�D�6��ƚ6	 ��&�8� J�\�"�����L�^�ȟ ڟ�گ����&�4� f�$�6�Wώ�����Ŀ ֿ����N���ߍ�f� ܸ���x�&�8� J�\�n������"e�w� 1�߭߿������߯� �+��O��s��� ���������������Ȅ�����.I�w i�'#?�x�qHռ� <@L���5�8D�1WF �0%I���40 ��z�s5L������_�?t��>��������* <N`9/���� ��/�&8J #?n�Y?���� ��?/"/�?F/X/j/ |/�/�/^O�/�/�/�/ ?�?0?B?_f?�<�� ��S_e_w_�U2��_��_�_�_m�Ob2 oCoUogoyo�o�o�o �o�o�o��~1QQD |�|�qL��̉̉�B�� ���O癟����vPD�P���y�QA�
-c�1>5�\��MS�8H��Ci�>L����x�?cr�I<#�
�1`Bpi��EթO�<r���1,E0A�� �A@��@����4�L��O �4�½?���e�B�?[BaA������� �B�T�K�>E�ń�����~sIt$ Z��$f>�Ƃ
���A}t򯚯���Ц�!�+���`�.����l� �$敕|�(4$܈�@�R��;��.��>��yH�� �5��еO8M�Yܵ(}=�� �� ��A	�/�	&�?� *�c�Nǜ��ϣϵ�����������$CCS�CH_GRP1J 2�����&� �\^��Y  �BI��鄔��y� a�8zf���ߗߩ߻�P�����<r�>�΃,�?333(���)�|ly��D/  CM@�G�P ?fff(�>�mt,�m�e�? �H>���L�T}(�C�P� ,��!�B�E�o��)�x���J��F@ ��0��)�H���DzW��������C��Q�_�Y ܑ������� ����E�W��?W i{������ �/ASew���y/�/
/��,� /��/���������� ��?|��/�/�??*? <?N?`?r?,O�?�?:O �?O�?OO&OpO�M_4_ _2_<� /JPVC��0��O�^�� js�O�_�%9⹐�"JP �b��0�Ԗ%��u�� �JBo�G���TJQ0�d �n����2hAT$�^�x�lx>���AT zq_�_�_�_�_�_�_ �oo%o7oeo�mo o�o�o�o�o���o�o ֏!3EWy3�� �x�����'�� ۟A�S�e�w���o��� �����5�_>_Я���
�2_�=�O�a�s���c���2����ҿ �����,�>�P�b� i�`��ή�Δ����� E-I�I�=�R/8'b�d�@�.�[�R�w�͔��@�������ת�j�>�A��t��"�"V���>L/��V���u�O<#�
��ݒp������%&��ֹ����j������⾐�@ j!�B��t�<�M":�@��E*�m���Bޑ ��h�����~�������n�>��B�m�c�$^��It$ =$��K>�C�
oA���o�;M��+�{���.����ޝ�$敕�(4�$���;��=.1>��H=���5��M8M�	YY��=�u��F���	����� / /2/D/V/h/w+��$CCSCH_�GRP1K 2�����!?&� \��RO>��  I��@ ��f��n��%�%���! ��??&?8?�O?=>ʹ���@K�E?3�33���"�����D�/  CʐG�P_ ?fff��>�� �ĩE�9�1�w��/dB �M�ͥ��7�I���O�O �O��y�,O�O _��?@F@ 2U>A�5��?@Dz�0ST>O0__p�J0��� �O  O2ODOVOozO�_Fo Xo�O�O���_�_�_
o  o.o`o0Q�o�o �o�o�o�o�oH���`����Or�  _2_D_V_h_z_���� _�q�+�������ˏݏ ��%���I���m� �����ퟛUʯ�_�������X�~Ǡӓ (��'c�!����r�k� B��26�F�Ǡ�咲2� ��Q��������	� .��ǡ�*���m�F6�������ǹό�>�������� � �$�6�H�Z�3�~��� ����⿄����� � 2�D��h�z�S�ϰ� �����ϰ�
����@� R�d�vߤߚ�X����� �������*�<�`쉯��M_q�2@�L������2=Oas� ������D�N . +K�v9v:k��}�9�9 ����w���I�/�/�/�/�&J�z 7{/�)(�;7'��>/�V?���M�B���c5>L�0�1��]"��<#�	
z�Z�pc?2?���66"����&�*��5B;�5@�q�4.� FO�����r��yF�z_O���B[�5O�O�__�O<_N_��0>�?A�4�/�/�_x#Itk$ �_$>��2	
�_�WAw$�_�_ox�_�V0+���Ze�.���fe1$�{��ve(4$܂e�:oLk;��.�e>���H�e15�=��e8M�Y�e"-�=�0�e2��)k	  o9$]Hw�o�� ����$[