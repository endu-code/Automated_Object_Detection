��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1d�DDd!OE4LA!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTc@�D5�F6�F7�F8�F9�G0�G�GJA��E�GbA�E�G1�G1��G �F�G2�B!S�BN_CF>"
 }8F CNV_J� �; �"�!_CMNT��$FLAGS<]�CHEC�8 �� ELLSETU�P � $H�O30IO�0� %��SMACRO�RR'EPR�X� D+�0��R{�T UTO�BACKU��0 �)DEV�IC�CTI*0��� �0�#�`B�S$�INTERVAL�O#ISP_UNI�O`_DO>f7ui�FR_F�0AIN��1���1c�C_�WAkda�jOFFu_O0N�DEL�h�L� ?aA�a1b?19a�`C?��P�1bE��#sATB�d���MO� �cE D [M�c���^qREV�BIL�rw!XI� QrR o � OD�P~�q$NO^PAM�Wp�t�r/"��w� �u�q�r�0D~`S p E �RD_E�pCq$�FSSBn&$CH�KBD_SE^eA�G G�"$SL�OT_��2=�� V��d�%��3 a_�EDIm   �� �"��PS<�`(4%$EP�1�1O$OP�0�2�an�p_OK�UST1P_C� ��d��U ^�PLACI4!�Q��4�( raCOMM� ,0$D����0��`��EOWBn�IGA�LLOW� (�K�"(2�0VAR�a��@�2ao�L�0OUy� ,Kvay�r�PS�`�0M_O]�����CCFS'_UT~p0 "�1 �3�#�ؗ`X"�}R�0  4F IMC	M�`O#S�`��up�i �_�p�BAw��a���M/ �h�pIMPEE_F�N��N���@O���r�D_�~�n�Dry�F� dCC_��r0  T� '��'�DI�n0"��pu�P�$I�������F�t XF� GRP0��M=q�NFLI�7��0U�IRE��$g"� S�WITCH5�AX�_N�PSs"CF_�LIM� �; �0EED��!���qP�t�`PJ_dVЦMODEh�.Z`��PӺ�ELBOF � ������p� ���3���� FB/���0�>�G� �>� WARNM�`/���qP��n�NST�� COR-0bF�LTRh�TRAT�PT1�� $AC�C1a��N ��r$�ORI�o"V�RT��P_S� CHG*�0I��rT2��1
�I��T�I1��>� x i#�Q\��HDRBJ; TCQ�2L�3L�4L�5L�6L�7L� N��9s!��O`S <F +�=�O��#92^��LLECy�"MULTI�b�"N���1�!���0T�� �STY�"�R`�=l�)2`����*�`T  |� �&$��۱m��P�̱�UT�O���E��EXT�����ÁB���"2Q� (䈴![0�������<�b+�� "D"���ŽQ��<煰kc!(�9�#���1���ÂM�ԽP��" q'�3�$ L� �E���P<��`A�$�JOBn�T���l�TwRIG3�% dK� ������<���\��+��Y�p�_M��&� t�pFLܐBN9G AgTBA� �� �M��
�!��p� �q��0�P[`��O�'[���0tna*4���"J��_R���ECDJ��IdJk�D�%C�`�Z���0���P_�P��@ ( @F RO.��&�t�sIT�c�NOM�0
����S�`TE)w@���Z�P�d���RA�0��2b"�����
$T����MKD3�T��`U31����p(5!HGb�T%1�*E�7�c�KA�b�WAb�cA4#YNT|���PDBGD��2 *(��PUt@0X��W���AX��a���eTAI^cBUF���0!+ � �7n�PIW�**5 P�7M�8M�9
0��6F�7SIMQS�@>KEE�3PATn�^�a" 2`#�"��L64FIX!,C ���!d��D�2B�us=CCI�:FPCH�P:BAD�aHCE hAOGhA]HW�_�0>�0_h@�f�Ak���F��q\'M`#�"�DE3�- l�p3G��@FSOES]FgHBSU��IBS9WC��. `{ ��MARG쀜���FACLp�SLEWxQe�ӿl��MC�/�>\pSM_JBM��Ԁ�QYC	g�ew3�w0 ā�CHN-�;MP�$G� Jg��_� #��1_FP$�!TCuf!õ#@�����d�#a��V&�0�r�a;�fJR���r�SEGFR�PIO�� STRT��N��cPV5���!41�r��
r>İ�b�B��O�2` + �[���,qE`&�,q`�y�Ԣ}t��yaSI!Z%���t�vT�s� ��z�y,qRSINF }Oбc���k��`���`�`L�ĸ T`7�C3RCf�ԣCC/�9���`a�uah�ub'�MI�N��uaDs�#�G�D
�YC��C�����e�0q0��� �EV�q�UF�_�eF��N3��s�ah��Xa+p,�5!�#1�!VSCIA?� A��s1�"!3 ��`F/k��_ �U��g��]��C�� a��s�"R�4� �����N����5a�R��HANC��$L�G��P�f1$+@NYDP�t�AR5@N^�`�a�q���c��ME�108���}0��RAө�CAZ 𨵰�%O��FCTK��s`"��S�PFADIJ�O J�ʠ�ʠ���<����Ր��GI�p�B�MP�d�p�Dba��AcES�@	�K�W_���BAS�� �G�5 � M�I�T�C�SX[@@�!62�	-$X���T9�{s�C��N�`�a~P_H�EIGHs1;�WI�D�0�aVT ACϰ�1A�Pl�<����EXPg���|��C}U�0MMENU���7�TIT,AE�%)�a2��a��g8 P� a�ED�E� ��PDT��R�EM.��AUTH?_KEY  ����R�� �b�O	���}1ERRLH� �9c \� �q-�OR�D�B�_ID�@l �PU�N_O��Y�$SCYS0��4g�-�I��E�EV�#q'�P�XWO�� �: �$SK7!f2 VR�(�Td�TRL��; �'AC�`��Ġ7IND9DJ.D���_��f1��f���P5L�A�RWAj��"�SD�A��!+r|>��UMMY9d�F�C10d�&���J�<��v}1PR� 
3��POS��J�= l�$V$�q
�PL~�>���SܠK�)?����CJ�@�����ENE�@T��A����S_�RECOR���BH 5 O��@=$LA�>$ ~�r2�R��`�q�b`�3_Du��0RO�@�aT[�Q��b������x! }У�PAUS��>�dETURN���MRU�  CR�p�EWM�b�AGNsAL:s2$LA��!?$PX�g@$P�y A ��Ax�C0 #ܠDO��`X�k�W�v�q�GO�_AWAY��MO��ae���]�CSS�_CCSCB C� �'N��CERI@��гJ`u�QA0�}��@�GAG� R�0�`��{`��{`OF�q�5���#MA��X���&шLL�D� �$���sU�D�)E%!`���OVR310W�,�OR|�'�?$ESC_$`�eDSBIOQ��l q��B�VIB&� �c,�����f�=p�SSW���f!VL���PL���ARMLO
��`����df7%SC �bALspH�MPCh �Ch P�#h �#h 5�UU� ��C�'�C�'�#�$'�d�#C\4�$�pH���Ou��!Y��!�SB ���`k$4�C�P3�Wұ46$VOL�T37$$`�*��^1��$`O1*�$,o��0RQY��2b4~�0DH_THE�����0SЯ4�7ALPAH�4�`���7�@ �0T�qb7�rR�5�8 8� ×���"��JFn�MӁVHBPFUAFLQ"D�s�`�THR��i2dBP�����G(��PVP������������1�J2`�B�E�C�E�CPSu� Y@��Fb3���H�(V �H:U�G�
X0��FkQw�[�Na�'B���C �INHBcFILT���$��W�2�T 1�[ ��$����H YАAF�sDO ��Y�Rp� fg�Q� +�c5h�Q�iSh�Q�PL���Wqi�QTMOU�#c�i�Q\��X@�gmb��vi�h�bAi�fI�aHIG��caB	xO��ܰ��W�"v�AN-u!��	#AVj�H!Pa8$P�(ד#p�R_:�A�a���B�N0�X�M�CN���f1[1�qVAE�p��Z2;&f�I�Q�O�u�rx�wGldDEN{G|d��aF>�!�9��aM:�U�FW	A�:�Ml���X�Lu���$!����!l�ZO ����0%O�lF�s�1&3�DI�W�@���Q���_��!CUgRVA԰0rCR41ͰZ�C<�r�H�v����<�`��<�(�f�CH �QR3�S���t���Xp�VS_�`�ד��F��ژ����?NSTCY_ OE L����1�tP�1��U��24�2B��NI O7������DwEVI|� F���$5�RBTxS�PIB�P���BY�X����T��HN�DG��G H tn���L��Q��C���5��Lo0 aH��閻�FBP�{tFE{�5�t��T���I�DO���uPMCS�v>�f>�t�>"HOTSW�`s��ІELE��J T���e�2��25�� O� ��HA7�E��3�44�0趘�A�K �� MDL� 2J~PE��	A��s��tːÈ�s�JÆG!�rD"�ó�����\�T�O��W�	��/��S�LAV�L  �0INPڐ���`%��_CFd�Mw� $��ENU��OG��b�ϑ]զP�0�`ҕ�]�IDMaA�Sa��\�WR�#���"]�VE�$a�SKI�STs��sk$��	2u���J�������p	��Q���_SVh�EXCLUMqJ2M!'ONL��D�Y��|r�PE ղI_V��APPLYZP��HcID-@Y�r�_M�2=��VRFY�0��xr�1�cIOC_f�D�� 1������O���u�LS���R$D_UMMY3�!��z�S� L_TP/B�v�"���AӞ�ّ �N ���RT_\u�� N�G&r�[�O D��P_B�A�`�3x�!IF ��_5���H���N���� �� P y$�KwARGI���� q�2O[�_S;GNZ�Q �~P/�/PIGNs�l�$��^ sQANNUN�@�T<�U/�ߴ�LAzp]	Z�Xd~N�EFwPI�@_ R @�F?�IT�	$TOT�A%��d���!ڙM�NIY�S�+���E�A[�
D7AYS\�ADx�@���	� �EFF/_AXI?�TI��0�zCOJAM�ADJ_RTRQ��Up��<P�1D D�r5̀Ll�T�0�? ]P�"p�� �A8tpd��V 0w��G��������SK��SU� ��CTR�L_CA�� W>�TRANS�6PIDLE_PW����!��A�V��V_��l�V �DI�AGS���X� �/$2�_SE�#TAC���t!�!0z*L@��RR��vPA��4�p ; SW�!�! �  ��ol�U��o3OH��PP� ��sIR�r��BRK'#��"A_Ak���x 2 x�9ϐZs2��%l��W�0t*�x%RQD�W�%MSx�t5AX��'�"��LIFEC�AL���10��N �1{"�5Z�3{"dp5�xZU`}�MOTN°9Y$@FLA�cZgOVC@p�5HE	>��SUPPOQ�ݑ�Aq� Lj (C�1_�X6�IEYRJZRJW�RJ�0TH�!UC��6�X�Z_AR�p��Y2��HCOQ��Sf6A�N��w$w��IC�TE�Y `��CACHE�C9��M�PLAN��UFFIQ@�Ф0<Ѩ1	��6
��M�SW�EZ 8�K�EYIM�p��TM~�SwQq�wQ#���}�OCVIE� ��[ A�BGL���/�}�?����D�?��D\p�ذST��!�R� �T� �T�� �T	��PEMAI�f�ҁ��_FAKUL�]�Rц�1��U�� �TRE��^< $dRc�uS�% IT�ӇBUFW}�W��N�_� SUB~d��C�|��Sb�q�bSAV �e�bu �B��� �gX��^P�d�u+p�$�_p~`�e�p%yOTT����sP��M��OtT�FLwAX � ��X~`�9#�c_G�3
�YSN_1�_�D��T1 �2M���T�F��H@ g�?`� 0p���Gb-sC_R�AIK ���r�t�RoQ�u�7h�qDSPq��rP��A�IM�c6�\��Ä�s2�U�@�A�sMF*`IP���s�!DҐ�6�TH�@n�)�OT��!6�HSDI3�AGBSC���@ Vyİ�� �_D�CONVI�G���@$3�~`F�!�pd��p�sqSCZ"���sM3ERk��qFB��k��pET���aeRFMU:@DUr`����x�CD,���@p;cH%R�A!��bp�ՔXՔ+PSԕCN�e�C��p��ғSp�cH *�LX�:cd�Rqa�|  ����W��U��U���U�	�U�OQU�7R�8BR�9R��0T�^�1k�U1x�1��1��1��U1��1��1ƪ2Ԫ�2^�k�2x�2��2���2��2��2��2*ƪ3Ԫ3^�3k�x��3���o���3��3���3ƪ4Ԣ�%�X9Tk!0�d <� 7h �p�6�pO��p����Na�FDRZ$eT^`V�Gr����䂴2�REM� Fj��BO�VM��A�TR�OV�DT�`-�MX<�IN��0,�W!'INDKЗ
w�׀�p$DG~q36���P�5�!D�6�RI�V���2�BGEAR��IO�%K�¾DN �p��J�82�PB@�CZ_MCM�@�1��r@U��1�f ,⑞�a? ���P\I�!?I�E��BQ����`m���g� j_0Pfqg RI9e�j�k!UP2_ 3h � �cTD�p�〪�! a���$��bB;AC�ri T�P�b��`�) OG��%p���p��IFI�!`�pm�>��	�PT�"���MR2��j ��Ɛ+"���� \��������$�B`x%J��_ԡ�ޭ_�İ�� M������DG�CLF�%DGDY&%LDa��5�6�ߨ�4@��Uk���� T�FS#p�Tl� P���e�qP�p�$EX_���1PM2��2� 3�5�s�G ���m ���֍�SW�eOe6DE�BUG���%GRt���pU�#BKU_��O1'� �@P�O�I5�5M�S��OOfswSM���E�bUP�0�0_?E n �0 ��TERM�o��XPO�ORI�+�p��&
�GSM_���b�q��   �TA�rڢE�UP�Rs� -�1�2n$|�' o$SEG,*�> ELTO��$wUSE�pNFIA�U"4�e1���#$p$UFR���0ؐO!��0����OT�'�TqAƀU�#NST��PAT��P�"PTHJ����E�P rF�V"ART�``%B`�a�bU!REL:�aS�HFT��V!�!�(_�SH+@M$���� ���@N8r����OV9Rq��rSHI%0���UN� �aAYLO����qIl����!�@��@ERV]��1� ?:�¦'�2��%��5��%�RCq��EAScYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba��
5aPo��0�p6OR��MY� `GR��t 2b5n� � ��UPaN�Uu Ԭ")���TOCO!S�1POP ��`�pC�����e��Oѥ`REP�R3��aO�P�b�"ePR�%WU.X1���e$PWR��IM�IU�2R_	S�$VI1S��#(AUD���D�v" v��$H|���P_ADDR��H�G�"�Q�Q�QБqR~pDp1�w H� SZ�a��e�ex��e��SE��r��H�S��MNvx ���%Ŕ��OL���p<P��-���ACROlP_!QND_C��ג�1�T �OROUPT��B_�VpQ�A1Q�v��c _��i���i��hx��i����i��v�ACk�I	OU��D�gfsu^d��y $|�P_�D��VB`bPRM�_�b�ATTPu_אHaz (���OBJEr��P��-$��LE�#�s`�{ � ��u�AKB_x�T~�S�@��DBGLV��K�RL�YHITCOmU�BGY LO a�TEM��e�>Ҙ+P'�,PSS|�P�J�QUERY_FLA�b�HW��\!ae|`u@�PU�b�PIO��"�]�ӂ/d�ԁ=dԁ�� �IO�LN��}����C�Xa$SLZ�$�INPUT_g��$IP#�P��'���S	Lvpa~��!�\�W��C-�B����pF_�ASv��$L  ��w �F1G�U�B0�m!���0HYp��ڑ����UOPs� `������[�ʔ[�і"�[PP�SIP��<�іI�2���P_M�EMB��i`� XƟ�IP�P�b{�_N�`����R��̬��bSP��p$F�OCUSBG�a4� �UJ�Ƃ �q  � o7JOG�'n�DIS[�J7�cVx�J8�7� Im!|�)�7_LAB�!��@�A��APHI�b�Q�]�D� J�7J\���� _KE}Yt� �KՀ�LMONa����$XR��ɀ��WATCH_��3���EL��}Sy~���s� �Ю!V�g� �CTR3򲓥��LG�D� �R��I�~
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�Gȴ I�F�%SO���q �Ɩ�@��v��ƴ��K�S�����w�k�N����E��\���'�"*�U�s5��@L>�4�7DAUZ�EA�pՀ�Dp�f�GH�B�q���BOO��� C���PIT���� REC��SCR�N����D_p�aMARGf�`��:����T�L���S�s��Wp�Ԣ�Iԭ�JGMO��MNCH�c��FNt��R�Kx�PRGv��UF��p0��FWDv��HL��STP���V��+���Є�RS"��H�@�몖Cr4�� ?B��� +�O�U�q��@*�a28����Gh�0PO��������M�8�Ģ��EX��TU%Iv�I��(�4� @�t�x�J0J�~�P��J0��N�a�#A�NA��O"�0VAI|A��dCLEAR�6?DCS_HI"��/c�O�O�SI��S��IGN _�vpq�uᛀT�d� 7DEV-�LLA Ѧ°BUW`���x0T<$U�EMH��Ł����0�A�R��x0�σ�a�@WOS1�2�3�p���� `� ����h�AN%-���-�ID%X�DP�2MRO��Ԭ�!�ST��Rq�Y�{b! �$E�&C+��p.&A&8���`� L��ȟ@%Pݘ��T\Q�UE�`��Ua��_ � ��@(��`�����# ?�MB_PN@ R`�r��R�w�TRIN8��P��BASS�a�	6IRQ6�aM�C(�� ��C�LDP�� ETRQ�LI��!D�O9=4FALʡh2�Aq3zD᱌q7��LDq5[4q5ORG�)�2�8P�R���4/c�4=b-4�t�� �rp[4*�L4q5SB�@TO0Qt�0*D2FRCLMC@D�?�?�RIAt,1ID`�D� Yd1��RQQprp�DSTB
`� �F�HAXD2���G��LEXCES?RR�EMhPa���B�D4�E�q`�`�F_A�J�C[�O�H:� K��� \���b2Tf$� ��LI�q�SREQUIRE�#�MO�\�a�XDEB�U��,1L� M䵔 �p���P�c�AA"$RN��
Q�q�/�&����-cDC��B�IN�a?�RSM�Gh� �N#B��N�iPST�9� � 4��L�OC�RI���EX�fANG��A,1�ODAQ䵗�@1$��9�ZMF���� �f��"��%u#ЖVgSUP�%QFX�@�IGGo�� � rq�"��1��#B��$���p%#by��rx���v<bPDATAK�p!E;����R��M��*�� t�`MD�qI���)�v� �t�A�wH8�`��tDIAE��sANSW��th��
�uD��)�bԣ(@$`�� PCU_�V06�ʠ�d�PLOr�$`��R���B���B�pp�����RRR2�E��  ��V�A�/A d$CALII�@��G~�2���!V��<$R�S�W0^D"��ABC~�hD_J2SE�Q\�@�q_J3M�
G�G1SP�,��@PG�Bn�3m�u�3p�@���JkC���2'AO)IyMk@{BCSKP^:�ܔ9�wܔJy�{BQ�ܜ�����`_A1Z.B��?�EL��YAOCMP�c|A)���RT�j���1�ﰈ��@1�������Z��SMG��pԕf� ER!��a[INҠACk�p�����b�n _���@����D�/R��3DIU��CDH�@
�:#a�q$V�Fc6�$x�$���`�@���b��̂�E��H �$BEL�P����!ACCEL����kA°IRCS_R�pG0�T!��$PS�@B2L����W3�ط9�< ٶPATH��.�Dγ.�3���p�A_ ��_�e�-B�`C����_MG�$DDx��ٰ��$FW�@��p����γ����DE���PPABN�R?OTSPEEup��O0��DEF>Q����$USE_���JPQPC��JYh����-A 6qYN�@�A�L�̐�L�MO�U�NG��|�OL�y�INCU��a���ĻB��ӑ�AENCS���q�B�����D�IN�I�����pzC��VE�����23�_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��PR9C����MOS� gT�MOpp�@-GPERoCH  M�OVӤ �����!3�yD!@e�]�6�<�� ʓA����LIʓdWɗ��:p83�.�I�TRKӥ�AY����?Q^���m��b��`p�CQ�� MOM�B?R�0u��D����y�0Â��DU�ҐZ�S_BCKLSH_C����o�n� ��TӀ���
c��CLALJ��A��/PKCHKO0�SNu�RTY� �q���M�1�q_
#c�_U�MCP�	C���SC�L���LMTj�_AL�0X����E� � �� ���m�0h���6��PC����!H� �P�ŞCN@�"sXT����CN_��1N^C�kCSF����V6����ϡj���nnCAT�SHs �����ָ1���֙����������PA���_	P���_P0� e���0O1u�$xJG� P�{#�OG���TORQU(�p�a�~���`�Ry������"_W�� ^�����4t�
5z�
5UI;I ;Iz�F�``�!��_8�1��VC��0�D�B�21�>	P�?�B�5JRK�<�2�6~i�DBL_SM�Q:&BMD`_DLt�&BGRV4
Dt�
Dz���1H_���31�8JCcOSEKr�EHLN�0 hK�5oDt�jI��jI<1�J�LZ1�5Zc@y��1cMYqA�HQBTHWM�YTHET09�N�K23z�/Rn�r@C�B4VCBn�CqPASfaYR<4gQt�gQ4V�SBt��R?UGTS���Cq��a��P#��<�Z�C$DUu ���R䂥э2�Vӑ��Q��r�f$NE�+pI�s@�|� �$R�#QA�'UPeYg7EBHBALP!HEE.b�.bS�E�c �E�c�E.b�F�c�j�F�R�VrhVghd��lV��jV�kV�kV�kV*�kV�kV�iHrh�f��r�m!�x�kH�kH��kH�kH�kH�iOJclOrhO��nO�jUO�kO�kO�kO�kO�kO�FF.bTQ����E��egSPBAL�ANCE��RLE6�PH_'USP衅F���F��FPFUL�C�3��3��E��1=�l�UTO_p �%�T1T2t���2N W�����ǡ��5�`(�擳�T�OU���>� INSEG��R��REV��R���DI�FH��1���F�1�;�OB��;C���2� �b�4LCHgWAR��;�ABW!~��$MECH]Q��@k�q��AXk�P���IgU�i�� 
p���!����ROB��CR��ͥ*�C���_s"T � �x $WEIGHh�9�$cc�� �Ih�.�IF ќ�LAGK�8SK��K�7BIL?�OD��U�&�STŰ�P�; �����������
�Ы�L��  2��`�"�DEBU.�L�&�n��PMMY9���NA#δ9�$D&���$��� Qw �DO_�A��� <	���~�H�L�BX�P�N�Ӣ+�_7�L�t�OH  ��� %��T����ѼT�����TgICK/�C�T1��%������N��c����R L�S���S��ž��PROMPh�E~� $IR� �X�~ ���!�MAI��0��j���_9�����t�l�R�0CO�D��FU`�+�ID�_" =�����G_�SUFF<0 h3�O����DO�� ِ��R��Ǔن�S���P�!{������	�H)��_FI��9��O�RDX� ����3�6��X�����GqR9�S��ZDTD���v�ŧ4 =*�L_NA4���|K��DEF_I[� K���g��_���i���0��š���IS`i  �萚����e��"��4�0i�Dg����D� O��LOCKEA!uӛϭ�0����{�u�UMz�K� {ԓ�{ԡ�{����}� ��v�Ա��g����� ��^���K�Փ����!w�N�P'���^����,`�W\�[R��7�TEFĨ ��OULOMB�_u�0�VIS�PITY�A�!O>Y�A_FRId��F(�SI���R��H����3���W�!W��0��0_,�EAS%��!�& �"���4p�G;穯 h ��7ƵC?OEFF_Om��H�m�/�G!%�S.��߲CA5����u�G�R` � � �$R� �X]�TME�$R�s�Z�/,)ËER�T;�:䗰��  ]�LL��S��_SV�($�~����@���� �"SETU��MEA��Z�x0�u���>��� � � �� ȰID�"���!�*��&P���*�F�'����)3��#�A��"�5;`*�ЧREC���!7�S�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I���0�MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X17ࡐMO�R�� H	�CU �A3�z�1Q�
��3���$��FV���2SbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų7�=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	����y��t�#�}1� @�@;���O&E�RI#A��
N��@X�s�f�tQ��PL}1�,RTv�m�ATU}SRBTRC_T(qR��B �����$ �pƱ��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���U1P(4����PX��؆��q��3�w� �P�G�5� $SUB������t�JMPWAITO�,�s��LOyCFt�!D=�CVF	ь�y����R`�0��CC_C�TR�Q�	�IGN�R_PLt�DBTeBm�P��z�BW)�d���0U@���IG�az��Iy�TNLN��"Z�R]aK� N��B�0�PE�s���r��f�wSPD}1� L	��A�`gఠ�S��UN��{���]�R!�BD�LY�2���P��H�_PK�E��2RETRIEt��2�b�v��FI�B� ��м�8� 2��0D�BGLV�LOGgSIZ$C�KTؑ�Uy#u�D7�_�_T,1@�EM�@C\1Aě���R��D�FCHgECKK�R�P�0ʳ���@&�(bLE,c�" PA9�T���PJ�C߰PN�����ARh�0���Ӯ�P�O�BORMATTnaF�f1h���2�S��UXy`	�tQP�LB��4�  ^rEITCH��7��9PL)�AL_ �� $��XPB�q� C,2D�!��+2��J3D��� T�pPDCKyp��oC>� _ALPH����BEWQo���� ���I�wp � �~b@PAYLOA�Öm�_1t�2t���J3AR��؀դ֏�^laTIA4��5��6,2MOMCP������������0BϐAD���������PUBk`R��;���;��Ғ��z4�` I$PI\Ds�oӓ1yՕ�w�T2�w�Z��I��I��I���p����n���y�e`�9S)bT�S/PEED� G��(� Е��/���Е�`/��e�>��M��ЕSAMP�6V��/���Е#MO�@ 2@�A�� QP���C��n������� ����LRf`kb�ІE9h�EIN09��7 S.В9
yPy�/GAMM%S���D$GET)bP�ciD]��2
�IB�:q�I�G$HI(0;�A��LREXPA8)LWVM�8z)��g���C�5�CHKKp]�0�I_��h`eT��n� q��eT,����� �$�� �1�iPI� RCH�_D�313\��30L�E�1�1\�o(Y�7 ¾t�MSWFL �M.��SCRc�7�@�&���%n�f�SV���PB``�'�!�B�sS_SAV&0ct5B3NO]�C\�C2^� 0�mߗ�uٍa��u� ��u:e;��1���8��D�P��������� )��b9��e�GE��3��V���Ml�� 7� �YL��Q
NQSRlbfqXG �P�RR#dCQp� $�S:AW70�B�B[�ȤCgR:AMxP�KCL �H���W�r�(1n�g�9M�!o�� �F�P@}t$WP�u�P r ��P5�R<�RC�R ��%�6�`��� ��qsJr X��OD�qZ�U�g�ڐ>D� ��OM#w�J?\?n?�?��?��9�b"�L]�_��� |��X0�� bf��qf��q`�ڏgzf"��Eڐ��Bf�"�����FdPB���PM�QU�� �� 8L�QCOU�!5�QTHI�HO�QBpHYSY�ES���qUE�`�"�O.���  �P�@�\�UN���Cf�O�� P��Vu�x�!����OGRAƁ�cB2�O�tVuITxe �q:pINFO������{�qcB�e�O�I�r� (�@SLEQS��q��p�vgqyS���� 4L��ENABDRZ�PTIONt�����Q����)�GCF��G�c$J�q^r�� �R���U�g��rS�_ED����� ��F��PK��E�'NU߇وAUT<$1܅COPY���(��n�00MN��^�PRUT8R ��Nx�OU��$G�[rf�e�RGAD5J���*�X_:@բC$�����P��W���P��} ��)�}�E�X�YCDR|�N�S.��F@r�LGO��#�NYQ_FREQR�W� �#�h�TsLAe#����ӄ ��CRE� s�I�F��sNA��%�a�_Ge#STAT�UI`e#MAIL �����q t��������ELEM�� ��/0<�FEASI ?�B��n�ڢ�vA�]� � I�p��Y!0q]�t#A�ABM����E�p<�VΡY�BA!SR�Z��S�UZ���0$q���RMS_TR;�qb �� �SY�	�ǡ��$���>C��Q`	� 2� _�TM���� ��̲�@ �A��)ǅ�Ni$DOU�s]$Nj����PR+@3���rG�RID�qM�BAR�S �TY@��OTIO�p��� Hp_}��!����d�O�P/��� � �p�`PO�R�s��}���SRV���)����DI&0T������ #�	�#�4�!�5!�6!�7!�8��e�F�2��Ep$VALUt��%���=b��/��� ;�1�q�����(_�#AN�#�ғ�Rɀ(�>��TOTAL��S��PW�Il��R�EGEN�1�cX���ks(��a���`TR��R��_S� ��1����V�����⹂Z�E���p�q��Vr���V_H��DA�S����GS_Y,1�R4�S� {AR�P2� ^�IG_SE	s����2å_Zp��C_�ƂѿENHANC�a_� T ;�������INT�.��@yFPsİ_OVRsP�`p�`��Lv��o���7�}��Z�@�SL)G�AA�~�25��	��D��S�BĤD�E�U�����TE|�P���� !Y���
�J��$2�IL�_MC�x r#_��`T�Q�`��q���'�BV�C�P_� 0�mM�	V1�
V1�U2�2�3�3�4�4�
�!���� �� m�A�2IN~V�IBP���1�2��2�3�3�4�4�A@-�C2����p� MC_F,p+0�0L	11d���M50Id�%"Eã S`�R/�@K�EEP_HNADED!!`$^�j)C�Q����$��"	��#O �a_$A�!�0�#i��#REM�"�$��¨�%�!�(U}�e�$HPWD  `#_SBMSK|)G�q�U2:�P	�COLLAB� �!K5�B��� ��g��pIT�I1{9p#>D� ,��@FLAP��$SSYN �<M�`C6����UP_DLYzAA�ErDELA�0�ᐢY�`AD�Q}	��QSKIP=E�� ���XpOfPN1Tv�A�0P_Xp�r G�p�RU@,G��:I+� :IB1:IG�9JT�9JaР9Jn�9J{�9J9<��{RA=s� X����4�%1�QB� NFGLIC�s�@J�U�<H�LwNO_H�0�"�?��RITg��@_�PA�pG�Q� )��^�U��W��LV|�d�NGRLT�0 _q��O�  " ��OS���T_JvA V	�AP�PR_WEIGH��sJ4CH?pvTOqR��vT��LOO�Ј]�+�tVJ�е�ғA0�Q�U�S�XOB'�'�M��J2P���7�X�T�<a43DP=`�Ԡ\"<a�q\!��RD�C��L� �рR"��R�`� �RV��j8r�b�RGE��*��cN�FLG�a�Z��ΒSPC�s�UM�_<`^2TH2N�H��P.a 1� gP�p�11��� lQ �!#� <�p3AT� g�S�&�Vr �p�tMq�Lr����HOMEwr�t2'r�-?Qcu�
�w3'r����(���w4'r�'�9��K�]�o����w5'r뀤���ȏڏ����w6'r�!�3�E�W�i�{�
�w7'r힟��ԟ(����w8'r��-� ?�Q�c�u��uS$0�q�  �� sF�`�`�1�"`P����a�`/���-�IO[�M�I֠��)aR�pW=E�� ��0rZa*��� �5ވ�$DSB GN�AL���0Cpm�Sw2323�� �~`r��� / ICEQP���PEp��5PIT�����OPBx0��F7LOW�@TRvP�X�!U���CU�M���UXT�A��w�ER�FAC�� U���ȳCH��� t�Q  _��>�Q$L����OM��A�`�T�P#UPD7 Ad�ct�T��UEX@8�ȟ�U EFA: X"΁1RSPT����)�T ��PPA�0o�l���`EXP�IOS���)ԭ�_���%Ќ�C�WR�A��ѩD�ag֕`ԦFRIE3NDsaC2UF7P��ޤ�TOOL��MY�H C2LENGT_H_VTE��I�<�Ӆ$SE����?UFINV_����RGI�{QITI5B��Xv��-�G2-�G17�w�S�G�X��_��UQQD�=#���AS��d~C��`��q�� �$$�C/�S�`������S0f�����VERsSI� ��f��5��I��������AAVM_Y�2� � �0  �5���C�O�@�r� r�	 ����S0�!����������������
?QY�B�S���1��� <-�� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O�OiCC�@XLM�T��C�  ��DIN�O�A�Dq�EXE�HPV_���ATQz
��L�ARMRECOV� �RgLM_DG *�5���OLM_IF 	*��`d�O�_�_�_ �_j�_'o9oKo]onm, 
��odb���o�o�o�o^��$� yz, A   2�D{�PPINFO7 u[ �Vw��������`� ������*��&��`�J���n�����DQ� ���
��.�@�R��d�v���������a
P�PLICAT��?��P��`�Handlin�gTool 
� �
V8.30P�/40Cpɔ_LI
883��ɕ$ME
F0G��4�-

39�8�ɘ�%�z�
?7DC3�ɜ^
�NoneɘVr����ɞ@6�d� Vq_ACT#IVU��C죴�MODP���C�I��?HGAPON����OUP�1*�� i�m�����Қ_����1*� ) �@������� ��Q���Կ�@�
������ ���5�Hʵl�K�HTTHKY_� �/�M�SϹ������� ��%�7ߑ�[�m�� �ߣߵ���������� !�3��W�i�{��� ������������/� ��S�e�w��������� ������+�O as������ �'�K]o �������� /#/}/G/Y/k/�/�/ �/�/�/�/�/�/?? y?C?U?g?�?�?�?�? �?�?�?�?	OOuO?O QOcO�O�O�O�O�O�O �O�O__q_;_M___ }_�_�_�_�_�_�_k�ƭ�TOp��
�DO?_CLEAN9�ꤾpcNM  !{ 衮o�o�o�o�o��DSPDRYRwo&��HI��m@�or ����������&�8�J���MAX@ݐWdak�H�h�XWd��d���PLUG�GW�Xgd��PRC*)pB�`�kaS��Oǂ2DtSEGF0�K� �+��o�o�r����������%�LAPOb�x�� �2� D�V�h�z�������¯�ԯ�+�TOTAL�����+�USENU
O�\� e�A�k­��RGDISPMM�C.���C6�z�@I@Dr\�OMpo�:��X�_STRING� 1	(�
�kM!�S�
���_ITEM1Ƕ  n������+� =�O�a�sυϗϩϻπ��������'�9��I/O SIG�NAL��Tr�yout Mod�eȵInpy�S�imulated�̱Out���OVERRLp =� 100˲In� cycl�̱�Prog Abo�r��̱u�Sta�tusʳ	Hea�rtbeatƷMH Faul	��Aler�L�:� L�^�p��������� ScûSaտ ��-�?�Q�c�u����� ����������)�;M_q��WOR .�û������ +=Oas� ������//'.PO����M � 6/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l?�~?�?�?�?�?H"DEVP.�0d/�?O*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_>n_PALT	��Q �o_�_�_�_�_oo )o;oMo_oqo�o�o�o��o�o�o�o�_GRIm�û9q�_as �������� �'�9�K�]�o�������'�R	�݁Q�� ��)�;�M�_�q��� ������˟ݟ����%�7�I�ˏPREG �^����[�����ͯ߯ ���'�9�K�]�o� ��������ɿۿ�Oݿ�$ARG_� D ?	���0���  �	$O�	[�D�]D��O�e�#�S�BN_CONFIOG 
0˃����}�CII_SA_VE  O������#�TCELLSETUP 0��%  OME_I�OO�O�%MOV�_H������REP���J��UTOBA�CK�����FRA:\o�c Q�o���'`�йo���� �� f�o�����*�p!�3�`�Ԉ��f� ����������o�{� �&�8�J�\�n���� ��������������" 4FXj|�������끁 � ��_i�_\AT�BCKCTL.T�MP 6.VD �GIF .TP �D_q��N.sE#��f�INI�P��Օ�c�MESSAG�����8��ODE_D����z���O�0�c�PAU�SM!!�0� (�73�U/g+(Od/�/x/�/�/�/�/ �/�/???P?>?t?�1�0$: TSK  �@-��T�f�UPD�T��d�0
&XWZD_ENB����6STA�0��5�"�XIS��UNT� 20Ž� �� 	 I�2�0�e���� ���z⶙�Eư2�џ�@�HsM�Oo�}C�5�� �D�O��O�O _�?5CMET�߀2CMPTA@4�;?���?��/�@5��@���@�]4���4��%4�cG.5q�24h�@4���8]�SCRDCFG }1�6����H _�_o@o(o:oLo��o�Q�� �_�o�o�o�o�o�o]o �o>Pbt��0�o9�i�GR<@MX/�s/NA�/�s	i��v_ED��1�Y� 
 ��%-5EDT-��'�GETDA�TAU�o�9�����?�j�H�o�f��\��A�􏕀��2`�&�!�E���:IB ބj��~�ŏ׏m����3��&۔��D_��ߟJ�����9�ǟ�4 ���ϯ�(����]�o�����5N����� �(�w��)�;�ѿ_��6ϊ�gϮ�(�C�@����ϝ�+��7�� V�3�z�(��z�����i����8��&���~�]���F�ߟ�5���B�9~������]�����Y�k�����CR�!ߖ���W�q����#�5���Y��p$�NO�_DEL��rGE?_UNUSE��t�IGALLOW �1��(�*SYSTEM*�S	$SERV�_GR�V� : REG�$�\� �NUM�
��P�MUB ULA�YNP\PM�PAL�CYC10#6 $\ULSU�8:!�Lr�BOX�ORI�CUR_���PMCNV6�10L�T4DLI�0��	����BN/`/r/�/��/�/�/�/���pLA�L_OUT ��;���qWD_AB�OR=f�q;0IT_R_RTN�7�o	�;0NONS�0�6� 
HCCFS_U?TIL #<�5�CC_@6A 2#; h ?�?�?O�#O6]CE_OPT;IOc8qF@�RIA_Ic f5�Y@�2�0F�Q�=2q&}�A_LI�M�2.� ��K �]B��KX�K 
K �2O�Q�R�B�r�qFK Q 5T1)TR�H�_:J�F_PARAMGoP 1�<g^�&S�_�_�_�_�VC��  C�d�`��o!o`�`�`�
`�Cd��Tii:ah:e>eBa�GgC�`~� D� D	�`m�w?��2HE �ONFI� E?�aG�_P�1#; ���o1C�Ugy�aKPAU�S�1�yC ,�������� �	�C�-�g�Q�w���@������я���rO�A��O�H�LLECT_�B�IPV6��EN. QF�3�ND�E>� �G�7�1234567890��sB�TR�����%
 H�/%) �������W���0� B���f�x���㯮��� ү+�����s�>�P� b����������ο� �K��(�:ϓ�^�|�:�B!F� �I|�IO #��<U%�e6�'�9�K���T-R�P2$��(9X�t�Y޼`%�̓ڥH���_MOR�3&��=�K XB2 �a��A�$��H�6� l�~���~S��'�=�r�_A?�a�a`��K K(��R�dP��)F�ha�-�_�'�9�%
�k��G� ��%yZ�%��`K ]c.�PDB��+����cpmidbag��	3 :��@%��@�QU��p��N�  �  +�o �/���V]܌0�0 w�<�^�`@N`��wg�$�V
`@Wwfl�q>��ud1:���:J��DEF *�ۈ��)�c�b?uf.txt�����_L64FIX ,������l/ [Y/�/}/�/�/�/�/ 
?�/.?@??d?v?U? �?�?�?�?�?�?,/>#__E -���<�2ODOVOhOzO�O6&I�M��.o�YU>�c��d�
�IMC��2/����dU�C���20�M.:Uw�Cz�  B�i�A����A�jA@���B3�*CG��B<�=w�i�B�.��B�v1B����B�$�D?�%B���ezV�Cit&C���C�n�D-lE\D�n أkJ��22o�D�|��0�0���0j� �� ����
ЙxObi�D4cdv`Dů�`/�`v`s]E��D D�` E�4�F*� Ec���FC��u[F����E��fE���fFކ3F�Y�F�P3�Z���@�33 ;��O>L���Aw�n,au@�0@e�5Y��H�a���`A��w�=�`<#���
��?�oz�JRSMOFST� (�,bIT1���D @3��
д�X���a��;��b�w?���<��M�NTEST�1O�CR@�4��>V�C5`A�w�Ia+ah�aORI`CTPB�U�3C�`4���r�0�:d����qI?�5���qT_�PROOG ��
�%$/�ˏ�t��NUSER�  �U������K�EY_TBL  �����#a��	
��� !"#$�%&'()*+,�-./��:;<=�>?@ABC�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~��������������������������������������������������������������������������������͓���������������������������������耇��������������������������LC�K�
����STA�T/��s_AUTO/_DO �	�c��INDT_ENB�P���Rpqn�`�T2����STOr`���;XC�� 26����8
SONY �XC-56�"b�����@��F( �А�HR5!0w���>�P�7b�t�Aff����ֿ� Ŀ����C�U�0� yϋ�fϯ��Ϝ�����p���-ߜ�TRL��oLETEͦ ���T_SCREEN� ��kc�s���U�MME�NU 17�� <ܹ���w����� ����K�"�4�� X�j���������� ��5���k�B�T�z� �������������� .g>P�t� �����Q (:�^p��� �/��;//$/J/ �/Z/l/�/�/�/�/�/ �/�/7?? ?m?D?V? �?z?�?�?�?�?�?!O �?
OWO.O@OfO�OvO��O�O(y��REG c8�y����`�M��ߎ�_MANUAyL�k�DBCO���RIGY�9�DBG�_ERRL��9��ۉq��_�_�_ }^QNUMLI�p�ϡ��d
�
^QP�XWORK 1:���_5oGoYoko}o�ӍDBTB_N� S;������ADB_AWA�YfS�qGCP r
�=�p�f_AL�pR��bbRY�[�
�WX]_�P 1<{y�n�,�%oc�P��h�_M��ISO��k@|L��sONTIMXכ�
���vy
���2sMOTNEN�D�1tRECOR�D 1B�� �<��sG�O�]�K� �{�b��������V�Ǐ �]����6�H�Z�� �������#�؟��� ���2���V�şz��� �����ԯC���g�� .�@�R���v�寚�	� ��п���c�χ�#� ��`�rτϖ�Ϻ�)� ��M���&�8ߧ�\� G�Uߒ�߶�����I� �����4�� �p7� n���ߤ������ ���"���F�1���|� �������[�����i� ��BTf���b�TOLERENC��dB�'r�`L���^PCSS_CCS�CB 3C>y�`IP�t}�~� <�_`r�K�� ���/�{��5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_��~�LL� D���fFY C�[C�`ZP^r_ +A� p� �sp���Q �\	 !A�p�Q�_�[? �_h�[oU�p��p��pSB�VHW�@�PWoio{h+�o�Xa�o�oY��[�	r�hN�>������AAs�<�h8<K��c���aD@VB���|�G����+��K� A�otGb^Gr�S�o����eB  _ =��Ͷa>�t&YB�� �pC�p�q
�aA"�H�S�Q-��q ���ud�v�����Af�P ` 0����D^P��p@�a
F�QX��\ a"W>� �a9P��b�e :�L�^�h���́Ha�R�Q�He�z�֟ �o\^��-�?��c��u����zCz��ů�b2�Щ�RE{�u��D��)�� ��S̡0��]�0�.��@����Q�p��F� X�ѿUҁп�VS���NSTCY 1)E��]�ڿ�� K�]�oρϓϥϷ��� �������#�5�G�Y��k�}ߏߒ��DEV�ICE 1F5� E_����	� ��?�6�c��V|㰟�����_HNDGD �G5�N`���R�LS 2H�ݠ��/��A�S�e�w����� ZPARAM I�����RBT [2K��8р<�߬O`pC�C��,`¢�P�Z�z��%>{�C*  �2�j�Edv�,`"nPB , s��M� }�gT�g��
B��!�bcy�[2Dch z����/���/gT#I%D��CǓ` b!�R��A���A,��Bd���A��P��_C14kP�!2�C��$Ɓ��]�ffA�À���B�� �| �0��/�/�T (�P5 4a5�}%/7/d?/ M?_?q?�?�?�?�?�? O�?OO%O7OIO�O mOO�O�O�O�O�O�O �OJ_!_3_�_�_3�_ �_�_�_�_o�_(oo Lo^oЁ=?k_IoS_�o �o�o�o�o�o�o #5G�k}�� �����H��1� ~�U�g�y�ƏAo�Տ ���2�D�/�h�S��� go����ԟ����ϟ� ��R�)�;���_�q� ���������ݯ�<� �%�7�I�[�m����� ����}�&��J�5� n�YϒϤϏ��ϣ�ѿ ������F��/�A� ��e�w��ߛ߭����� ����B��+�x�O�a� �����������,� ��%�b�M���q����� ����������L #5�Yk}�� � ��61 CUg����� ���	//h/���/ w/�/�/�/�/�/
?�/ .?@?I/[/1/_?q? �?�?�?�?�?�?�?O O%OrOIO[O�OO�O �O�O�O�O&_�O_\_ 3_E_W_�_?�_�_�_ �_�_"ooFo1ojoE? s_�_�om_�o�o�o�o �o0f=Oa �������� ��b�9�K���o��� Ώ��[o��(��L��7�I���m������$�DCSS_SLA�VE L��}�ё���_4D  љ�~�CFG Mѕ���������FRA:\ĐL�-�%04d.CS�V��  }�� ����A i�CHq�z������|�����"������Ρޯ̩硞Ґ-��*����_�CRC_OUT �N������_�FSI ?њ ����k�}� ������ſ׿ ���� �H�C�U�gϐϋϝ� ���������� ��-� ?�h�c�u߇߽߰߫� ��������@�;�M� _����������� ����%�7�`�[�m� ��������������� 83EW�{� ����� /XSew��� ����/0/+/=/ O/x/s/�/�/�/�/�/ �/???'?P?K?]? o?�?�?�?�?�?�?�? �?(O#O5OGOpOkO}O �O�O�O�O�O _�O_ _H_C_U_g_�_�_�_ �_�_�_�_�_ oo-o ?ohocouo�o�o�o�o �o�o�o@;M _������� ���%�7�`�[�m� �������Ǐ����� �8�3�E�W���{��� ��ȟß՟���� /�X�S�e�w������� �������0�+�=� O�x�s���������Ϳ ߿���'�P�K�]� oϘϓϥϷ������� ��(�#�5�G�p�k�}� �߸߳����� ���� �H�C�U�g���� ���������� ��-� ?�h�c�u��������� ������@;M _������� �%7`[m ������� /8/3/E/W/�/{/�/ �/�/�/�/�/??? /?X?S?e?w?�?�?�? �?�?�?�?O0O+O=O OOxOsO�O�O�O�O�C��$DCS_C_�FSO ?�����A P �O�O_?_ :_L_^_�_�_�_�_�_ �_�_�_oo$o6o_o Zolo~o�o�o�o�o�o �o�o72DV z������� 
��.�W�R�d�v��� ����������/� *�<�N�w�r������� ��̟ޟ���&�O� J�\�n���������߯ گ���'�"�4�F�o� j�|�������Ŀֿ�������G�B�T��OC/_RPI�N_j� �����ς��O����1�XZ�U��NSL��@&� h߱���������"�� /�A�j�e�w���� ����������B�=� O�a������������� ����'9b] o������� �:5GY�} ������// /1/Z/U/g/y/�/�/ �/�/�/�/�/	?2?-? ??Q?z?u?��ߤ߆? �?�?�?OO@O;OMO _O�O�O�O�O�O�O�O �O__%_7_`_[_m_ _�_�_�_�_�_�_�_ o8o3oEoWo�o{o�o �o�o�o�o�o /XSew��� �����0�+�=� O�x�s���������͏ ߏ���'�P�K�]��o����� �PRE_?CHK P۪��A ��,8��2��� 	 18�9�K���+�q� ��a�������ݯ�ͯ �%��I�[�9���� o���ǿ��׿���)� 3�E��i�{�Yϟϱ� ������������-� S�1�c߉�g�y߿��� �����!�+�=���a� s�Q�������� ������K�]�;��� ��q������������� #5�Ak{� ����� CU3y�i�� ����/-/G/ c/u/S/�/�/�/�/�/ �/??�/;?M?+?q? �?a?�?�?�?�?�?�? �?%O?/Q/[OmOO�O �O�O�O�O�O�O_�O 3_E_#_U_{_Y_�_�_ �_�_�_�_�_o/oo SoeoGO�o�o=o�o�o �o�o�o=- s�c����� ��'��K�]�woi� ��5���ɏ������� �5�G�%�k�}�[��� ����ן�ǟ���� C�U�o�A�����{��� ӯ����	��-�?�� c�u�S�������Ͽ� ������'�M�+�=� �ϕ�w�����m���� ��%�7��[�m�K�}� �߁߳��߷����!� ��E�W�5�{��ϱ� ��e�������	�/�� ?�e�C�U��������� ������=O- s����]�� ��'9]oM �������/ �5/G/%/k/}/[/�/ �/��/�/�/�/?1? ?U?g?E?�?�?{?�? �?�?�?	O�?O?OO OOuOSOeO�O�O�/�O �O�O_)__M___=_ �_�_s_�_�_�_�_o �_�_7oIo'omoo]o �o�o�O�o�o�o! �o1W5g�k} ������/�A� �e�w�U�������я ��o����	�O�a� ?�����u���͟��� ��'�9��]�o�M� ��������ۯ��ǯ� #�ůG�Y�7�}���m� ��ſ�����ٿ�1� �A�g�E�wϝ�{ύ� ������	�߽�?�Q� /�u߇�e߽߫ߛ��� �����)���_�q� O���������� ���7�I���Y��]� ��������������! 3WiG��} ����%�A �1w�g��� ���/+/	/O/a/ ?/�/�/u/�/�/�/�/ ?�/9?K?�/o?�? _?�?�?�?�?�?�?O #OOGOYO7OiO�OmO �O�O�O�O�O_�O1_ C_%?g_y__�_�_�_ �_�_�_�_o�_+oQo /oAo�o�owo�o�o�o �o�o);U__q ������� �%��I�[�9���� o���Ǐ�����ۏ!� 3�M?�i��Y����� ��՟�ş����A� S�1�w���g�����������ӯ�+�=��$�DCS_SGN �QK�c��7m�� 18-J�AN-19 12?:59   O�l�}4p�08:38}������ N.DѤ���������h��x,rWf*�o��^M��  O��VERSION �[�V3.�5.13�EFLOGIC 1RK���  	���P�?�P�N��!�PROG_EN/B  ��6Ù��o�ULSE  �TŇ�!�_ACC�LIM�����Ö��WRSTJ�NT��c��K�E�MOx̘��� ���I?NIT S.�G��Z���OPT_SL� ?	,��
 ?	R575��YЫ74^�6_�7_�50��1��2_�@ȭ�|�<�TO  H�跿��V�DEXҚ�dc����PA�TH A[�A�\�g�y��HCP�_CLNTID y?��6� @�������IAG_G�RP 2XK� ,`� ��� �9�$�]�H������1234567890����S�� |�������!�� ��H���@;�dC�S���6 �����.� Rv�f��H ��//�</N/� "/p/�/t/�/�/V/h/ �/?&??J?\?�/l? B?�?�?�?�?�?v?O �?4OFO$OjO|OOE� �Oy��O�O_�O2_���_T_y_d_�_,
�B^ 4�_�_~_`O o�O&oLo^oI��Tjo �o.o�o�o�o�o �O '�_K6H�l� ������#���G�2�k�V���B]���}OF�ƠV��ۣf��� ?�{#�>!6�=��2�>+���{O�B_�
���G�� �Ƈ����(��L�B\�ډC*�@�b�.f�>���:������ߟʟܟ���C�T_CONFIG� Y��Ӛ��egU���ST�BF_TTS��
@��b����Û�u�O��MAU��|��MS/W_CF6�Z��6�~�OCVIEW��3[ɭ������ -�?�Q�c�u�G�	��� ��¿Կ������.� @�R�d�v�ϚϬϾ� ������ߕ�*�<�N� `�r߄�ߨߺ����� ����&�8�J�\�n� ���!���������� ���4�F�X�j�|�����RC£\�e��! *�B^������C�2g{�SBL_FAULT ]��|ި�GPMSKk���*�TDIAG �^:�աI���UD1: 67�89012345�G�BSP�-? Qcu����� ��//)/;/M/t
J��
@q��/$��TRECP��

 ��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOi/{/�xO�/UMP_OP�TIONk���AT�R¢l��	�EPM�Ej��OY_TEM�P  È�33B�J�P�AP�D�UNI��m�Q��Y�N_BRK _�ɩ�EMGDI_STA"U�aQK�XP�NC_S1`ɫ ��FO�_�_�^
�^d pOoo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{�E �����y�Q�� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d��z����� ��˟����%�7� I�[�m��������ǯ ٯ����!�3�E�W� i���������ÿݟ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�{�iߗ� �߻�տ������'� 9�K�]�o����� ���������#�5�G� Y�s߅ߏ�����i��� ����1CUg y������� 	-?Qk�}�� �������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?u?�?�?�?� �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_m?w_ �_�_�_�?�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9Ke_W����_ �_����#�5�G� Y�k�}�������ŏ׏ �����1�C�]o y��������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;���g�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�_� i�{ߍߟ߹������� ����/�A�S�e�w� ������������ �+�=�W�E�s����� �ߧ�������' 9K]o���� ����#5O� a�k}�E���� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-?GYc?u?�? �?��?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ Q?[_m__�_�?�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/I_Sew ��_������ �+�=�O�a�s����� ����͏ߏ���'� A3�]�o������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����9�K�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� ��C�M�_�q߃ߝ��� ����������%�7� I�[�m������� �������!�;�E�W� i�{��ߟ��������� ��/ASew ������� 3�!Oas��� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?+=G? Y?k?!?��?�?�?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O 	_#?5??_Q_c_u_�? �_�_�_�_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o-_7 I[m�_���� ����!�3�E�W� i�{�������ÏՏ� ���%/�A�S�e� q�������џ���� �+�=�O�a�s����� ����ͯ߯���� 9�K�]�w��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� �����'�1�C�U�g� ���ߝ߯��������� 	��-�?�Q�c�u�� ����������m�� )�;�M�_�y߃����� ��������%7 I[m���� ����!3EW q�{������ �////A/S/e/w/ �/�/�/�/�/�/�/ �/+?=?O?i_?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O��O�O�O? �$E�NETMODE �1aj5��  00�54_F[PRROR�_PROG %�#Z%6�_�YdUTA�BLE  #[�t?�_�_�_gdRSE�V_NUM 2R?  �-Q)`�dQ_AUTO_ENB  PU+SaTw_NO>a b#[�EQ(b  *�*�`��`��`��`4`�+�`�o�o�oZdHI�S%c1+PSk_AL�M 1c#[ �24�l0+�o;@M_q���o_b.``  #[aFR��zPTCP_VE/R !#Z!�_��$EXTLOG_7REQ�f�Qi,��SIZ5�'�STK�R�oe�)�TOoL  1Dz�b��A '�_BW�D�p��Hf��D�_D�I�� dj5�SdDT1KRņSTE�Pя�P��OP_�DOt�QFACTORY_TUN�g�d<�DR_GRP� 1e#YNad 	����FP��x�̹ ���� �$�f�?�� ��� ǖ��ٟ�ԟ���1� �U�@�y�d�v������ӯ����LW
 JG$�o�,��tۯ��j�U���y�B� � B୰���$ � A@��s�@UU�UӾ�������E��� E�`F@ �F�5U/�,��L����M��J�k�Lzp�JP��Fg�f��?�  s��9��Y9}�9���8j
�6̿�6�;���	�\�鉵 ��� 
H 	ȥ�ma͜[�FEATURE �fj5��JQ�Handlin�gTool � �"
PEn�glish Di�ctionary��def.4�D St�ard��  
! h�Analog �I/OI�  !�
IX�gle S/hiftI�d�X��uto Soft�ware Upd�ate  rt �sѓ�matic �Backup�3�\st��gr�ound Edi�t��fd
Camera`��Fd�e��CnrROndIm���3��Common calib UI��_ Ethe�n���"�Monitor��LOAD8�tr~�Reliaby��O�ENS�Data Acquis>���m.fdp�ia�gnos��]�i�D�ocument �VieweJ��8�70p�ual �Check Saofety*� cy�� �hanced Us��Fr�����C �xt. DI�O :�fi�� m�8���end��ErrI�L��S������s  t Pa��r[�� ���J9�44FCTN_ Menu��ve��M� J9l�TP �InT�fac{� � 744��G��p� Mask Ex�c��g�� R85��T��Proxy� Sv��  15� J�igh-S�pe��Ski
� �R738Г��m�munic��on�s�S R7��uqrr�T�d�022���aю�connecwt 2� J5���Incr��str�u,Қ�2 R�KAREL Cmod. L��ua���R860hRunw-Ti��EnvL��oa��KU�el u+��s��S/W����7�Licensye���rodu� �ogBook(S�ystem)�A�D pMAC�ROs,��/Of�fs��2�NDs�M�H�� ����M�MRC�?��ORD�E� echSto�p��t? � 84�fMi$�|� 13dx��]е�׏����Modz�witc�hI�VP��?��.� sv��2Op�tm�8�2��fi�l��I ��2g �4 !+ulti�-T�����;�PCM funY�Po|���4$�b&/Regi� r �Pri��FK+7����g Num Se-lW  F�#��� Adju���6�0.��%|� fe<���&tatu�!$�6���%��  9 �J6RDM �Robot)�sc�ove2� 561N��RemU�n@�� 8 (S�F3Se�rvo�ҩ�)�SNPX b<�I�\dcs�0}��Libr1��H� �5� f�0��[58��So� tr��ssag4%G 91��p ��&0����p/I��  (�ig TMILIBx(MӋ�Firm�����gd7���s�Ac�c����0�XATX��Heln��*LR�"1��Spac��Arquz�imu�laH��� Q���Tou�Pa��I���T��c��&��ev�. f.sv?USB po��"��iP�a��  r�"1Unexcep�t��`0i$/����H[59� VC&�r��[6���P{��RcJ�PRIN�V�; d� T@�TSP C�SUI�� r�[X�C��#Web P9l6�%d -c�1R�@4d�����I�R66?0FV�L�!FV�GridK1play C�lh@���і5RiR�R.@���R-35iA���Ascii���"�η� 51f�cUp9l� � (T�����S��@rityA?voidM �`���CE��rk�C�ol%�@�GuF� 5P��j}P����
 B�zL�t� 120C C� o�І!J��P�Бy��� o=q�b �@DCS b ./��c��O��q��`�;� ���qckpaboE4�DH@�OT�~��main N��r�1.�H��an.�t�A> aB!FRLM����!i ���MI 7Dev�  (�1�G h8j��spiJP@��� �@��Ae1/�r����!hP� M-A2� i��߂^0i��p6�PC��  �iA/'�Pass�wo�qT�ROS� 4����qeda�SN��Cli�����G6x Ar�� 47��!���5s�DER\��Tsup>RtОI�7 (M�a�T2�DV�
�3D Tri-���&��_�8;�
�A�@Def�?����Ba: d7eRe p 4t0���e�+�V�st6�4MB DRAM��h86΢FR�O֫0�Arc� v#isI�ԙ�n��7|� ), �b�He�al�wJ�\h��C'ell`��p� �sh[��� Kqw�c�� - �v���pX	VCv�tyy�s�"^Ѐ6�ut� �v�m���xs ���TD_0��J�m�` �2��a[�>R ts=i�MAILYk��/F2�h��ࠛ 9�0 H��F02]�q2�P5'���T1C��5���@FC��U�F�9�GigEH�S�t8�0/A� if�!2v��boF�dri=c� �OLF�S�����" H5k�OgPT ��49f88���cro6���@��l�ApA�Sy�n.(RSS) �1L�\1y�rH�L� �(2x5�5�d�pCV�x9����est�$S�Р��> \pϐSS�F�e$�tex�D �o���A�	� BP����a�(R00�Qi#rt��:���2)�D���1�e�VKb@l �Bui, n��WACPLf��0��Va��kT�XCGM��D��L8����[CRG&a&�YBU��YKfL�p�pf��k�\sm�ZCTAf�@�О�Bf2�и��V#�s���� r���CB���
Pf���WE��!��
���T�p��DT�&4 Y�V�`���EH����
�61�Z��
�R=2�
�E 	(Np��F�V�PK�B����#��Gf1`?GD���H�р?I�e ����LD�L��N��7\s@���`����M��dela�<,��2�M�� "L[P��`?��_P�%�����S��-F��TSO�W�J5�7��VGF�|�V;P2֥ 5\b�`0�&�cV:���T;T�� �<�ce,?V{PD��$
T;YF��DI)�<I�'a\so<��a-�6J�c6s6�4L�M�V9R�h���Tri�� ���5�` �f�@��������P
� ����`��IOmg PH�[l�6�I/A  VP�S��U�Ow��!%S|�Skastdpn)���t�� SWIMEkST�BFe�00��-Q� �_�PB�_�RGued�_�T�!�_��S ��_bH573�o2c2��-oNbJ5�N�Iojb)�Cdo�cx E��o�_�lp��o�TdP �o�c�B�or�2.r�ٱ(Jsp�EfrSE�o�f1�}�r3 R�GoeELS��sL ����s�����B	�0�S\ $�F�ryz�ftl�o~�g�o����������?�����P   �n�&�"�l ��T �@<�^��Y��e�uy8Z���alib���Γ��ɟ3���埿�\v ��e\c�6�Z�qf�T�v�R VW�r��8S��UJ91��0��i�ů[c91+o�wy8���847� :��A4�j��Q��t6�<m���vrc.����0HR���ot�0ݿN��  ��8ޯf�460�>eS0L�97���U�ЄϦ�60.� g�н�+���'�ܠ�Ϻ�8co��D	M߱U"�����ߕp�i�߲T! ��n	a;�� ���u%��ⅰI��loR�d��1a59gϱŭ�&��95�ϔ�R����1��?��o�#��1A��/���vt{�UWe0ǟ���ￇ73[���97�ρ�C W���62K�=fR���8���������d����2 �ڔ����@�@y" "http������t7 �� v 3R7��78�����4�� ��TTPT��#	��ePCV�4/v߀�j�Q�Fa�7��$N�0�/2�rI�O�)/;/M/6.sv�3�64i�oS�l? torah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4c.K?�g'�)�s24g?�� (B�O�d�\iOA5sb�?U_�?vi�/i��/��/Wn��`�o%�F o�4l�$of��oXF� I)xo�cmp\�7��mp���duC`��lh����o(A�_Bt� �o]6P��m�I?0�w�@���naO��	4*O0wi�%P�?"�bsg?�]7�YE$M���8woVJ�/ե311?o��DMs�BC��7J�\���r(�52�XFa AP��ڟ<�v�`/şaqqs����/Of���1�9�VR`K���ph�քH5+��=�IN/¤SkiW�/�IF��_�%��fs�I�O�l����"<𜿚$�`�����\jԿz5bO�vr�ouς�3(�ΤH (DϮ��?sG��|� �F�Ou�������D)O��*�3P$�FӅ�@k��ϻ���럴� �P�L��ʿ��pbox��ߦebo���Sh$ �>�R.�0wT{����fx6��P��D`��3��#_I\m;YEe�OԆM�hxW��=Ete,���dct\���O$kR���d���Xm*���ro30��D�l�j9��Vx'�  FC����|@�ք f?6K�ARE0�_�~ (1Kh��.cf����WpoO�_K�up���a���H/j#- 3Eqd/�84���$qu�o��/ o2o?DVo<�7C�)�s�NJ�Ԇ�|?�3l\sy`�?�40�?Τwio��u]?�w58�?,F�a$OJ�
?Ԇ"io��!�V��u&A��P�R�ߩ5, s��v1�\  Hg552B�Q21p�0R78P5�10.R0  n�el J61�4Ҡ/WA�TUP��d8P54�5*�H8R6��9_VCAM�q97P�CRImP\1tPUI�F�C8Q28  i�ngsQy0��4P P6�3P @P PSCH~��DOCVڀD �PCSU���08Q�0=PqpVEIcOCr��� P54Pwupd�PR69aP܄��PSET�pt\!hPQ`Qt�8P7`Q�!?MASK��(P?PRXY���R�7B#POCO  /\pppb36���@PR�Q��b1Pd60Q^$cJ539.eHsb~��vLCH-`~(�OPLGqK\bPQ0]`��P(`GHCR��4`S�awund�PMCSIPR`e0aPle5=Ps�p(`DSW� �  qPb`0`�aPa��(`PRQ``Tq�RE`(Poa601P�<cPCM�PHcR0@q\j23b�V�`pE`�S`UPvisP�`E` c�`UPcPR9S	a�bJ69E`s�FRDmPsRMC�N:eH931PHcS�NBARa�rHLB��USM�qc�Pg5�2�fHTCIP0cT�MIL�e"P�`eJ� �PA�PdSTPT�X6p967PTEL��p��P�`�`
Q8P8$Q48>a"PPX�8Pc95�P`[�95qq�bUEC-`F
�PUFRmPfahQCvmP90ZQVCO�`�@PVIP%�53�7sQSUIzVSX��P�SWEBIP�SH�TTIPthrQ6�2aP�!tPG���cI�G؁�`c�PGSξeIRC%��cH7�6�P�e Q�Q|�Ror��R51P s:PL�P,t53=P8u8=P
y�C�Q6]`�b�P�I��q52]`sJ5�6E`s���PDsCLt�qPt5�\rd�q375UP cR8���u95P sR55]`,s � P8s��P�`CP�P�P�SJ77P0\o�6��cRPP�cR6�ap�`�QtaT�379P`�64�Pd387]`�d90P0c ��=P,���5�9ta�T91P� ��1P(Sܒ��Qpai�P06�=P- C�PF�T`	���!aLP PTS�p.L�CAB%�I Б�IQ` ;�H�UPPa[intPMS�Pa�иD�IP|�STY%�t7\patPTO�b8�P�PLSR76�`�5�Q��WaNN�Pa�ic�qNNE`�OsRS�`�cR681Pwint'�FCB�P"(�6x�-W`M�r���!(`OBQ`pluug�`L�aot �`GOPI-���PSP�Z�PPG�Q7�`7�3ΒPRQadv�RL��(Sp�P�S��n�@�E`��� �PTS-��q W��P�`apw�`8��P`cFVR�Plc�V3D%�l�PBV�I�SAPL�Pcy�c+PAPV1�pa�_�CCGIP - uU��L�Prog+PGCCR�`�ԁB�Pi �PԁK=�"L�PH��p��(h�<�P���h�̱�@g�Bـ
�TX�%���CTC��ptp��2��P927"0ҝPs2�Qb��;TC-�rmt;�	`�#1ΒTC9`HcC[TE�Perj�EIPp.p/�E�P�c�ЮI�use��Fـverv�F%���TG�Pp� CP��%�d -h��H-�Tra�PCT�I�p��TL� TRS���p�@נ��IP�PTh�M%�lex�sQTMQ`ver, �p�SC:���F��P�v\e�PF�IPSV�"+�H�$cj�ـtr��aCTW-���CPVsGF-��SVP2mPOv\fx���pc�bؚ�e��bVP4�fx�_m��-��SVPD�-��SVPF�P_m�o�`V� cV��t�\��LmPove4���-�sVPR�\t|�tPV�Qe5.W`V6�*u"��P}�o`�М�`��CVK��N�I�IP��CV����IP=N9�Gene���D���D�R�D����  ��f谔�pos.^��inal��n�D�DeR���`��d�P��omB���on,����R�D�R��\��T�Xf��D$b��omp��� "N��P��m����! ��=C-qf����=FXU�����g F��(��Dt II��r�D���u�� "����Cx_ui X�������f2��h	Crl02��D,r9ui�Ԣ>� it2c�0�co��e"���Խا(.)� ����� ���� IQnQ �{I[ ��_= �wo��,bD�� ��|GG�� �����{4 �e� �vʷ� ��&�� 2��Z u{z������ ��TW&q~q� 5�׷&�o�? ;0��  ��2� �y�� ���W&��� ?�3� {A��e�/> ��\�3&T���� 77߸ ��{�� ���� �ֵ��&��8� �l1��S��) ���d *�J� F's� ~��� 6:0ݙ ��,��s�{�- Q�v� ���� �,սT �ZBLx6�ۯ�6 ��6����Par ��s�>�E��j�6dsq��F  ���������Dhel�����ti-S�� �Ob��Dbcf�O���V��t OFT��P< A�_�V�ZI��D���V\�qWS��= d7tle�Ean�(b{zd��titv�JZ�z�Ez XWO� H6�6���5 �H�6H691�E4܀TofkstF� Y�682�4�`�f8�04�E91�g�`3<0oBkmon_�E��xeݱ�� qlm��W0 J�fh��B�__  ZDTfL0��f(P7�Eckl`KV� �6|��D85��ّ�m\b����xo܊k�ktq��g2`.g���yLbkLV�ts��IF�bk������Id I/�f��GR� �han�L��Vy��%���%ere�����io��� ac�- A��n�h���cuA2Cl�_�^ir��)�dg��	.�@�& G��R630���p v��p�&H�f��un���R57v�OJa�vG�`Y��owc��-ASF��O��7���SM������
af��rafLa�vl�\F c�w a���?VXpoV� �30��NT "L�FFM��=����yPh	a�G-�w�� �m2.�,�t��̹π6ԯ��sdF_�MC'V����D����fslm�is�c.  �H5522��21�&dc.pR7�8����0�708J614V�ip ATUtu�@�OL�545Ҵ�INTL�6�t8 ?(VCA����sseCRI���ȑ��UI���rt�\rL�28g��N�RE��.f,�63�!��,�SCH�d =Ek�DOCV���p���C,�<�L�0Q�i;sp��EIO��xEF,�54����9���2\sl,�SETp���lр�lt2��J7�ՌMA�SK��̀PR�XY҇��7���O[CO��J6l�3�<l�� (SVl�A��H�L�@Օ��539fRsv���#1���LCH���OPL]Gf�outl�0���D��HCR
sv�g��S@�h��CSa�!�{�50��D�l�q5!�lQ��DSW��aS����̀��OP����7��PR���L<�ұ�(Sgd���gPCM���R0 �\s��5P՝���0����n�q� AJ�1��N�q�2��PRS�a���69�� (A?uFRD�Խ���RMCN���9�3A�ɐCSN�BA�F9� HLB��� M��4���h��2A�95z�HTC�aԈ�TMIL6�j�95,��857.v,PA1�ito��oTPTXҴ JK�'TEL��piL��i XpL�80�I)��p.�!��P;�J95�ԏs "N���H�U{EC��7\cs��FR��<Q��C��5;7\{VCOa�,����IP1jH��S;UI�	CSX1�A�WEBa��HsTTa�8�R62���m`��GP%�IG� %tutKIPG�Sj�| RC1_m�e�H76��7�P�ws_+�?x�R;51�\iw�N�L��H�53!��wL�98!�h�R66��H����Ԡ���@;J56��1���N0��9�ej��L���R5`%��A|�5q�r�`,�8 5��{165!��@�"�5��H84!�29���0��PJ���n; B[�J77!ԨӃR6�5h3n���y36P��3R6��-`;о pԨ@��exeK�J87��#J90�!�stu+�~@!�۵�k90�koAp�B����@!�p�@|BA�g*�n@!��Q��#06!�@[�F�FaPb�6��́,�TS�w NC[�CAB$iiͰl1I��R7��p@q�y�CMS1�rog+QM�� �� sTY$x�CTOa�nv\+��1�(�,�6�con�~0�Ի15��JNN�%ep:��P��9ORS%tx���8A�815[�FCBaUnZQ�P!�p�p{��CMOB���"G��OL��x�O�PI�$\lr[�S�Š�T	D7�U��CP�RQR9RL���S��V�~`���K�ETS�$1��0���3\�Ԩ�FVR1�LZQ�V3D$ ���BV�a�SAPL1�CL�N[�PV��	rCC1Gaԙ��CL�3�CCRA�n "Wr!B�H�CSKQ�n\0�p��)�0CTPn�ЌQe��p.!$bCt�aT0U��pCTC�yЋRC�1�1 (�s��trsl,�r��
TX��;TCaerrm�r��MC"�s��#CT]E��nrr�REa��XPj�^��rmcH�^�a"�P�QF!$����$p "�rG,1�tTG$c8��Q�H�$SCTI�!� s��CTLqdACCK�Rp)��rLa�R82��M��YPk�.���OF��.���e��{�CN���^�1�"M�^�a�С�Q`US���!$��M�QW�$m�VGF�$R M�H��P2�� H5�� ΐq��ΐ�$(M-H[�VP�uoY���h�$)��D��hg���VPF��"MHG�̑`e!�+�V/vpcm�N��ՙ�N��$��VPRqd)��CV�x�V� "�X�,�1��($TIa�t\mh:��K��etpK��A%Y�VP%ɠ�!PN����GeneB�rip����8��extt���Y�m�"�(��HB� ��)��x��������Ȣ�res.�yA�ɠn����*���p�@M�_�N��6L���Ș�yAvL�Xr�Ȉ2��"R;�Ƚ\rax��	P�� h86���Gu+ʸ�Ͽ�Se0Lɨm�9�69�P����r�Ȩ2�ɹ1��n2��h� �0L�XR}�R�I{�e� L�x���c �Ș���N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1��/�k�@���A���ruk�ʘ L�scop��H�}�ts{������s��9��j7965��Sc��h���5 J9�{�
t�PL�J	een���t I[
x�comr��Fh�L�4 J���fo��DIF�+�6�Q����rat�i|��p��1�0�
R	8l߾�M�����PB��8� �j�mK�@X�HZ����N��oڠ��3�q��v�i���80�~�l� Sl�yQ��tpk�xb�j�.�@�R� d������,/n(�8�A8�0���
:�O8��<�Q}�CO���PT.��O (��.�Xp�|�~H���?�v� �wv��8�228�pm���722�j7�^�@ƙ���c�f�=Yvr���vcu���O�O�O�O�_#_5_7�3Y_��w3v4{_�_w�ʈ��ust_�_�cus�_�Z��oo,o>opPo�io��nge���(pLy747�jWe�lʨHM47ZKE�q {���[m�MFH�?�(wsK�8J��n���o��fh9l;��wmf���?� :�}(4	<g 9J{��II)̏މ9w��X�774kﭏ&/7ntˏ݊e+���3se�/�aw��8ͤɐ��EX \�!+: X�p��~�00��nh��,:Mo+�xO��1 �"K�O��\a��# 0��.8���{h�L?��j+�mon�:��tL�/�st�?-�w�: ���)�;��(=h��;
d Pۻ�{: 7 ��� �J0֛�re�����STD�!treLANG���81�\tqd����<���rch.��x����htwv��WWָ� R79��"Lo�51 (�I�W�h�Ո�4֧aww� �v�y �623c�h a?�cti�֘!�$X�iؠ�t �Ձn,�։����j<��"AJP@�3�p�vr{�H�6��!���- SeT� Ex3�) G�J934��{LoW�4 (S������� <���91 ��8!4�j9�所+�d��y�
��	�btN�ite{�R ��I@ Ո�����P��������	 ����Z�vol ��X ��9�<�I�p����ld*���F�86!4{��?��K�	��k扐�֘1�wmsk��M�q�Xa�Ae����p���0RBT�1ks.?OPTN�qf��U$ RTCam T��y��U��y�� U��UlU6L�T@�1Tx����SFq��Ue�6T��USP; W�b DT�qT2h�T�!/&+��8TX�U\j6&��U U�Usfd�O&�&ȁT���662DPN�abi��%�Q�%62V� �$���%�� �#(�(6{To6e St�%���#5y�$�)5(To�%tT0�%5�W6�T���%�#�#orc���#I���#���%c�ct�6ؑ?�4\W6965"p6}"�#\j536���4�"��?kruO O,Im ?Np�C �?t�0<O�;�e �%���?�
;gcJ7 "AV<�?�;avsf�O__&_8WtpD_V_0GT�F|_:UcK6�_�_9r�O�3e\s�O2^�y`O:�migxGvNgW! m�%��!�%T�$E A{6�po6̀�#37N�)5R5�_2E���$0���$Ada�Vd���V�?;Tpz7�_�e7DDTF9���#8�`�%��4~y�ted Z@0�A}�@�}�04N�}�0}���}�dc& }����u 6�v��v1�u1\b�u$2}�<��}� R83�u�"x}��"}�valg���Nrh�&�8�J��Y�o�ue��� j7q0�v=1��MIG�uerfa��{q����E�N�ء��EYE�ce A���� �pV�e�A!���2Յ�Q �%��u1�e�i�@��@H�e����J0� '��b��T��E In��B�  W�|��5�37g����(MI�t�Ԇr��ݟ�Cam���nеv!g�U -�v J߆8⹖0F���P�y�ac���28���Rɏ jo��2�� djd�8r}�� og\k�0��gܕ�wmf�Fro/� Eq'�4"}��3 J8��oni[��ᅩ}Ĵ��C o� ��ʛ��m@�R�e��{n�Д�V��o������  �����裆"P�OS\����ͯ mcenϖ�⑥OMo��43��� �(Coc� An[�t���"Fe�a\�vp��.��ocflx$�le��`8�hr�tr�NT�w CF+�x E/�at	qi�M�ӓxc�֌p�f�lx����Z�c�x��
0 h��h8f��mo��=� H����)� (�vSER�,���g�0߆0\�r�vX�= ��I � - �ti��H���VC�828�5ص�L"�RC��n �G/���w�P�y�\v�vm "o�lϚ��x`��=e�ߠ-�R-3?������vM [��AX/2�)�S�r�xl�v#�0��h8�߷=� RAX�AТ����9�H�E/�Rצ����h߶"R�Xk��F�˦85ή�2L/�xB88�5_�q�Ro�0iA��5\rO�9�K��v����8���.�gn "�v��88��8s�i ?�9 �����/�$�y O�MS"����&�9R H784&�`�745�	pp��p��ycr0C�Rc�hP0� j�-�a�%?o��6D950R7tsrl��ctlO��APC���j�ui�"�L���  ����K^棆!�A��qH���&-^7����� ��616C�q�794h����� M�ƔI��99���(��$F�EAT_ADD �?	���Q~%P  	�H ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n���������TDEMO �fY   WM_��� �����//%/ R/I/[/�//�/�/�/ �/�/�/�/?!?N?E? W?�?{?�?�?�?�?�? �?�?OOJOAOSO�O wO�O�O�O�O�O�O�O __F_=_O_|_s_�_ �_�_�_�_�_�_oo Bo9oKoxooo�o�o�o �o�o�o�o>5 Gtk}���� ����:�1�C�p� g�y�������܏ӏ� ��	�6�-�?�l�c�u� ������؟ϟ���� 2�)�;�h�_�q����� ��ԯ˯ݯ���.�%� 7�d�[�m�������п ǿٿ���*�!�3�`� W�iϖύϟ������� ����&��/�\�S�e� �߉ߛ��߿������� "��+�X�O�a��� ������������� '�T�K�]��������� ��������#P GY�}���� ��LCU �y������ /	//H/?/Q/~/u/ �/�/�/�/�/�/?? ?D?;?M?z?q?�?�? �?�?�?�?
OOO@O 7OIOvOmOO�O�O�O �O�O_�O_<_3_E_ r_i_{_�_�_�_�_�_ o�_o8o/oAonoeo wo�o�o�o�o�o�o�o 4+=jas� �������0� '�9�f�]�o������� ��ɏ�����,�#�5� b�Y�k���������ş ����(��1�^�U� g������������� ��$��-�Z�Q�c��� ����������� � �)�V�M�_όσϕ� �Ϲ���������%� R�I�[߈�ߑ߫ߵ� ��������!�N�E� W��{�������� �����J�A�S��� w������������� F=O|s� ����� B9Kxo��� ���/�/>/5/ G/t/k/}/�/�/�/�/ �/?�/?:?1?C?p? g?y?�?�?�?�?�? O �?	O6O-O?OlOcOuO �O�O�O�O�O�O�O_ 2_)_;_h___q_�_�_ �_�_�_�_�_o.o%o 7odo[omo�o�o�o�o �o�o�o�o*!3` Wi������ ��&��/�\�S�e� ������������� "��+�X�O�a�{��� �������ߟ��� '�T�K�]�w������� ���ۯ���#�P� G�Y�s�}�������� ׿����L�C�U� o�yϦϝϯ������� �	��H�?�Q�k�u� �ߙ߫��������� �D�;�M�g�q��� ��������
���@� 7�I�c�m��������� ������<3E _i������ �8/A[e �������� /4/+/=/W/a/�/�/ �/�/�/�/�/�/?0? '?9?S?]?�?�?�?�? �?�?�?�?�?,O#O5O OOYO�O}O�O�O�O�O �O�O�O(__1_K_U_ �_y_�_�_�_�_�_�_ �_$oo-oGoQo~ouo �o�o�o�o�o�o�o  )CMzq�� �������%� ?�I�v�m����������ُ���;�  2�Q�c�u��� ������ϟ���� )�;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����� ��1CUg y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����'>9  :> Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{��������/=C6Yk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A���$FEAT_D�EMOIN  VE��q��>�Y�_INDEXf�u���Y�ILECOM�P g������t�T���S�ETUP2 h������  �N ܑ��_AP2�BCK 1i��  �)B���%�C�>���1�n� E����)���M�˯�� �����<�N�ݯr�� ����7�̿[��ϑ� &ϵ�J�ٿWπ�Ϥ� 3�����i��ύ�"�4� ��X���|ߎ�߲�A� ��e�����0��T� f��ߊ�����O��� s�����>���b��� o���'���K������� ��:L��p��� �5�Y�}�$ �H�l~�1 ��g�� /2/� V/�z/	/�/�/?/�/ c/�/
?�/.?�/R?d? �/�??�?�?M?�?q?@O�?O<O���P�� 2�*.V1RCO�O�0*�O�O`�3�O�O�5w@PC�O|_�0FR6:�O"=^�Oa_�KT���_ �_&U�_�\h�R_�_�6�*.FzOo�1	�(SoEl�_io�[STM �b�o�^+P�o��m�0iPen�dant Panel�o�[H�o �g��oYor�ZGIF |��e�Oa��ZJPG �*��e���z��JJS�����0�@���X�%
Ja�vaScriptُ�CSʏ1��f��ۏ %Casc�ading St�yle Shee�ts]��0
ARGNAME.DT��
�<�`\��^���Д�៍�АDISP*ן���`$�d��V��e��CLLB.cZI��=�/`:\���\�����Col�labo鯕�	P�ANEL1[�C�%��`,�l��o�o�2 a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V���zό��!ߘ�TPEINS�.XML(�@�:\�<����Custo�m Toolba�r}��PASSW�ORD���>FR�S:\��� %�Password Config� �?J���C��"O��3� ����i����"�4��� X���|�����A��� e�����0��Tf �����O�s ��>�b�[ �'�K���/ �:/L/�p/��/#/ 5/�/Y/�/}/�/$?�/ H?�/l?~??�?1?�? �?g?�?�? O�?�?VO �?zO	OsO�O?O�OcO �O
_�O._�OR_d_�O �__�_;_M_�_q_o �_�_<o�_`o�_�o�o %o�oIo�o�oo�o 8�o�on�o�!� �W�{�"��F� �j�|����/�ďS� e���������T�� x������=�ҟa��� ���,���P�ߟ񟆯 ���9����o���� (�:�ɯ^�����#� ��G�ܿk�}�ϡ�6� ſ/�l�����ϴ��� U���y�� ߯�D��� h���	ߞ�-���Q߻���߇��,��$FI�LE_DGBCK� 1i������ (� �)
SUMM?ARY.DG,���OMD:`�����Diag Su�mmary���
CONSLOG���y����$���Co�nsole lo�g%���	TPACCN��%g������TP Acco�untinF����FR6:IPKD?MP.ZIP�����
��)����Exc?eption-�����MEMCHEC�K�����8�M�emory Da�ta��LN�=)�RIPE����0�%� �Packet L�E���$Sn�S�TAT*#�� %LSta�tus�i	FTAP�/�/�:��mment TB�D=/� >)ETHERNE��/o�/�/��Et�hernU<�fi�guraL��'!DCSVRF1//)/�B?�0 verify allE?��M(5DIFF:? ?2?�?F\8diff�?}7o0CHGD1�?�?�?�LO �?sO~3&��
I2BO)O;O�O� bO�O�OGD3p�O�O�OT_ �O�{_
VUPDAT�ES.�P�_��FORS:\�_�]���Updates �List�_��PS�RBWLD.CM�o���Ro�_9�P�S_ROBOWEyL^/�/:GIG��o>_�o�Gig�E ��nosti�cW�N�>�)}�aHADOW�o�o�ob�Sha�dow Chan�ge��8+"rNOTI?=O���Notif�ic�"��O�A=�PMIO�o���h��f/��o�^U�*�UI3�E�W��&{�UI������B� ��f��_�������O� ��������>�P�ߟ t������9�ί]�� ���(���L�ۯp��� ���5�ʿܿk� Ϗ� $�6�ſZ��~��w� ��C���g���ߝ�2� ��V�h��ό�߰��� Q���u�
���@��� d��߈��)��M��� ������<�N���r� ���%�����[���� &��J��n� �3��i��" �X�|�� A�e�/�0/� T/f/��//�/=/�/��/�$�$FILE�_�PPR�P���� �����(MDONLY� 1i5�  
 �z/Q?�/u?�/ �?�?t/�?^?�?O�? )O�?MO_O�?�OO�O �OHO�OlO_�O_7_ �O[_�O_�_ _�_D_ �_�_z_o�_3oEo�_ io�_�oo�o�oRo�o vo�oA�oew �*��`�����&�O��*VIS�BCK,81;3*�.VDV����F�R:\o�ION\�DATA\��/���Vision� VD file ̏��&�<�J�4�n� �����3�ȟW���� ��"���F�՟�|�� ����m�֯e������ 0���T��x������ =�ҿa�s�ϗ�,�>� ��b���ϗϼ�K� ��o��ߥ�:���^�����ϔ��*MR2_�GRP 1j;��C4  B�}�	 71�������E�� E�  �F@ F�5U�������L����M��Jk��Lzp�JP���Fg�f�?� � S����9�Y�9}�9���8j
�6���6�;��A� � ���BH��B���B���$�������������@UUU#�����Y�D�}� h����������������
C��_CFG� k;T �M���]�NO {:
F0�� � \�RM_CHKTYP  0��}�000��O=M_MIN	x�g��50X� �SSBdl5:0��bx�Y����%TP_DEF'_OW0x�9��IRCOM���$GENOVRD�_DO*62�T[HR* d%d�o_ENB� �/RAVC��mK�� ��՚�/3�/���/�/�� ��M!OUW s���}��ؾ��8��g�;?�/7?Y?[? 7 C��0����(7l�?�<B�?B�����2��*9�N SMT�T#t[)��X�4�$�HOSTCd1u�x���?�� kMCx��;zO�x�  27.0z�@1�O  e�O �O	__-_;Z�O^_p_��_�_�LN_HS	anonymous�_ �_�_oo1o yO��FhFk�O�_�o�O�o �o�o�oJ_'9K ]�o�_���� �4o�XojoG�~�o ^�������ŏ��� ��1�T���y��� ��������,�>�@� -�t�Q�c�u������� ��ϯ���(�^�� M�_�q�����ܟ� � ݿ��H�%�7�I�[� ��ϑϣϵ����l� 2��!�3�E�Wߞ��� ¿Կ����
������ �/�v�S�e�w��� �����������+� r߄ߖ�s�����߻� ���������'9K ]�������� �4�F�X�j�l>�� }������ //1/T��y/�/��/�/�/.D\AENT� 1v
; P!\J/?  ��/ 3?"?W??{?>?�?b? �?�?�?�?�?O�?AO OeO(O�OLO^O�O�O �O�O_�O+_�O _a_ $_�_H_�_l_�_�_�_ o�_'o�_Koooo2o {oVo�o�o�o�o�o �o5�oY.�R�v��zQUICC0���3��tA14��"����t2���`�r�ӏ!ROU�TERԏ��#�!?PCJOG$����!192.168.0.10�~�sCAMPRTt�P�!d�1m������RT폟�����$N�AME !�*!�ROBO���S_CFG 1u�)� �A�uto-star�tedFTP&��=?/֯s�� ��0�B��f�x��� ������S������ ,���������ϼ�ޯ ���������ʿ'�9� K�]�oߒ�ߥ߷��� ������(:~� k�Ϗ�������� ����1�C�f���y� �����������,�>� R�?��cu�� `�����(� $M_q������  /H%/7/I/ [/m/4�/�/�/�/�/ �~/?!?3?E?W?i? ����?�/�?/�? OO/O�/�?eOwO�O �O�?�ORO�O�O__ +_r?�?�?�?�O|_�? �_�_�_�_o�O'o9o Ko]ooo�_o�o�o�o �o�o�oF_X_j_~o k�_������o ���1�TU��y����������U�)�_ERR w3�я��PDUSIZ  �g�^�p���>~�WRD ?r��Cq�  guestb�Q�c��u�������"�SCD�MNGRP 2x�r�����Cqg�\�b�K� 	�P01.00 �8(q   ��5p�5pz�5pB�  �{ ���H���L���L��L������O8�����l�����Ua4� x��Ȥ�x���8���\���)j�`�;�������d�.�@�R�ɛ__GROUېy�����	ӑ���QUPD  ?u�����İTYg�����TTP_A�UTH 1z��� <!iPen'dan��-�l����!KAREL�:*-�6�H�KC�]�m��U�VISION SET�� �ϴ�g�G�U������ R�0��H�Bߏ�f�x���ߜ߮���CTRL� {����g�
�S�FFF9E�3��AtFRS:DEFAULT;��FANUC �Web Server;�)����9�K� �ܭ���������߄�WR_CONFI�G |ߛ �;��IDL_CP�U_PCZ�g�B��Dpy� BH_�M�INj�)�}�GNR_IO��g���a��NPT_SIM_�D_�����STA�L_SCRN�� ����TPMODN�TOL������RT�Y��y���� �EN�O���Ѳ]�OLN/K 1}��M���������eM�ASTE��ɾeSLAVE ~��|c�O_CFG�ٱBUO�O@C�YCLEn>T�_?ASG 1ߗ+�
 ����/ /+/=/O/a/s/�/�/p�/�/��NUM���
@IPCH��^RTRY_CNZ���@��������� @kI��+E�z?E�a�P_�MEMBERS �2�ߙ� $���2���ݰ7�?�9a��SDT_ISOL�C  ����$�J23_DSM�+�3JOBPRO�CN��JOG��1�+�d8��?��+�O�/?
�LQ�O__/_@�OS_e_w_�_`�O� Hm@��E#?&BPO�SREQO��KANJI_���a[�?MON ����b�yN_goyo�o�o�oH�Y�`3�<� ��e�_ִ��_L���"?�`EYLOGGI�NLE��������$LANGUA�GE ��<�T� {q�LGa2��	�b���g�xP��W  ��g��'��b���>��MC:\RSCH�\00\<�XpN_DISP �+�G�J��O�O߃LOClp�Dz���As�OGBOOK ������󑧱����X�����Ϗ�����a�*��	 p�����!�m��!����=p_BUFF 1-�p��2F幟����՟D� Co�llaborativǖ���F�=�O� a�s�������֯ͯ߯����B�9�K���D�CS �z� =���'�f��?ɿۿ����H@{�IO 1�� ~?9ü��9�I�[�mρϑϣ� �����������!�3� E�Y�i�{ߍߡ߱���h�����E��TMNd�_B�T�f�x��� ������������,� >�P�b�t�������L�N�SEVD0��TYPN1�$6���QRS"0&��><2FL 1�"�J0��������GTP:pO}F�NGNAM1D��mr�tUPS�G�I"5�aO5�_L�OADN@G %v�%�pIND�`�5SE� ��$MA?XUALRM�'��8�(��_PR"4F0�d��1�B_PN�P� V 2�C�	MDR077�1ߕ�BL"80{63%�@ �_#�?�ߒ|/�C���z�6��/���/Po@Pw 2��+ �ɖ�	T 	t  ��/�%W?B?{? �k?�?g?�?�?�?O �?*OONO`OCO�OoO �O�O�O�O�O_�O&_ 8__\_G_�_�_u_�_ �_�_�_�_o�_4oo XojoMo�oyo�o�o�o �o�o�o0B%f Q�u����� ���>�)�b�M��� ��{��������Տ� �:�%�^�p�S��������D_LDXD�ISApB�ME�MO_APjE {?C
 �, �(�:�L�^�p�����~�ISC 1�C ����4��������4��X���C_MSTR ���~w�SCD 1���L�ƿH��տ��� 2��/�h�Sό�wϰ� ���Ͽ���
���.�� R�=�v�aߚ߅ߗ��� ��������<�'�L� r�]��������� �����8�#�\�G��� k��������������� "F1jUg� ������ B-fQ�u����h�MKCFG �����/�#LTAWRM_��7"�0�0N/V$� M�ETPUᐒ3�����ND� ADCO�Lp%� {.CMNT�/ �%� �����.E#>!�/4�%P�OSCF�'�.PgRPM�/9ST� {1��� 4@��<#�
1�5�? �7{?�?�?�?�?�?�? )OOO_OAOSO�OwO��O�O�O�O_�A�!S�ING_CHK � �/$MODA�Q,#����.;UD�EV 	��	�MC:o\HSIZ�Eᝢ��;UTAS�K %��%$1�23456789� �_�U9WTRIGW 1���l3%%���9o��"ocoFo5#�VY�P�QNe��:SEM_INF 1�3'� `)�AT&FV0E�0po�m)�aE0�V1&A3&B1�&D2&S0&C�1S0=�m)A#TZ�o;"tH?g�a[o�xA��z���� �o>��o '��K����� ��я:�L�3�p� #�5���Y�k�}���� ��$�[�H���~�9� ����Ưد�������� ӟ�V�	�z������� c�Կ����
��.�� �d��)�;��Ͼ�q� ������˿<���`� G߄ߖ�IϺ�m�ϑ� �����8�J��n�!߀��M�������h_N�ITOR� G ?��[   	EOXEC1�/�25�35�45�55��P7�U75�85�9�0� �Қ�4��@��L�� X��d��p��|��P������2��2��U2��2��2��2��U2��2��22�3��3��3@�;QR�_GRP_SV �1��k (�A����??���4[Ͻཌ���q���j]��Q_D��^�PL�_NAME !�3%,�!De�fault Pe�rsonalit�y (from �FD) �RR2�� 1�L6(�L?�,0	l d������ ��//(/:/L/^/ p/�/�/�/�/�/�/�/ZX2u?0?B?T?f?@x?�?�?�?�?\R<? �?�?O O2ODOVOhO�zO�O�O�OZZ`\R�?�N
�O_\TP�O:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHo_)_~o�o�o�o �o�o�o�o 2D Vhz�[omo�� ��
��.�@�R�d��v���������Џ�� Ef  Fb�� F7���  G ��!��d� �@�R�6�t����獀�l���ʝ����� ݘ����"�@� F�d���� "𩯹�ݐA�  ϩU[�$n�B�oE �� �� @D�  �?��� �?�@��A@��;f��FH� ;��	l,�	 �|��j�s�d�>���� ��� K(���Kd$2K ���J7w�K�YJ˷�Ϝ�J�	�ܿ�� @I����_f�@�z���f�γ��N������	X�l������W�S�ĽÔ��I �����5����  ����A?o�i#�;��A��� ���l� �Ϫ�-���ܛG��G�Ѳ��@n��@a   �  ��ܟ*�͵	'� � H��I� �  ��Рn�:�È~l�È=��̈́�в@�ߚЕ�����/�����̷N<P�  ',����-�@
�@�U��?=�@A���?B�  Cj�a��Be�Ci��@#��Bи�� L �,ee��^^ȹBР��P��`��̠�����ADz՟ �n�3��C�i�@�R�pR�Yщ��  �@O� ��Ż���?�ff������n� ɠ#ѱy9�G
(���I�(�@uP@~����t�t���>�����;�Cd;���.<߈<�g�<F+<L�������,�d�,�̠�?fff?��?&�&��@��@x���@�N�@�?��@T�H�� ��!-�ȹ�|�� 
`�������/ /</'/`/r/]/�/��eF���/�/�/�/@m?��/J?�(E���G�#�� F Y�T?�?P?�?�?�?�? �?O�?/OO?OeOk� ��O�IQOG�?�O1?��OmO_0_B_T_������A_�_	_�_P�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�ol�o���W�����o;C�E� q�H�d��؜a@q��e��F�BµWB]��NB2�(A����@�u\?��D�������b�0��|�uR�����
x~�ؽ���Bu*C���$�)`�$ ����GC#����rAU�����1�eG��D�I�mH��� I:�I��6[F���C��I��J�:�\IT�H
~�QF�y��p���*J�/ I8�Y�I��KFjʻCe�o��s��� ��Џ���ߏ�*�� N�9�r�]��������� ���۟���8�#�\� G�����}�����گů ���"���X�C�|� g�����Ŀ������ �	�B�-�f�Qϊ�u� ���ϫ��������,� �P�b�M߆�qߪߕ� �߹�������(��L� 7�p�[����������s($���3:�����$���3���d�,�4��x@�R��񴲚�l�<~�wa���e����wa4 �{����@��(L:ueP�	P~�A�O�������	���� G2W}h� �����/�� �O�O7/m/[(d=�s/ U/�/�/�/�/�/?�/�1??U?C?y?�=  �2 Ef9gFb-��77�9fB)aa�)`C9A`�&`w`@ -o�?9de�O-OOQOpn�?�?�O�O�O�O�9c?�0�A7ht4Rw`w`!w`xn
 �O9_K_]_o_ �_�_�_�_�_�_�_�_po#ozzQ ��h���G���$MR�_CABLE 2}�h �a:�T� @@�0�A�e��a�a�a��`���0�`C�`�aO8��tB����bo}GT D�D�F��o�f�#��0���0�DO���`����0��CbD�%���o�h8  ����C�07�d�4�`���P�}�T D��R"�4��`y`By`C\�p�bHE��`�,�w��И5D��#z�lҠ`��0�q�pήb0��abr3E}�T D�R��y /o�c-���H� �2��� V�����������'��"���D���^q��o <�\���������������*,�**} \cOM �ii�����h2���q%% 2345?678901i�{�! f�����������15����
��`��not se�nt 5���;��TESTFE�CSALGupeg�`��1d.�š
:�� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.x�ml��ֿ�`Z��DEFAULT�-��4\bGRP 2�M�  =�U[�  �%For�ce�sor c?heck  ������z��p����h5-���ϻ��������%�!1st cle�aning of� cont. v��ilation��}�Rߗ+��[��Дߦ߸���me;ch�cal`������0��h5k�@�R�d�v����>(�rolle_Ƶ����/���(��:�L��Basi�c quarte�rly�������,�������������M��:(�"GpP(�X_h5�������#C���M"��{Pbt�|��Suppq�greasq� ��?/&/8/J/�\/��C+ ge��./ batn�y`/��/h5	/�/�/�/?� ?_�ѷen'�v��/�/��/��?�?0�?�?�?�G=?O��ap"CrB1O��0 �/`OrO�O�O�O�t$,��Lf��C-(��A�O:�OO$_6_H_Z_�l_�t*cabl,�O(���S<(��Q�_:�
_�_�_oo�0oo)(Ӂ/�_�_����_�o�o�o�o�o��O@hau1�l�2r x(�<qC:��op������_ReplaW�fU��2�:�._4�F�X�j�|�(�$%���ߟ ����#���
��.�@� ��d���ŏ׏����П ����U�*�y����� r���������	�q�� ?�߯c�8�J�\�n��� ϯ�����ڿ)���� "�4�Fϕ�jϹ�˿�� ����������[�0� ϑ�fߵϊߜ߮��� ��!���E�W�,�{�P� b�t����߼��� ��A��(�:�L�^��� ������������  $s�H������q �����9] o�Vhz��� U�#�G/./@/ R/d/��/�/��// �/�/??*?y/N?�/ �/�?�/�?�?�?�?�? ??Oc?u?JO�?nO�O��O�O�O+Jkb	 H �O�O__6M2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o�*<ND@ ̾bA?�  @!Q _���Fwp�� �H* �** @A>F�pRT��f�x�:�������ҏ��eO^C7�Տ#�5� G�	�k�}���ُ��� c�����W��C�U� g���ß)�����ӯ� ��	��-�w�����9� ������m�Ͽ��=��O�E!Q�$MR�_HIST 2��>EN�� 
 \�
B$ 2345678901^�f�#�
�]�9O���φ� ��O�)�;����q� �ߕ�L�^߬����ߦ� ���7�I� �m�$�� ��Z���~������!� ��E�W��{�2������h�����:�SKCF�MAP  >EKQ��r5�!P�����ONREL7  .�3����EXCFENB�8
��QFNC�XJJOGOVL�IM8dNá ��K�EY8��_�PAN7����R�UN����SFSPDTYPx<C��SIGN8J�T1MOT�G���_CE_GRP7 1�>EV� �@�����/Ⱥ ��/�/U//y/ 0/n/�/f/�/�/�/	? �/???�/c??\?�? P?�?�?�?�?�?O)O�OMO,���QZ_E�DIT5 )TC�OM_CFG 1����[�O�O�O }
�ASI �yB3�
__+[_�O_��>O�_bHT__ARC_U.���	T_MN_MO�DE5�	UA�P_CPL�_gN�OCHECK ?��� ��  o.o@oRodovo�o�o �o�o�o�o�o*�!NO_WAITc_L4~GiNT�A����EUwT_E�RRs2���3��@ƱJ�����>_�)��|MO�s��}x�:E�~$�A��	�������Z§�C	~��E�8�?��4���4� �~�rPA�RAM�r�����s_��5�5�G� = ��d�v�~�X� �����������֟�0����b�t������SUM_RSPACE�����Aѯۤ��$ODRDSP��S7cOFFSET_CARt@�_��DIS��PEN_FILE:�7�A�F�PTION_�IO��q�M_P�RG %��%$�*����M�WORK� �yf C��춍���  '� �������G	 ������It���RG_DS�BL  ��C��{u��RIENTkTO7 �C� �A �UT_S/IM_Dy����V�LCT ���}{B �٭��_P�EX�P=��RAT��W dc��UOP ���`����e�w�]ߛߩ��$��2r�L6(�L?���	l d������&�8� J�\�n������� �������"�4�F�X���2�߈���������@����*�<w� Tfx��������J` [ˣG���Tz��Pg������ /"/4/F/X/j/|/�/ �/�/���/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?�/�/,O>O PObOtO�O�O�O�O�O �O�O__(_:_��O���y_�]2ӆ� �_�^�_�_�W^]^]��/ooSog��Hgro hozo�o�o�o�o�oF`��#|G`A� � 9y����OK�1��k������<�E�A�nq @D�C  �q����nq?���C��s�q1� ;��	l��	 �|�Q�s�r�q>���u
��qF`H<�zH~�H3�k7GL�zH?pG�99l7�0k_B�T�F`C4��k��H���t��-�Ae����k�����~s���  �ሏ�����EeBVT����dZ=���ڏ ���q�-�Fk�y�{FbU��= n@6�  ���z�Fo���Be	'� � ���I� � � �:p܋=��q�ڟ웆�@�@��B�,���B����g�AgN����  '�|���g��B��
p�BӀC׏����@?  #�Bu�&��ee�^^މB:p2���>�m�06p�Z�=Dz?o}� ܏������׿�������Ǒ��� f�  ȧ �M���*�?��ff�_8�J�ܿ !3pϑ�ñ8= �ϐ�ʖq.·�(= ��P@���'��s�tL�>���/�;�Cd;���.<߈<�g�<F+<L ��^oiΚrd@��r6p�?fff?�?&��п�@��@x���@�N�@�?��@T싶�Z ���ћtމ�u�߈w	� x��ti�>�)�b�M�� q����������� ��:�%�^�������W����S�E�  G}�=F�� Fk� ��������1U@ yd������q ��	��{�A��h@�����a��ird��A{/w/J/(5/n/	�A��A���":t�/ C^/�/Z/ ލ?���/�/1?,?���W����g��pE� ~1�?0�4�0
1�1@I�Ӏ��BµWB]��NB2�(A���@�u\?����������b��0�|�uR�����
�>�ؽ���Bu*C��$�)`�?� ���GC#����rAU�����1�e�G���I�mH��� I:�I��6[F���C�4OI��J��:\IT�H
?~QF�y�Ol@��*J�/ I�8Y�I��KFjʻC��-?�O�O __>_)_b_M_�_�_ �_�_�_�_�_o�_(o o%o^oIo�omo�o�o �o�o�o �o$H 3lW�{��� ����2��V�h� S���w�����ԏ���� ���.��R�=�v�a� ������П����ߟ� �<�'�`�K�]����� ����ޯɯ��&�8��#�\��3(J���3�:a������J�3Ï�c4�����������������xڿ�n����e�<�n�4 �{2�2ɀr�`ϖτϺϨ��%PR�P���!�h��!�K�6�o�Z�����u�|ߵߠ������� ���3��W�B�{�f�@4���������d�A ����!��1�3�E�{��i������������� � 2 Ef�7F[b�7��6B�!,�!� C9� �� n�@�/`r������#x��+D=�3?, V�8v�n�n��n��.
 D��� ��//%/7/I/[/�m//�/�:� ���ֻ�G���$P�ARAM_MEN�U ?2���  �DEFPULSE��+	WAITT�MOUT�+RC�V? SHE�LL_WRK.$�CUR_STYLv� 4<OPTJNJ?PTB_?Y2C/?R_DECSN 0 �Ű<�?�?�?�?�?O O?O:OLO^O�O�O�O��O�O�!SSREL?_ID  .�����EUSE_PR_OG %�*%�O0_�CCCR0�B���#CW_HOST !�*!HT�_=ZAT��O_�Sh_zQ�S|�_<[_TIME
2��FXU� GDEB�UG�@�+�CGINP_FLMSKo�5iTRDo5gPGA�b` %l�tkCH�Co4hTYPE�,� �O�O�o#0 Bkfx���� �����C�>�P� b���������ӏΏ�� ���(�:�c�^�p������7eWORD �?	�+
 	�RSc`n�PNS2��C4�JOv1���TE�P�CO�L�է�2��gLP �3��n��OjTR�ACECTL 1�2��! .��m n����|��q�DT Q�2��Ǡ��D � _: Ԡؤؤ��ڢׯ� ����1�C�U�g�y����������ӿ���':�����X}`���1�<���&�@.�K�uJ�qJ�H�EH�	H�?�K�H�UH�H�H�H�T�@J�H�H�H��E�W�i�{ύϟϰ�������;��a�ߞ߰����� ���'��������� ������'���/��� 7���?���G�3�ݿ� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������С �*<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6@ubt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀�V�߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z?��?�?�?�?�1�$P�GTRACELE�N  �1  ����0���6_UP �����A@�1�@�1_CFG ��E�3�1

@�<D�3UOaHSO��0$BDEFSPD� �/L�1�0���0H_CONF�IG �E�3� �0�0d�D�&�2 �1�APpDsAl�A�0��0IN'@?TRL �/MOA�8pEQPE�E��G�A<D�AIWLID(C�/M	bT�GRP 1ýI� l�1B � �����1A��33FC� F8� E�� @eN	�A�AsA�Y�Y�A�@?� 	 vO�Fg�_ ´8cokB;`baBo,o>oxobo��o�1>о�?B�/�o�o~�o =%<��
 C@yd��"�������  Dz@�I�@A0�q� � ������ˏ���ڏ� ��7�"�4�m�X���|����Ú)ґ
V7�.10beta1�HF @�����Aq��Q�  �?� �B���P�p �C��~&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@p���f������ҡr�R�ܣ�Rљ����1�i�������t<B!CeQKNO?W_M  lE7F�bTSV ĽJ�BoC_�b�t��������������1�]aSM��SŽK ���	�NB�0����ĿK���-�bb��A�RP���`�0�Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1=�K
 4MU�iǨj� K�]�oߠ� �ߥ߷�������2�� #�h�G�Y��}������
������,�2r7�I��1�<t�H��P3^�p�����,�A4��������,�5(:,�6Wi{�,�7����,��8�!3,�MA�D�6 F,�OV_LD  KD��xO.�PARNUM�  ��C/%�S+CH� E
9'!8G)�3Y%UPD/���E�/P�_CMP_0��0@�0'7E�$�ER_CHK�%05H�&�/�+RS����bQ_MO�+?=5_�'?O�_RES_G6��:�I�o�?�?�? �?O�?O7O*O[ONO OrO�O�O�{4]��<�?�Oz5���O__ |3 #_B_G_|3V b_ �_�_|3� �_�_�_|3 � �_�_o|3Oo>o<Co|2V 1�:�k1�!�@c?�=2T?HR_INRc0i!�}�o5d�fMASS6�o Z�gMN�o�c�MON_QUEUE �:�"�j0��Ut4N� U1Nv�+DpENDFqd?`y�EXEo`u� BE�npPAsOPTIO�Mwm;DpPROGR�AM %$z%�Cp}o(/BrTASK�_I��~OCFG� �$��K�D�ATA��T���j12,ź�̏ޏ�� ���&�8�J�\�n���������ȟ{�INFO�͘��3t��!� 3�E�W�i�{������� ïկ�����/�A�@S�e�w�����Θ�a '��FJ�a K_N���T��˶ENB�g ڽw1��2��G�N�2�ڻ P(O�=���]�ϸ�@���v� ��u�uɡdƷ_E?DIT �T���|��G�WERFL�x��c)�RGADJ {Ҷ�A�  $Ձ?j00��a�Dqձ���5�?�D�ʨ�<u�j0�%e`������FӨ�2�R�V�	H;pl�G�b�_�>�pAod�t$��*�/� **:�j0�$�@킆5Y�T���^��q �߈b~�L��\�n�� ������������ ��4�F�t�j�|����� ��������bL BT�x���� :��$,�P b���/��� �/~/(/:/h/^/p/ �/�/�/�/�/�/V? ? ?@?6?H?�?l?~?�? �?�?.O�?�?OO O �ODOVO�OzO�O_�O �O�O�O�Or__._\_ R_d_�_�_�_�_�_�_�f	g�io�pWo�o{d �o�~o�ozo�B�PREF ��Rږp�p
�IOORITY�w[���MPDSP�q��pw�UT6����ODU[CT3���v��OG��_TG���8��ʯrTOENT� 1׶� (!AF_INE�p�,�7�!tcp|7�_�!udN�~��!icmv���ޯrXYK�ض���q)� ,�����p��&�	��R� 9�v�]�o�����П�������*��N�`�*�sK��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b��t����u�w�HANCE �R��:�Bwd��连�2s�9�Ks��PORT_WNUM�s�p����_CARTR�EP{p�Ω�SKS�TA�w d�LGmS)�ݶ��t���pUnothing�������{��TEMP ޾y���'e��_a_seiban�o\��o lߒ�}߶ߡ������� ��"���X�C�|�g� ������������� 	�B�-�f�Q���u��� ����������, <bM�q��� ����(LٟVERSIyp�w�} disa�bledWSAV�E ߾z	2600H768S	?�!ؿ�����/ 	5(�r)og+^/y�e{/�/�/�/�/"�*�,/? �p����_�p 1�Ћ�� ������Wh?z?�W*pURG�E��B�p}vgu,�W�F�0DO�vƲ�vW�%��4(�C�WRUP�_DELAY ��\κ5R_HOT %Nf�q׿GO�5�R_NORMAL�&H�r6O�OZGSEM�IjO�O�O(qQSKKIPF3��W3x= _98_J_\_]�_�_ {_�_�_�_�_�_�_	o /oAoSoowoeo�o�o �o�o�o�o�o+= aOq���� ����'��7�]��K�������)E�$R�A{���K/�zĀ~Á_PARAM�A�3��K @.�s@`�61�2C<�5�y��C�6$�=BÀBTIF�4`�RCVTMOUu��c��ÀDCR�F3��I ��+QB�s�D��ߚD�J:��ϗ9±"Z¹{�ޅ��_�1��J��_��k_ �;�Cd;���.<߈<�g��<F+<L�A��Ѱ��d�u�L� ������ϯ�����)�;�M�_���RDI�O_TYPE  �M=U�k�EFPO�S1 1�\�
 x4/�œS����0� )/T��x��uϮ�I� ��m��ϑ�ߵ����� �t�_ߘ�3߼�W��� {�����:���^��� ���/�A�{����� � ��$���H���E�~�� ��=���a������������D/h��S2 1�KԿX��T�x��3 1� ����nY�S4 1�'9K��/�'/�S5 1���/�/�/|�/:/S6 1�Q/�c/u/�/-??Q?�/S7 1��/�/
?D?��?�?�?d?S8 1�{?�?�?�?WOBO{O��?SMASK 1�L��O�D�GXN�O���F&�^��MOCTEZ�Ż��Q_ǁ��%]pA݂��PL_RANG!Q]�_QOWER �ŵ��P1VSM_DRYPRG %ź�%"O�_�UTART� �^�ZUME_PRO�_�_4o���_EXEC_EN�B  J�e�GS�PD`O`WhՅjbT3DBro�jRM�o�h�INGVERSI�ON Ź�#o�)I_AIRPURhP �O(�M�MT_�@T�P#_�ÀOBOT_ISOLC�NTVő'q�huNAME�l���o�JOB_ORD_NUM ?�X�#qH76�8  j1Zc@n�r
�rV�sw��r�?�r�?�r�pÀPC�_TIMEu�a�x�ÀS232>R1��� LTE�ACH PENDcANw�:GX��!O Maint�enance C�onsj2����"���No UseB�׏������1�8C�y�V�NPO�P@��YQ�cS�C7H_L`�%^ ��	ő��!UD�1:럒�R�@VA#IL�q@�Ӏ�J�Q�SPACE1 2�ż ��YRs�i�@Ct�YRԀ'{��?8�?��˯ ����"���7�2�c� u�����G���߯ѿ� ���(��u�AC�c� u�����Ͻ�߿���� ���(��=�_�qσ� ��C߹������߱�� $��9�[�m�ߑߣ� Q������߭��� ��� 	�W�i�{���M��� ����5���.S� e�w�����I����� ��*?as ��E����� /&//;/]o�� ����/2/�/?"? �/7?Y/k/}/�/�/O? �/�/�?�?�?O0OO~KA��*SYPp�M*�8.302�61 yB5/21�/2018 A� �WPfG|�H�_�TX`� !$C�OMME��$USAp �$ENABLED�Ԁ$INN`QpI�OR�B�@RY�E_�SIGN_�`�AP��AIT�C�BWRKz�BD<�_TYP�CRINDXS�@W��@%VFRI{�_G�RPԀ$UFR�AM�rSRTOOL�\VMYHOL�A�$LENGTH_�VTEBTIRST��T  $SE�CLP�XUFINV�_POS�@$�MARGI�A$�WAIT�`�ZX2l�\�VG2�GG1�AAI�@�S�Q	g�`_WR��BNO_USE_�DI�BuQ_REQ��BC�C]S$CUR_TCQP�R"a^f� �GP_STA�TUS�A @ ��A3`�BLk�H$�zc1�h�P@���@_��FX �@E_MLT_CT�C�H_�J�`CO�@O�L�E�CGQQ$W��@w�b#tDEA�DLOCKuDELAY_CNT�a�3qGt�a$wf �2 R1[1T$X<�2[2�{3[3$Zwy�q%Y�y�q%V0�@�c�@�b$V�`�R�V�UV3oh>b�@� � �d�0arMSKJ�LgWaZ�C`�NRK�PS_RATE�0$���S
`�Qv�TAC��PRD��$�e�S*��a4�A�0:�DG�A 0�P�f�lp bquS2�ppI�#`
`�P 
��S\`  ؾA�R_ENBQ ��$RUNN�ER_AXI�<`A�LPL�Q�RU�THI�CQ$FLIP�7��DTFEREN|��R�IF_CHS�U�IW��%V)�G1�����$PřA�Q�Pnݖ_JF�PR_P��	�RV_DA�TA�A  =$�ETIM���_$VALU$�	��OP_   ��A  2 ��SC*�	�� �$ITP_0!�SQ]PNPOU}�o��TOTL�o�DSP>��JOGLIb��P'E_PKpc�Of�i���PX]PTAS��$KEPT_MI�R��¤"`M�b�A	Pq�aE�@�y�q��g@١c�q�PG�BCRK6�x���L�I��  ?�SJ�q�P��ADEz�ܠBSO�Cz�MOTNv�D�UMMY16Ӂ�$SV�`DE_O�P��SFSPD_�OVR
���@L�D����OR��TP8�LE��F������OV��SF��F����bF�d�ƣ&c)�fQ~c�LCHDLY��RECOV���`���W�PM��gŢ�ROȲ�����_F�?� �@v�S �NVER\�@�`OFS�PC,�CSWDٱc�ձ���B,����TRG�š�`�E_FDO��MB�_CM}���B��BALQ�¢	�Q�̄VzaF�BUP�g��G
��AM���@`KՊ�fe�_M!�d�AMf�<Q��T$CA����uDF���HBKd��v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�Dd�9�1A��9�3A�^��ATIO�0���͠��US����WaAB��R+c�`tá`Dؼ�A��_AUXw�S�UBCPUP���S �`����3Եжc����3�FLA�B�HW�_Cwp"�Ns&�]sA�a��$UNIT�S�M�F�ATTR�Iz�Z�CYCL��CNECA���F�LTR_2_FI~��TARTUPJp0����A��LP����ޖ�_SCT*cF_�F�F_P���b�FS8��+�K�CHA/Q��p*�d�RSD��`Q����Q���_TH��PROr���հEM�PJ���G�T�c �Q�DI�@~y�RAILAC/��bMX�LOf�xS���ځ���拁���P�R#�S`app�C�� 	��FUsNC���RIN``QQP� ԱRA)]R ��AƠ��AgWAR֓��BLZa�WrAkg�ngD�AQ�B�rkLD@�र&q�M�K����TI���j���$�@RIA_SWV��AF��Pñ#���%%�p9r1��MO9IQ���DF_~P(��PD"LM-�FA��PHRDY�DORG�H; _QP�s%MULSE~Pz���**�� J��Jײ���FAN_ALMsLVG��!WRN�%�HARDP��UcO��� K2$SHADOW]�kp�a02��N� STOf�+�_^�w�AU{`R��eP_SBR�z5���:�F�� �3MPIN�F?�\�4��3R3EGV/1DG�+c1Vm �C�CFL(��?�DAiP���Z`Ɨ� �����Z�	 ��P(Q$�A$�Z�Q V�@�[�
7� ��EG��o����kAAR���㌵2p�axG��AXE��wROB��RED���W�QD�_�Mh�SY�A��AF��FS�GWRqI�P~F&�STR��(��E�˰EH�)��D�a\2kPB6P��=V���Dv�OTO�1)���ARYL�tR��v�3���FI&�ͣ$LINKb!\��Q%�_3S���E�N�QXYZ2�Z5�V'OFF���R�R�X%xPB��ds�G�cFI�03g�h������_J���'�ɲ�S&qR0LTV[6����aTBja�"�bCL���DU�F7�TUR� X��e�Qb�2XP�ЊgFL�@E���x@�`�U9Z8��^�� 1	)�K��	Mw��F9��劂����ORQj��G;W3���#�Ґd ���upz����1�tOVE�q_�M��ё?C�uEC�u KB�v'0�x-�wH��t ���& `��qڠ� B�ё�u�q�wh�ECh�L���ER��K	�!EP����AT�K�6e9e�W���AXs�'��v�/�R  ����!�� ��P ��`��`�3p�Yp�1�p�� �� � � (�� 8�� H�� X� � h�� x�� ������oDEBU�$`%3�I��·RAB�ȱ�ٱ�sV��� 
d�J、��@񘧕� ������Q���a���a ��3q��Yq+$�`%"<�.cLAB0b�u��'�GRO���b<��B_s��"Tҳ*`��0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθu�ݸ��PNT0����SERVE �Z@� $`EAV�!�PO����nP!��P@�$!Y@ w $>�TRQ�b�
=��BG�K�%"2�\��� _ � l��5�D6ERRVb(�I��V0`;���'TOQ:�7�L�@
�(R��e G�%�Q��q <�50F� ,��`�z�>�RA� �2 d!�����S�  M��px�U ����OCuG��  ��COU�NT6Q��FZN_wCFGF� 4#��6��TG4�_�=������Î�VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@HE�L�0�� }5b`B_BAS��RSR�6�CSHH����1�Ǌ�2��U3��4��5��6���7��8��}�ROO0����P�PNLEA�c�AB)ë ��ACK�u�INO�T��(B$�UR0� =�_PUX��!0��OU+�Pd��8j��� V��TPFWD_KAR��L� ��RE(ĉ P�Pܺ>QUE�:RO �p�`r0P1I� x��j�P�f��6�QSE�M��0��� A��S�TYL�SO j�D�IX�&�����S!_�TMCMANRQ܉�PENDIt$�KEYSWITCaH���kHE�`�BEATM83PE�{@LE��>]��Uү�F��SpDO/_HOM# O�@�EF�pPRaB�A#PY�C� O�!��яOV_M|b<0 I�OCM�dFQk��h�HKYA DH�Q�7��UF2��M�x��p�cFORC�3gWAR�"�OM|@  @S�#o0UU)SP�@1�2&�3&4E���T�O���L���8UN�LOv�D4K$ED�U1  �SY�HwDDNF� M��BLOB  p��SNPX_AS�� 0@�0��81�$SIZ�1$�VA{���MULTKIP-��# A� � $���� /4`�BS��0�C<���&FRIFBO�aS���3� NF�ODBUP߰�%@3�;9(��ҋ�Z@ x6��SI��TEs�r.�cSGL�1T�Rp�&�Н3B��@�0ST�MTq�3Pg@VByW�p�4SHOW�5n@�SV��_G��; 3p$PCJ�PЬ����FB�PHS�P AW�EP@VD|�0WC� ���A00��PB XG �XG XG$ XG5VI6�VI7VI8VI9VIAVIBVI�XG�YF�0BXGFVH��XbI1oIU1|I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1YU1Y2UI2bI2oI2|I2�I2�I�`�XP�I2p�X�I2�I2�IU2�I2�I2Y2Y��p�hbI3oI3|I3��I3�I3�I3�I3��I3�I3�I3�I3��I3�I3Y3Y4��i4bI4oI4|I4��I4�I4�I4�I4��I4�I4�I4�I4��I4�I4Y4Y5��i5bI5oI5|I5��I5�I5�I5�I5��I5�I5�I5�I5��I5�I5Y5Y6��i6bI6oI6|I6��I6�I6�I6�I6��I6�I6�I6�I6��I6�I6Y6Y7��i7bI7oI7|I7��I7�I7�I7�I7��I7�I7�I7�I7��I7�I7Y7TiցVP� UD��y"ՠ��
<A62��t�R��CMD� ��M5�Rv�]��Q_h�R���e�����<�YSL���  � �%\2��+4��'��W�BVA�LU��b��'���F�H�ID_L���H�I��I���LE_���㴦�$0C�S�AC�! h ��VE_BLCK���1%�D_CPU5ɧ 5ɛ ������C�� ��R " � PWj��#06��LA�1SBћ������RUN_FLG�Ś����ĳ ����������H���ХĽZ�TBC2��#/ � @ B��e ��S�8=�FTD	C����V���3dՆQ�THF�����R��L�ESERVE9��F��3�2�E�|�Н�X -$��LEN9��F��f�cRA��W"G�W_5��b�1��д2�MO$-�T%S60U�Ik�0�`ܱF����[�DEk�21LACEi0�CqCS#0�� _MA� pj��z��TCV����z�T�������.B i�'A�z�'AJh�#E�M5���J��@@i�V�z���2Q �0&@�o�h��JK��VK�9��{���щ�J0l����JJ��JJ��AAL���������e4��5�ӕ N1��P����.�LD�_�1�* �CF�"%{ `�GROU��(�1�AN4�C�#m ?REQUIR���EBU�#��6�$Tk�2$���z�܏ #�& \�AP�PR� C� 0�
$�OPEN�CLO�S�St��	i�
\��&' �Mf�p����W"-_MG�7CB@�A���B�BRK@NOLD|@�0RTMO_5�H�p1J��P�� ������������6��1�@ �)!�#�(� ������'��+#PATH''@!6#@!��<#� � '��1SCaA���6IN�ңUCJ�[1� C0@UM�(Y ��#�"������*���*��� PAYwLOA~J2LؠOR_AN^�3L���91�)1AR_F�2LSHg2B4LO�4�!F7�#T7�#ACRL_�%�0�'�$r��H��.�$HA^�2FLEX��J!�) P�2�D��߽���0��* :����z�FG]D��`��z���%�F1]A �E�G4�F�X�j�|���BE���������� ��(��X�T*�A���@�XI�[�m�\At�T$g�QX<�=��2TX ���emX���������� ��������+	�J>+ �-�K]o|�٠AT�F�4�CELFPѪs�J� �*� JEmCTR��!�ATN�vzH�AND_VB.���1��$, $8`Fi2Av���SW��
"-� $$M*0.�]W�lg��PZ����A��� 1�����:AK��]A�kAz��LN�]D*kDzPZ G��C�CST_K�lK�N}DY��� A����0 ��<7]A<7W1�'��d�@g`�P����0���" 1B$. M�2D%"��H�<���ASYMj%0�	� j&-��-W1�/_�{8� �$���� �/�/�/�/ 3J<��:9�/�89�D_VI��v����V_UCNI�ӛ��cD1J�� ��╴�W<��n5Ŵ� w=4��9��?�?<�ucI�4�3P�%�H����/�j��0�D)IzuO��L�k�N>0 �`��I��A��#���@ģ���@���IPl� 1 �� /�ME.Q�p��9�ơT}�PT@�;pG �+ Gt� ����'��T�0� $DUMMY}1��$PS_�@�RF�@;�$b�n'FLA@ YP(c�|��$GLB_TP�ŗ���9 P�q��2 X� z!�ST9�� SBR�M M21_V�T�$SV_ER*0O��p����CL����A�GPO��f�GL~�E�W>�3 4H �+$YrZrW@�x��A1+�A���";�"�U.&�4 8`NZ�"��$GI�p}$�&� -� �Y�>�5� LH {��}$Fz�E��NEAR(P�N�CF��%PTAN9C�B;�JOG�@�� 69�$JO�INTwa?pd�MS�ET>�7  x�E��HQtpS{r��up>�_8� �pU.Q�?�� LOCK_�FOV06���BGL�V�sGLt�TES�T_XM� 3�EM�P�����_�c$U&@%�w`24� �Y��5��2�d��3���CE- ���� $�KAR�QM��TP�DRA)�����VE�Cn@��IU��6���HEf�TOOL��C2V�DRE I�S3ER6��@ASCH� 7?Ox L�Q�29Z�H I��  @$RAI�L_BOXEwa��ROBO��?�~�HOWWAR�1x�_�zROLMj� �:qw�jq� �@ �O_Fkp! �  �l>�9�� +�R O8B: �@��c�OU�;��Һ�3ơ�r�q_�/$PIP��N&`H��l�@��#@CO�RDEDd�p >S�f�fpO�� < 7D ��OB⁴s d���Kӕ���qwSYS�ADR�q�f��TCHt� 7= ,8`ENo��1Ak�_{�-$Cq7��f�VWVA��>� �  &��P�REV_RT��$EDITr&VSHWRkq�֑ &RJ:�v�D��JA�$~�a$HEAD�h6�� �z#KE:�E�CPSPD�&JKMP�L~�R*PF��?��1%&I��5S�rC�pNE; �q��wTICK�C��M��1��5HN��@� @� 1Gu�!_GqPp6��0STY'"xLO��:�2l2?�_A t 
m G3%S%$R!{�=��S�`!$��w`���ճ�r��Pˠp6SQU��x�E��u�TERC�����TSUtB ����hw&`gw�Q)b�pO����@IZ��4{��^�PR�kј�B1XPU���E_�DO��, XS�KN~�AXI�@���UR�pGS�r� ^0�d&��p_) �ET�BQPm��o��0Fo�2�0A|���Rԍl��a<�SR�Cl>@P��b_� yUr��Y��yU��yS�� yS���UЇ�U���U�� �U�]��Ul[��Y�bXk�]Cm������YRSC�� D �h�DS~0��Q�S�P���eATހ���A]0,2N�ADDR�ES<B} SHIyF{s��_2CH�p��I��=q�TV
srI��E"���a�C*T�
��
;�VW�AN��F \��q��0l|\A@�rC�_B"R�{zp�ҩq�TXS�CREE�Gv��1TINA���t�{����A�b?�H T1�ЂB�����I���A��BE�y RRO������� B���1UE4I �g�!p�9S��RSM]0�GUNEX(@~Ƴ�j�S_S�ӆ��Á։�ģ��ACY�0� [2H�pUE;�J�¸���@GMT��L�ֱ�A��O	�BB�L_| W8���K ���0s�OM��L1E/r��� TO!�s��RIGH��BRD<
�%qCKGR8л��TEX�@����WIDTH�� �B�|�Z<��I_��Hi�� L 8K���_�!=r���R:�_���Yґ��O6q�M�g0紐U��h�Rm��LUMh��FpGERVw��P����`�N��&�GEKUR��FP)�)� �LP��(RE%@�a)�ק�a�!��f �5*�6�7�8Ǣ#B@�É@���tP�fW��S@M�USR�&�O <����U8�Qs�FOC)��PRI;Qm� :����TRIP�m�SUN����Pv��0 ��f%�~Œ����@�0� Q����AG ��0T� �a>q�O	S�%�RPo���8�R/�A�H�L4����U¡�SU�g��8¢5��OFF����T�}�O�� �1R�����S�G�UN��6�B_�SUB?���,�SR	TN�`TUg2��mCsOR| D�RAUrP�E�TZ�#'�VCCܵ�	3V AC3�6MFB1��d�P=G �W (#��ASTEM����䦒0PE��T3G�X� �\ ��MOVEz�A��AN�� ����M���LIM_X ��2��2��7�,���`��ı�
�BVF�` E���~��04Y���IB�7���5S��_�Rp� 2��� WİGp+@��}СP|��3�Zx ���3���A�ݠ9CZ�DRID��B��Vy08�90� De�?MY_UBYd�� �6��@��!��X���P_S��3��L��KBM,�$+0DEY(#EX`�����_UM_MU� X����ȀUS�� ���=G0`PACI���� �@��:��:,�:�����RE/�3qL�+���:[��TAREG��P�r��R<�\ d`��A��$�i	��AR��SW2 $��-��@Oz�%qQA7p�yREU�U�0�1�,�HK�2]g0�qP� N� �sEAM0GWOR����MRCV3�^� ���O�0M�C��s	���|�REF_���x(�+T�  ���������3_RCH4(a�P �І�hrj�NAۑXQ��0�_ ��2����L@4��n�@@OU~7w�6���Z��a2[ư�RE�p�@;0\��c�a'2K�@SUL���]��C��0�^��� NT��L�3��@(6I�(6q�(3� L��@Q5��Q5I�]7q�}�)Tg`4D`�0.`0ПAP_HUC�5S]A��CMPz�F�6(�5�5�0_�aR��a��1I\!X�9��GF}S��ad ��qM��0p�UF_x�0�B� �ʼ,RO��Q���'����UR�3GR�`.�3IDp���)�D�;��A��~�IEN��H{D���V@A J���S͓UWm�i=�����TYLO�*�5����b�t +�cPA�= �cCACH�vR��UvQ��Y��p�#CZF�I0sFR�XT����Vn+$HO��� �P!A3�XBf�(1 ���$�`VPy� ^bO_SZ313he6K3he12J�eh chG�6chWA�UMP�j���IMG9uPAD<�iiIMRE�$�b/_SIZ�$P�����0 ��ASYNBU=F��VRTD)u5t�qΓOLE_2DPJ�Qu5R��C��U���vPQuECCUlVEMV �U�r�W�VIRC�aIuVTPG���rv1s��5qFMPLAqa��v�V�0�c��� CKL�AS�	�Q�"��dC  �ѧ%ӑӠ@}���$�Q���Ue | �0!�rSr�T�#0! �r�iI��m�v6K�BG��VE�Z��PK= �v�Q�&�_�HO�0��f � �>֦3�@Sp�SL�OW>�RO��A�CCE���!� 9�V�R�#���p:���AD�����PAV�j�� uD����M_B"����^�JMPG ��g|:�#E$SSC�� F�vPq��hݲvQ�S�`qVN��LEXc�i T`�sӂ��Q�FLD �DEsFI�3�02����:��VP2�VjO� �A��V�4>[`MV_PIs���t���A�@��FI��|�Z��Ȥ�����A0���A��~�GAߥ1 �LOO��1 JCB����Xc��^`�#PLCANE��R��1F�c �����pr�M� [`�噴��S����f�����Af��R�Aw�״t�U��pRKE��d�V�ANC�A���� �k���ϲ�R;_AA� l��2�� ��p�#|"�m h�@��O K�$������kЍ0OU&A�"A��
p�pSK�TM�@FVIEM 2l ���P=���n <�<��dK�UMMYRK1P��`D倛�ACU��#AUކ�o $��TI}T�$PR�����OP���VS�HIF�r�p�`J�Qsԙ�fOxE-$� _R�`U�#�� ��s��q������G�"G�޵'�T�$�SsCO{D7�CNTQ  i�l�>a�-�a�;�a�H�a�V���1�+�2�u1��D���� � 5��MO�Uq���a�JQ������a_�R[�r�n��*@LIQ�AA/`�XKVR��s�n�TL�ޡ�ZABC�tВt�c�
AZIeP��u���LVbc�Ln"���MPC5Fx�v:�$�� ����DMY_LN��������@y�w �p�(a�u� MCM�@}CbcCART_��DPN� $	J71D��=NGpg0Sg0�BUXW� >��UXEUL|ByX���	���|!Z��x P	���m�YH�Db  y 80���0�EIGH�3n�?(�� H����$z a���|�����$B� �Kd'��_��L3�R�VS�F`���OVC�2'�$|�>P&���
q���5D�T�R�@ �V�1�SP9HX��!{ ,� �*<�$R�B2 �2 ���C!��  �@V+| b*c%g!(H�b)g"�`V*�,?8�?�V+�/ V.�/�/?�/�/V(7%3@/R/d/v/�/6?�/ �/�?�?�?O4OOION;4]?o?�?�?�?SO �?�?�O_�O0_Q_8_f_N;5zO�O�O�O�O p_�O_o8o�_MonoUo�oN;6�_�_�_�_ �_�oo%o4Uj�r�N;7�o�o�o �o�o� BQ�r�5� ��������N;8�� ���Ǐ=�_�n����R���ş��ڟN;G ;� џ�
������W�i� {�������ï�.��@�����A��dW� <�N�|�������Ŀֿ �ޯ���0�B�_� R�d�꿤϶������� ������*�L�^�� rτ�
������������&�8�J�l�~�; `ҟ @�з�@���ߩ��-��� �&�,���9�{��� ��a������������� ��A'Y�� �������a#1�
��N;�_MODE  ���S ��[�Y�B���
/\/�*	|/�/R4CWO�RK_AD�	�{#T1R  ����� �/� _INOTVAL�+$���R_OPTION�6 �q@V_�DATA_GRPg 27���D��P�/~?�/�?�9��? �?�?�?OO;O)OKO MO_O�O�O�O�O�O�O _�O_7_%_[_I__ m_�_�_�_�_�_�_�_ !ooEo3oioWoyo�o �o�o�o�o�o�o /eS�w�� �����+��O� =�s�a�������͏�� �ߏ��9�'�I�o��]�����$SAF�_DO_PULS�� �~������CAN_TIM�����ΑR ��Ƙ��5�;#U!P"�Z���� �?E�W�i�{� ����.�ïկ������'(~�T"2�F���dR�I�Y��2�o+@a얿�����)�u��� k0ϴ��_ ��  T�� � �2�D�)�T D��Q�zόϞ� ����������
��.� @�R�d�v߈ߚ�/V�������������B�;�o� �W�p��
�t��Diz$� �?0 � �T"%! ��������� ��������*�<�N� `�r������������� ��&8J\n ��������@"4FX ��� �������� /`4�=/O/a/s/�/ �/�/�/�/�/�!!/ �0޲k�ݵu�0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ ok$o 6oHoZolo~o�o�o�o �o1/�o�o 2D Vhz�/5?��� �����&�8�J� \�n���������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ���`Ò�ϯ� ���)�;�M�_�q� ��������˿ݿ� �����3� ����&2,��	12�345678v��h!B!��*2�Ch���0�� �����������!�3� 9ѻ�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�h�K߰����� ����
��.�@�R�d� v�������������� *<N`r� ������ &��J\n��� �����/"/4/ F/X/j/|/;�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�/ �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_�?L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o=_�o�o �o�o�o�o 2D Vhz�����h������u�o.��@�R���Cz  �B��   ����2&� � �_�
���  	�_�2�Տ�����_�p������ ďi�{�������ß՟ �����/�A�S�e� w���������N���� ��+�=�O�a�s��� ������Ϳ߿���'�9�K�_�������<v�_��$SCR�_GRP 1
�� �� t� ��� ���	 ���������� ������_������)��a����&�DE� DW8���l�&��G�CR-35�iA 901234567890��_M-20��8��?CR35 ��:�#
��������������:֦�Ӧ�G�D��&������	���]�o����:����H���>�� ���������&���ݯ:��j����g��,����B�t�����������A����  @��`��@� ( ?�=��Ht�P
���F@ F�` z�y������  �$H��G`s^p��B�� 7��/�0//-/ f/Q/�/u/�/�/�/8�@��P�� 7%?�����"?W?-2?<����]? H�1�?t���7�������?�-4A, �&E@�<�$@G�B-1 3OZOlO-:HA�H�O�O|O P�B(�B�O�O�_��EL_DEFAULT  ����`~SHOTSTR#]�JA7RMIPOWE?RFL  i�/U�YTWFDO$V� /URRVENT? 1����NU� L!DUM�_EIP_-8�j�!AF_INEx#P�_-4!FT�_�->�_;o!��`o ��*o�o!RP?C_MAIN�ojhq�vo�o�cVIS�o�ii��o!TP&pPU�Ydk�!
PMON_POROXYl�VeZ��2r��]f��!�RDM_SRV���Yg�O�!R���k��Xh>���!
��`M��\i���!RLSYNC��-98֏3�!R3OS�_-<�4"���!
CE4pMTC�OM���Vkn�˟!=	��CONS̟�W�l���!��WA'SRC��Vm�c�;!��USBd��XnR���Noӯ����� ��!��E��i�0����WRVICE_K�L ?%�[ (�%SVCPRG1��-:Ƶ2ܿ�˰3�	�˰4,�1�˰5T�Y�˰6|ρ�˰�7�ϩ�˰�����9����ȴf�!�˱ο I�˱��q�˱ϙ�˱ F���˱n���˱��� ˱��9�˱��a�˱� ���7߱��_���� �����)����Q� ���y��'���O� ���w������ ���˰��İd� c������ =(as^��� ���/�/9/$/ ]/H/�/l/�/�/�/�/ �/�/�/#??G?2?k? V?}?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O�O�O�O	_�O�-_��_DEV ��Y�MC:�5Xd�GTGR�P 2SVK ��b�x 	� 
 ,�P5_�_�R�_�_ �_�_�_�_3ooWo>o {o�oto�o�o�o�o�o �o/A�_e� ��������  �=�$�6�s�Z���~� ��͏���H�'�ޏ K�2�o���h�����ɟ ۟���#�5��Y� @�}�d�v���
�ׯ� Я���1��*�g�N� ��r��������̿	� ��?�&�c�u�̯�� PϽ��϶������)� �M�4�q�X�jߧߎ� �߲������%�|�� [���f������ �������3��W�i� P���t���������>� A(eL^ �������  =O6sZ��  ���/�'// K/]/D/�/h/�/�/�/ �/�/�/�/#?5??Y? �N?�?F?�?�?�?�? �?O�?1OCO*OgONO �O�O�O�O�O�O�O�O,_kT �"V		_R_�=_v_a_�_�_�_�[%���_�_�S��� a�Qeo)goIo7o mo[o�o�i�_�oi�o �o�o%'9o �o��o_���� ��!�w�n��G� ����ŏ���׏�O� 4�s���g���w����� �����'��K�՟?� -�c�Q�s��������� �#�����;�)�_� M�o���ׯ������� ݿ��7�%�[ϝ��� ��K�m�Gϵ������ ��3�u�Zߙ�#ߍ�{� �ߟ߱������M�2� q���e�S��w��� ����%�
�I���=�+� a�O���s�������� !���9']K ������q�m� �5#Y��� I�����/� 1/sX/�!/�/y/�/ �/�/�/�/	?K/0?o/ �/c?Q?�?u?�?�?�? ?�?O�?�?�?)O_O MO�OqO�O�?�OO�O _�O__%_[_I__ �O�_�Oo_�_�_�_�_ oo!oWo�_~o�_Go �o�o�o�o�o�o	_o �oV�o/�w�� ���7�[�O� �_���s�����͏� �3���'��K�9�[� ��o����̟����� �#��G�5�W�}��� ���m�ׯů���� �C���j�|�3�U�/� ��ӿ������]�B� ���u�cυχϙ��� ����5��Y���M�;� q�_߁߃ߕ������ 1߻�%��I�7�m�[� }�������	������ !��E�3�i������ Y���U������� A��h��1��� ����[@ 	sa����� �3/W�K/9/o/ ]/�/�/�/��/�/�/ �/�/?G?5?k?Y?�? �/�?�/?�?�?�?�? OCO1OgO�?�O�?WO �O�O�O�O�O�O	_?_ �Of_�O/_�_�_�_�_ �_�_�_G_m_>o}_o qo_o�o�o�o�o�oo Co�o7�oGm[ ���o��� �3�!�C�i�W���� ���}��Տ���/� �?�e�����ˏU��� ���џ���+�m�R� d��=��������߯ ͯ�E�*�i��]�K� m�o�������ۿ�� A�˿5�#�Y�G�i�k� }ϳ�����ϣ���� 1��U�C�e߻��ϲ� �ϋ�����	���-�� Q��x��A��=�� �������)�k�P��� ���q����������� C�(g���[I m���� ? �3!WE{i� �������// /S/A/w/��/�g/ �/�/�/�/�/+??O? �/v?�/??�?�?�?�? �?�?�?'Oi?NO�?O �OoO�O�O�O�O�O/O UO&_eO�OY_G_}_k_ �_�_�__�_+_�_o �_/oUoCoyogo�o�_ �oo�o�o�o	+ Q?u�o��oe� �����'�M�� t��=�����ˏ��� ݏ�U�:�L��%��� m�����ǟ���-�� Q�۟E�3�U�W�i��� ��ï��)����� A�/�Q�S�e���ݯ¿ ��������=�+� Mϣ�ɿ��ٿs��ϻ� ������9�{�`ߟ� )ߓ�%ߣ��߷����� �S�8�w��k�Y�� }�������+��O� ��C�1�g�U���y��� �����'���	? -cQ�����w �s�;)_ ���O���� �//7/y^/�'/ �//�/�/�/�/�/? Q/6?u/�/i?W?�?{? �?�?�??=?OM?�? AO/OeOSO�OwO�O�? �OO�O_�O_=_+_ a_O_�_�O�_�Ou_�_ �_o�_o9o'o]o�_ �o�_Mo�o�o�o�o�o �o5wo\�o%� }�����="� 4����U���y��� ��ӏ���9�Ï-�� =�?�Q���u����ҟ �����)��9�;� M���ş���s�ݯ˯ ��%��5������� ��[�����ٿǿ��� !�c�Hχ��{�ϋ� �ϟ�������;� �_� ��S�A�w�e߇߭ߛ� �����7���+��O� =�s�a�������� �����'��K�9�o� �����_���[����� ��#G��n��7 ������� aF�yg�� ����9/]� Q/?/u/c/�/�/�/� %/�/5/�/)??M?;? q?_?�?�/�?�/�?�? �?�?%OOIO7OmO�? �O�?]O�O�O�O�O�O !__E_�Ol_�O5_�_ �_�_�_�_�_�_o__ Do�_owoeo�o�o�o �o�o%o
�o�o�o =sa����o��!+q�$SERV�_MAIL  �+u!���OUTwPUT�$�}@�RV 2�v;  $� (�q�<}��SAVE7�	��TOP10 2>W� d 'ݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w�������0��ѿ�u��YP����FZN_CFG ;�u$�~�����GRP 2��D� ,B �  A[�+qD;�� B\��  B�4~�RB21ފ�HELL��u��j�k�2�����%RSR������ �
�C�.�g�Rߋ�v� ���߬�����	���-��?�Q��  �_�%Q���_����,p�������g�2,pd�����HK 1�� ��E�@�R�d����� �������������*<e`r���OMM ������FTOV_ENB��_���HOW_R�EG_UI�	�IMIOFWDL� ��^�)WAIT����$V1��^�NTIM����VA�_)_�UNIT����L]CTRYB���MB_HDD�N 2W�  2�:%0 �pQ/�qL/ ^/�/�/�/�/�/�/�/��"!ON_ALI_AS ?e�	f�he�A?S?e?w?�: /?�?�?�?�?�?OO &O8OJO�?nO�O�O�O �OaO�O�O�O_"_�O F_X_j_|_'_�_�_�_ �_�_�_oo0oBoTo �_xo�o�o�o�oko�o �o,�oPbt �1������ �(�:�L�^�	����� ����ʏu�� ��$� Ϗ5�Z�l�~���;��� Ɵ؟����� �2�D� V�h��������¯ԯ ���
��.�ٯR�d� v�����E���п��� ϱ�*�<�N�`�r�� �ϨϺ���w����� &�8���\�n߀ߒߤ� O�����������4� F�X�j�|�'����� �������0�B��� f�x�������Y����� ����>Pbt ������ (:L�p�� ��c�� //$/ �H/Z/l/~/)/�/�/ �/�/�/�/? ?2?D?�V?]3�$SMON�_DEFPRO ����1� *S�YSTEM*0�m6RECALL �?}9 ( ��}4xcopy �fr:\*.* �virt:\tm�pback�1=>�147.87.1�49.40:15172 �2�>	OO+L}5�5a�?�?�6��?O�O�O}J�2m�db:schin�del_5sem�.tpMEemp\��M_O�O_)_ }9��4s:orderfil.datML`�OuO_�_�_}0�F JOc_�1p_�_o%o8C �?QO�_�_o�o�o<O Mo_orO�o'�O�O �O�O��8_J_�_ n_��#��_�o��_ �����4oFo�ojo|� ���o�oՏ�o���� ��0BTfc�	�� �����v����,� >�Y�b�t����)��� O�ܯ������:�K� ]�p����%ϸ�ʟܟ � ϑϣ�6�H�ѯl� ~��!ߴ�Ư����� �ߟ�2�D�׿h�z�� ﰿ¿����߉���.�
xyzrate 11 J�\�n�Ѐ��#�6���61 ����I��������9� K�]�oρ�$���� R�������5�G�b k�} �������� ���1�C�Tg�y 
//���������+/ �/-?Qt/��/? *?��/��/?�?�? ;�[?q�?O&O� �?�?�O�O�O�/�/ R?�/O_"_5?G?�O k?�O�_�_�?�?XO�? {_oo1OCO�_gO�_ �o�o�O�O�Oaowo�o -_?_�oc_�o����$SNPX_�ASG 2�����q�� P 0 '�%R[1]@1�.1��y?��s% �!��E�(�:�{�^� ������Տ��ʏ�� �A�$�e�H�Z���~� ��џ����؟�+�� 5�a�D���h�z����� ů�ԯ���
�K�.� U���d�������ۿ�� ����5��*�k�N� uϡτ��ϨϺ����� �1��U�8�Jߋ�n� ���ߤ���������� %�Q�4�u�X�j��� �����������;�� E�q�T���x������� ����%[> e�t����� �!E(:{^ ������/� /A/$/e/H/Z/�/~/ �/�/�/�/�/�/+?? 5?a?D?�?h?z?�?�? �?�?�?O�?
OKO.O UO�OdO�O�O�O�O�O �O_�O5__*_k_N_ u_�_�_�_�_�_�_�_ o1ooUo8oJo�ono�o�o�d�tPARAoM �u�q_ �	��jP�dU9p�ht��p�OFT_KB_CFG  �c�u�s�OPIN_SIM  �{vn���p�pRVQST_P_DSBW~r�"t�HtSR �Zy � & �SCHINDEL�_5SEM�u��vTOP_ON_?ERR  &�Dx~8�PTN Zu�k�A4�R?ING_PR�D���`VCNT_GOP 2Zuq�!px 	r��ɍ����׏��wVD��RP' 1�i p�y ��K�]�o��������� ɟ۟����#�5�G� Y���}�������ůׯ �����F�C�U�g� y���������ӿ�� 	��-�?�Q�c�uχ� �ϫ����������� )�;�M�_�qߘߕߧ� ����������%�7� ^�[�m������� ������$�!�3�E�W� i�{������������� ��/ASew ������� +=Ovs�� �����//</ 9/K/]/o/�/�/�/�/ �/�/?�/?#?5?G? Y?k?}?�?�?�?�?�?��?�?OO)�PRG�_COUNT8vq�k�GuKBENB���FEMpC:t}O_UP�D 1�{T  
4Or�O�O�O_ _!_3_\_W_i_{_�_ �_�_�_�_�_�_o4o /oAoSo|owo�o�o�o �o�o�o+T Oas����� ���,�'�9�K�t� o���������ɏۏ� ���#�L�G�Y�k��� ������ܟן���$� �1�C�l�g�y����� ����ӯ����	��D� ?�Q�c���������Կ Ͽ����)�;�d��_�q�=L_INFO� 1�E�@ �2@����������� ��±_�B+��!w'���2��mn��£n<LYSDOEBUGU@�@����d�If�SP_PA�SSUEB?x�L_OG  ���C���*ؑ�  ���A��UD1:�\�ԘΥ�_MPC �ݵE&�8�A��V�� �A�SAV �!�������X����SVZ�TEM_TIME 1"��]�@ 0�Љ���RX�X����$T1SVGUNS�@�VE'�E��AS�K_OPTION�U@�E�A�A+�_D�I��qOG�BC2_?GRP 2#�I�������@�  C����<Ko�CFG %z��� ������`��	�.>d O�s����� ��*N9r] �������/ �8/#/\/n/��Z+�/ Z/�/�/H/�/?�/'? ?K?]�k?=�@0s?�? �?�?�?�?�?O�?O O)O_OMO�OqO�O�O �O�O�O_�O%__I_ 7_m_[_}__�_�_�X � �_�_oo/o�_So Aoco�owo�o�o�o�o �o�o=+MO a������� ��9�'�]�K���o� ��������ɏ���#� �_;�M�k�}������ ��ß�ן��1��� U�C�y�g��������� ������	�?�-�c� Q�s����������Ͽ ����)�_�Mσ� 9��ϭ�������m�� �#�I�7�m�ߑ�_� �ߣ����������� !�W�E�{�i����� ����������A�/� e�S�u�w��������� ����+=O��s a������� 9']Kmo �������#/ /3/Y/G/}/k/�/�/ �/�/�/�/�/??C? ��[?m?�?�?�?-?�? �?�?	O�?-O?OQOO uOcO�O�O�O�O�O�O �O__;_)___M_�_ q_�_�_�_�_�_o�_ %oo5o7oIoomo�o Y?�o�o�o�o�o3 !CiW��� ������-�/� A�w�e���������� я���=�+�a�O� ��s�������ߟ͟� �o�-�K�]�o�ퟓ������ɯ���צ���$TBCSG_G�RP 2&ץ�  ��� 
 ?�   6�H�2�l�V���z���@ƿ�������(��d�E+�?~�	 HC����>���G����C�  A�.�e�q�wC��>ǳ33��"S�/]϶�Y��=Ȑ� C\  Bȹ���B���>���X�P���B�Y�z�"�L�H�0�$���� J�\�n�����@�Ҿ ���������=�Z�%�07����?3������	V3.0�0.�	cr35��	*����
���0������ 3���4�   {�CaT�v�}��J2��)������CFG� +ץ'� ,*������I����.<
� <bM�q��� ����(L7 p[����� �/�6/!/Z/E/W/ �/{/�/�/�/�/.�H� �/??�/L?7?\?�? m?�?�?�?�?�? OO $O�?HO3OlOWO|O�O ����Oӯ�O�O�O!_ _E_3_i_W_�_{_�_ �_�_�_�_o�_/oo ?oAoSo�owo�o�o�o �o�o�o+O= s�E���Y�� ���9�'�]�K�m� ������u�Ǐɏۏ� ��5�G�Y�k�%���}� ����ßşן���1� �U�C�y�g������� ӯ������	�+�-� ?�u�c���������� Ͽ���/�A�S��� ��qϓϕϧ������ ��%�7�I�[���m� �ߑ߳������߷�� 3�!�W�E�{�i��� �����������A� /�e�S�u��������� ������+a O�s��e��� ��'K9o] ������� #//G/5/k/}/�/�/ [/�/�/�/�/�/?? C?1?g?U?�?y?�?�? �?�?�?	O�?-OOQO ?OaO�OuO�O�O�O�O �O�O___M_�e_ w_�_3_�_�_�_�_�_ oo7o%o[omoo�o Oo�o�o�o�o�o! 3�o�oiW�{� ������/�� S�A�w�e�������я �������=�+�M� s�a���������ߟ� �_	���_ן]�K��� o�������ۯɯ��� #���Y�G�}�k��� ��ſ׿������� �U�C�y�gϝϋ��� ���������	�?�-� c�Q�s�u߇߽߫��� �����)��9�_�M� ����/����i���� ��%��I�7�m�[��� ���������������� EWi{5�� ������A /eS�w��� ��/�+//O/=/ _/a/s/�/�/�/�/�/ �/?'?��??Q?c?? �?�?�?�?�?�?�?O �?5OGOYOkO)O�O}Op�O�O�O�N  �@�S V_R��$TBJOP_G�RP 2,�E��  ?��V	-R4S.;\=��@|u0{S~PU >��U�T @�@LR	� �C� �Vf?  C���ULQ�LQ>�33�U�R�����U�Y?�@=��ZC��P�����R��P  Bȸ�W$o/gC��@g��dDb�^�㙚eeao�P&ff~�e=�7LC/kFaB o�o�P��P��efb-C�p�B�^g`�d�o�PL�P�t<�eVC\ � �Q@�'p�`��  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�anaaF`C�;�`L�w��aQoxp�x�p:���XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb����X �	��1��)�W��� c������������ 󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSc7r35QT*�QT��A�� E��'E�i�F�V#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG��G#
�D���E'
E�MKE���E��ɑE�ۘE���E���F���F��F���F(��F�5��FB��F�O��F\��F�i��Fv��F���vF�u�<#�
<t����ٵ=�_��V �R�p�V9�~ ]ESTPARtp��HFP*SHR\�A�BLE 1/;[$%�SG�� �W�
G�G�G� WQG�	G�
G�GȖ�QG�G�G�ܱv�'RDI~�EQ�ϧ� ��������W�O_�q�@{ߍߟ߱���w�S]�CS !ڄ������ ������&�8�J�\� n������������� ] \�`��	��(�:� ����
��.�@�w��NUM  �EUEQ�P	P ۰�ܰw�_CFG �0��)r-PIMEBF_TTb��CSo�,VERڳ-B�,R 11;[' 8��R�@� �@&  ��� ����//)/;/ M/_/q/�/�/�/�/�/ ?�/?J?%?7?M?[? m?>�@�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_��_l_�Y@c�Y�MI_CHAN�8 c cDBGLV��:cX�	`�ETHERAD �?f�\`���?�_uo�oQ�	`RO�UTV!	
!��d�o�lSNMAS�KQhcba255.uߣ'9ߣY��OOLOFS_D�Ib��U;iORQCTRL 2		�Ϸ~T��� ��#�5�G�Y�k�}� ������ŏ׏�����.��R�V�PE_�DETAI/h|zP�GL_CONFI�G 8�	����/cell/$�CID$/grp1V�̟ޟ�������o?�Q�c�u����� (���ϯ������ ;�M�_�q�����$�6� ˿ݿ���%ϴ�I� [�m�ϑϣ�2����� �����!߰���W�i� {ߍߟ߱�%}F��� ����/�A�C�i�H�Eߞ�������� ��?��.�@�R�d�v� ������������� ��*<N`r� ������& 8J\n��!� ����/�4/F/ X/j/|/�//�/�/�/ �/�/??�/B?T?f? x?�?�?+?�?�?�?�? OO�?>OPObOtO�O��O�O���Us�er View ���}}1234567890�O�O�O�_#_5_=T�P��]_���I2�I:O�_�_�_@�_�_�_X_j_�B3�_ GoYoko}o�o�o o�op^46o�o1CU�ovp^5�o������	�h*�p^6 �c�u����������ޏp^7R��)�;�M� _�q�Џ��p^8�˟ ݟ���%���F�L�� lCamera�J���� ����ӯ���E~�� !�3��OM�_�q��������y  e��Yz��� 	��-�?�Q���uχ� ��俽���������>��e�5i��c�u߇� �߽߫�d������P� )�;�M�_�q��*�<� �i���������)� ��M�_�q�������� ��������<�û��= Oas��>��� �*'9K] f�Q������ �/�%/7/I/�m/ /�/�/�/�/n<�� ^/?%?7?I?[?m?/ �?�?�? ?�?�?�?O !O3O�/<׹��?O�O �O�O�O�O�?�O_!_ lOE_W_i_{_�_�_FOXG9+_�_�_oo(o :o�OKopo�o)_�o�o@�o�o�o ��	g�0�oM_q��� No����o�%�7� I�[�m�&l�n�� Ə؏���� ��D� V�h���������ԟ 柍�g�ڻ}�2�D�V� h�z���3���¯ԯ� ��
��.�@�R���3u F�鯞���¿Կ��� ���.�@ϋ�d�vψ� �ϬϾ�e�w���U�
� �.�@�R�d�ψߚ� ������������*� ��w���v���� ����w�����c�<� N�`�r�����=�w�� -�����*<�� `r�������x���  �� 1CUgy��������    -/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_�i_�  
��( � �%( 	 y_�_�_�_�_�_�_ o	o+o-o?ouoco�o�o�o�Z* � Q&�J\n ������o��� 9�(�:�L�^�p�� �������܏� �� $�6�}�Z�l�~�ŏ�� ��Ɵ؟���C�U�2� D�V���z�������¯ ԯ���
��c�@�R� d�v�����᯾�п� )���*�<�N�`ϧ� ���ϨϺ������� �&�8��\�n߀��� �߶���������E�"� 4�F��j�|���� ��������e�B� T�f�x����������� ��+�,>Pb ���������� (o�^p� ������ /G $/6/H/�l/~/�/�/ �/�//�/�/?U/2?�D?V?h?z?�?�/�`@� �2�?�?�?�3��7�P��!frh�:\tpgl\r�obots\m2�0ia\cr35?ia.xml�?;O MO_OqO�O�O�O�O�O�O�O ���O_(_ :_L_^_p_�_�_�_�_ �_�_�O�_o$o6oHo Zolo~o�o�o�o�o�o �_�o 2DVh z������o� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟�ݟ��&�8� J�\�n���������ȯ ߟٯ���"�4�F�X� j�|�������Ŀ־�8�.1 �?@8?8�?�ֻ� ֿ�3�5�G�iϓ�}� ���ϳ��������5߀�A�k�U�wߡ߿���$TPGL_OUTPUT ;�!��! �� ������,�>�P�b� t����������� ��(�:�L�^�p������������2345678901�� �������"�� BTfx��4�@����
}$ L^p��,>� �� //$/�2/Z/ l/~/�/�/:/�/�/�/ �/? ?�/�/V?h?z? �?�?�?H?�?�?�?
O O.O�?<OdOvO�O�O �ODOVO�O�O__*_ <_�OJ_r_�_�_�_�_ R_�_�_oo&o8o�_ �_no�o�o�o�o�o`o �o�o"4F�oT�|����\��} �����0�B�T�e��@������� ( 	 ��Џ��� ���<�*�L�N�`� ��������ޟ̟�� �8�&�\�J���n��� ������ȯ���"�������*�X�j�F��� ��|�¿Կ��C���� ��3�E�#�i�{�忇� ��S����������/� ��S�e�߉ߛ�y߿� ��;�������=�O� -�s���ߩ��]��� �����'����]�o� �����������E��� ��5G%W}�� ����g��� 1�Ug	w�{ ��=O	//�?/ Q///u/�/��/�/_/ �/�/�/�/)?;?�/_? q??�?�?�?�?�?G? �?O�?OIO[O9OO �O�?�O�OiO�O�O�O !_3_�O_i_{__�_�_�_�_�_�R�$T�POFF_LIM� >�op:�y�mqbN_SV`�  l�jP_�MON <6�)dopop2l�a�STRTCHK �=6�f� bVTCOMPAT-h��afVWVAR �>Mm�h1d ��o �oop`b�a_DEFPRO�G %|j%S�CHINDEL_�5SE`Nif_D?ISPLAY`|n�"rINST_MSwK  t| ^z?INUSER�odt�LCK�|}{QUI�CKMEN�dtS7CRE�p6��b?tpscdt�q���b*�_.�ST��jiRACE_C_FG ?Mi�du`	�d
?�u��HNL 2@|i����k r͏ߏ���'�9�K�]�w�I�TKp2A�� ��%$123456�7890����  �=<��П��  #!���p��=� �c��^��������� �.���R��v�"�H� ί��Я������*� ֿ���r�2ϖ����� 4�޿�ϰ���&���J� \�n���@ߤ�d�v��� �������4���X�� *��@�����ߨ� ������T���x�� �����l�������� ,�>�P�������FX ��d������: �p"��o� ����F6HZ t~��N/t/�/� �// /2/�/V/?(? :?�/F?�/�/�/j?�? ?�?�?R?�?v?�?QO �?lO�?�O�OO�O*O |O_`O _�O0_V_h_ �Ot_�O__�_8_�_ 
oo�_@o�_�_�_Lo do�_�o�o4o�oXojo 3�oN�or��o�P�s�S�B��>�z�  h��z� ��C�:y
 �P�v�]����UD�1:\�����qR_GRP 1C���� 	 @ Cp���$��H�6�l�Z��|�����f����˟���ڕ?�   
���<�*�`�N��� r�������ޯ̯���&��J�8�Z���	�u�����sSCB ;2D� ��� ��(�:�L�^�pς���|V_CONFIG E���@�����ϖ�OUTPUT� F�������6�H�Z�l�~ߐ� �ߴ������������ #�6�H�Z�l�~��� ������������2� D�V�h�z��������� ������
�.@R dv������ �)<N`r �������/ /%8/J/\/n/�/�/ �/�/�/�/�/�/?!/ 4?F?X?j?|?�?�?�? �?�?�?�?OO/?BO TOfOxO�O�O�O�O�O �O�O__+O>_P_b_ t_�_�_�_�_�_�_�_ oo'_:oLo^opo�o �o�o�o�o�o�o  $����!�bt�� �������(� :�-o^�p��������� ʏ܏� ��$�6�G� Z�l�~�������Ɵ؟ ���� �2�D�U�h� z�������¯ԯ��� 
��.�@�Q�d�v��� ������п����� *�<�M�`�rτϖϨ� ����������&�8� J�[�n߀ߒߤ߶��� �������"�4�F�W� j�|���������� ����0�B�S�f�x� �������������� ,>Pa�t�� �����(�:L/x��� k}gV�K�� �//&/8/J/\/n/ �/�/�/W�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�/�?�?�?OO 0OBOTOfOxO�O�O�O �?�O�O�O__,_>_ P_b_t_�_�_�_�O�_ �_�_oo(o:oLo^o po�o�o�o�o�_�o�o  $6HZl~ ����o����  �2�D�V�h�z����� ���ԏ���
��.� @�R�d�v��������� Ϗ�����*�<�N� `�r���������˟ޯ ���&�8�J�\�n����������Ż�$T�X_SCREEN� 1G�g�}ipn�l/��gen.htmſ�*�<�N�`���Panel� setupd�}�dϥϷ����������ω�6�H�Z�l�~� ��ߴ�+��������  �2�߻�h�z��� ����9�g�]�
��.� @�R�d��������� ������}���<N `r��;1� �&8�\� ������QȾ�UALRM_MS�G ?��� �Ȫ-/?/p/c/�/ �/�/�/�/�/�/??�6?)?Z?%SEV � -�6"E�CFG I���  ȥ@��  A�1   B�Ȥ
 [?ϣ� �?OO%O7OIO[OmO�O�O�O�G�1GRPw 2J�; 0Ȧ�	 �?�O I_�BBL_NOTE� K�:T���lϢ�ѡ��0RDEFPROz %+ (%N? u_Ѡc_�_�_�_�_�_ �_o�_o>o)oboMo��o\INUSER�  R]�O�oI_�MENHIST �1L�9  (� _P��(/S�OFTPART/�GENLINK?�current=�menupage?,955,1�oC�Ugy,15�30�����p2��uedit(rD�EMOPICKPLACE�S�e�w�2�x'�~71B�̏�ޏ����q)��$�ZERO��R�d�v���� �3�$�SCH�INDEL_TEST,18�����������wintp �p��B�e�w����*���5SEMA���� ��g9Rq|oB�T�f� x������s1�ƿؿ� ��� ϯ�D�V�h�z� �Ϟ�-���������
� ߫Ͻ�R�d�v߈ߚ� ��;���������*� ��N�`�r����7� I�������&�8�#� \�n������������� ����"4F��j |����S�� 0BT�x� ����a�// ,/>/P/�t/�/�/�/ �/�/�/o/??(?:? L?^?I��?�?�?�?�? �?�?�/O$O6OHOZO lO�?�O�O�O�O�O�O yO_ _2_D_V_h_z_ 	_�_�_�_�_�_�_�_ o.o@oRodovoo�o �o�o�o�o�o�o* <N`r�o?� �����8�J� \�n�����!���ȏڏ ��������F�X�j� |�����/�ğ֟��� ����B�T�f�x��� ��+�=�ү����� ,���P�b�t���������z�$UI_PA�NEDATA 1�N���ڱ�  	�}�/frh/cg�tp/wided�ev.stm _���th=800&�_height=�92&_��ice�=TP&_lin�es=11&_c�olumns=4~�font=3��page=who�l����7�)prsimYς�  }����ϻ�������� ) �)��M�4�q߃�j� �ߎ����������%��7��[�7����    �(�X���doub��2�������8����>�ual��"� ��F�X�j�|�����G� ����������B T;x_������i� ݰܳ7� <N`r���� -���//&/8/� \/n/U/�/y/�/�/�/ �/�/?�/4?F?-?j? Q?�?�?%�?�?�? OO0O�?TO�xO�O �O�O�O�O�OKO_�O ,__P_b_I_�_m_�_ �_�_�_�_oo�_:o �?�?po�o�o�o�o�o o�o sO$6HZ l~�o����� �� �2��V�=�z� ��s�����ԏGoYo �.�@�R�d�v�ɏ�� ��П������ <�N�5�r�Y������� ̯���ׯ�&��J� 1�n�������ȿڿ ����c�4ϧ�X�j� |ώϠϲ���+����� ���0�B�)�f�Mߊ� �߃��ߧ�������� ����P�b�t���� ������S���(�:� L�^����i������� ���� ��6Z�lS�w�'�9�}���"4FX)�}��l��� ��/j'//K/2/ D/�/h/�/�/�/�/�/ �/�/#?5??Y?��C��=��$UI_PO�STYPE  �C�� 	� e?�?�2QUI�CKMEN  �;�?�?�0RESTORE 1OC��  ��*defa�ult�;  O�UBLE�=P�RIM�?med�itpage,S�CHINDEL_?5SEM,1fO�O��O�OjLmenu~B955�O__+_ =_pFF_j_|_�_�_�_ EAL?�_�_G_�_"o4o FoXojoo�o�o�o�o �oyo�o0B�_ Oas�o���� ���,�>�P�b�t� �������Ώ���� �����L�^�p����� 7���ʟܟ� ���$� 6�H�Z�l��!����� ������� �2�կ V�h�z�����A�¿Կ����
��=SCRE��0?�=uw1sc+@u2K�U3K�4K�5K�6K��7K�8K��2USE1R-�2�D�ksMì�U3��4��5��6���7��8���0NDO_CFG P�;�� ��0PDATE� ���N�one�2��_IN_FO 1QC�@��10%�[���Iߊ� m߮��ߣ�������� ��>�P�3�t��i����<-�OFFSET T�=�ﲳ$@ ������1�^�U�g� ��������������� $-ZQcu����?�
����UFWRAMO@�����*�RTOL_AB�RT	(�!ENB�*GRP 1U�I�1Cz  A��~��~���������0U�J�9MSK  �M@�;N%�8�%��/�2VCC�M��V�ͣ#RG��#Y�9���/��Z��D�BH�p7�1C���3711?ـC0�$MRf2_��*S�Ҵ�	����~XC56 �*�?�6���1$��5���A@3C���. ��8 �?��OOKOx1FOsO"�5�51��_O�O��� B��� �A2�DWO�O7O_�O 8_#_\_G_�_k_}_�_ _�_�_�_�_"o�OFo\Xo�%TCC�#`mPI1�i������ �GFS��2aZ;� �| 2345678901�o�b�� ���o��!5a�$4BwB�`56 311?:�o=L�Br5 v1�1~1�2��}/��o �a��#�GYk }�p������� ُ�1�C�U�6�H��� 5�~���ߏ���	��|�4�dSELEC)�M!v1b3�VIR�TSYNC�� ����%�SIONT�MOU�������F��#bU���U�(u �FR:\H�\�A�\�� �� �MC��LOG�� �  UD1��E�X����' B@ ����̡m�|�̡  OBCL��1�H� � � =	 1- �n6  -�������[�,S�A�`=���͗��ˢ>��TRAIN⯞b(�a1l�
0d�$j�:T2cZ; (aE2 ϖ�i��;�)�_�M� g�qσϕϧ���������	��F�STAT' dm~2@�z�Č�*j$i߾��_GuE�#eZ;�`0��
� 02��HO�MIN� fU��U� ~������БC�g�X���JMPERR 2gZ;
  ��*jl�V� 7�������������� 
��2�@�q�d�v�B�-_ߠRE� hWޠ$�LEX��iZ;�a1�-e��VMPHA�SE  5��c&��!OFF/�F��P2n�j�0�㜳E1@��0ϒ<E1!1?s33�����ak/�kxk��!W�m[�䦲�[�����o3;� [i{� ���/�O� ?/M/_/q/��/��/ /�/'/9/�/=?7?I? s?�/�?�/�/�?�?? Om?O%O3OEO�?�? �O�?�O�O�?�O�O�O __gO\_�OE_�O�_ �O�O/_�_�_�_oQ_ Fou_�_|o�o�_�oo �o�o�o�o;oMo?qo f-�oI���� �7�[P�� �������ˏ��!� 3�(�:�i�[�ŏg�}�������TD_FI�LTEW�n�� �ֲ:���@��� +�=�O�a�s������� ��֯�����0��B�T�f�x���SHI�FTMENU 1-o[�<��%��ֿ ����ڿ����I� � 2��V�hώ��Ϟϰ��������3�
�	L�IVE/SNAP�'�vsfliv���E����IO�N * Ub�h�menu~߃�����ߣ�l����p���	�ؘ��E�.�50�s�P�@� ��AɠB8z�z��}��rx�~�P�� ,���MEb���<��0���MO��q����z�WAIT�DINEND�������OK1�O�UT���SD��T�IM����o�G ���#���C���b�������RELEAS1E������TM����{���_ACT[������_DATA' r��%L��<��xRDISb�E��$XVR�s����$ZABC_�GRP 1t�*Q�,#�0�2���ZIP�u'�&����[MPCF�_G 1v�Q�0�/� w�ɤ�� 	�Z/  85�/�/H/�/l$?��+�/�/�/?��/�/???r?�?  �D0�?�?�?�? �?�;���x�]�hYLIND֑y�� ��� ,(  *VOgM.�SO0�OwO�O�M i?�O �O^PO1_�OU_<_N_ �_�O�_�_�__�_�_ x_-ooQo8o�_�o�o�Y&#2z� ���oC�e?a?>�N|�oq����qA��$DSPHERE 2{6M��_�;o� ��!�io|W�i��_ ��,��Ï���Ώ@� �/�v���e�؏��p�����������ZZ�� �N