��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �� �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LAJ1R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B�ASBNw_CF>"
 8F CNV_J� ; �"��!_CMNT�?$FLAGS]��CHEC�8 � E�LLSETUP {� $HO30�IO�0� %�SM�ACRO�RREP	R�X� D+�0��R�{�T UTOBA�CKU�0� �)DEVIC&�CTI*0�� �0�#�`B�S$IN�TERVALO#I?SP_UNI�O`�_DO>f7uiFR3_F�0AIN�1����1c�C_WAxkda�jOFF_O0]N�DEL�hL� p?aA�a1b?9a��`C?��P�1E���#sATB�d���MO� �cE �D [M�c��^qR;EV�BILrwJ1�XI� QrR � � OD�P�q_$NO^PM�Wp�t�r/"�w� ��u�q�r�0D`S� p E RD�_E�pCq$FS�SBn&$CHKBoD_SE^eAG �G�"$SLOT!_��2=�� V�d�%���3J0a_ED�Im   � )�"��PS�`(4�%$EP�1�1$�OP�0�2�a�p_�OK�UST1P_�C� ��d��U �PLACI4!�Q�4�<( raCOMM� ,0$D����0�`���EOWBn�IGALL;OW� (K�":(2�0VARa��@h�2ao�L�0OUy�� ,Kvay��PS�`�0M_O]�����CCFS_U	T~p0 "�1�3�#��ؗ`X"�}R0 { 4F IMCM�`O#S�`��upi �)_�p�BAJ1����M/ h�pI?MPEE_F�N���N���@O��r�DQ_�~�n�Dy�F�� dCC_�r0 � T� '��'�DI��n0"��p�P�$I�������F�t X� GR�P0��M=qNFL�I�7��0UIRE��$g"� SWIT{CH5�AX_N�P�Ss"CF_LIM~� � �0EED��!��qP�t��`PJ_dVЦMODEh�.Z`�PӺ�ELBOF� ��� ���p� ���3���� FB/��0�>��G� �� WA'RNM�`/��qPܚ�n�NST� CO�R-0bFLTR^h�TRAT�PT1�>� $ACC1a���N ��r$ORIأo"V�RT�P_S\�J0CHG�0I�E�rT2��1�I���T�I1��� �x i#�Q��H�DRBJ; CQ�2�L�3L�4L�5L�6�L�7L� N�9s!z��O`S <F �+�=�O��#92��LL�ECy�"MULTI�b�"N��1�!�Ѻ�0T�� �S�TY�"�R`�=l�)�2`����*�`T  �|� �&$��۱m�0�P�̱�UTO���E��EXT����Á8B���"2� (�
��![0������<�8b+�� "D"�� �ŽQ��<煰kc��'�9�#���1��ÂM8�ԽP��" '�3�$ L� E���P�<��`A�$JOB�n�T���l�TRIG3�% dK��������<���\��+�Y�p�_yM��& t�p3FLܐBNG AgTBA� ���M��
 �!��p� �q��0�aP[`��O�'[����0tna*���"J���_R���CDJ���IdJk�D�%C��`�Z���0��P_��P��@ ( @F RaO.��&�t�IT�c�NOM�
���P�S���`T)w@����Z�P�d���RA��0��2b"����
$�T����MD3�TD��`U31���p(5!YHGb�T1�*E�7�c�KAb�WAb�cA�4#YNT���PD'BGD�� *(��PUt@X��W����AX��a��eTAI^cBUF��0!�+ � 7n�P�IW�*5 P�7M��8M�9
0�6F�7S�IMQS@>KEE�3PATn�^�a"� 2`#�"�L64F;IX!, ���!dĶ�D�2Bus=CCI��:FPCH�P:BAD�aHCEhAOGhA]H"W�_�0>�0_h@�f �Ak���F�q\'M`#��"n HE3�- l�p3G��@FSOES]FgHBSU�IBS9W|C��. ` ���MARG쀳��F�ACLp�SLEW�xQe�ӿ��BM�C�/�\pSM_JBM����QYC	g��e#�0 �n��CHN-�MP�G$G� Jg�_� <#��1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�fJR���rSEG�FR�PIO� S�TRT��N��cP!V5���!41�r�Ӏ
r>İ�b�B�O�2` +�[��� ,qE`&�,q`y�Ԣ}t8��yaSIZ%����t�vT�s� �z�y,qRSINF}Oбc����k��`��`�`Lp�ĸ T`7�CRCf�ԣCC/�9��`a�ua8h�ub'�MIN��uaPDs�#�G�D�YC��C�����e�q0��� ��EV�q�F�_
�eF��N3�s�ahƔ�Xa+p,5!�#=1�!VSCA?� �A��s1�"!3 ��`F/k��_�U��g�@�]��C�� a�s��}R�4� �ߠ��N����5a�R�HwANC��$LG��lP�f1$+@NDP�t�AR5@N^��a�q���c��ME�18����}0��RAө�AZ� 𨵰�%O��FCATK��s`"�S�P.FADIJ�OJ�ʠ �ʠ���<���Ր���GI�p�BMP��d�p�Dba��AESآ@	�K�W_��BA�S�� �G�5  �M�I�T�CSXh[@@�!62�	$X�K��T9�{sC���N�`�a~P_HEIsGHs1;�WID�06�aVT ACϰ��1A�Pl�<���EXqPg���|��CU�0_MMENU��7�TIT,AE�%�)�a2��a��8 YP� a�ED�E.`��PDT��REM�.��AUTH_K�EY  ������ ��b�O	��}1E�RRLH� �9 \�� �q-�OR�DB�_�ID�@l �PUN_�O��Y�$SYSP0��4g�-�I�E��EV�#q'�PXW�O�� �: $S�K7!f2&�Td�T�RL��; �'AqC�`��ĠIND9�DJ.D��_��f1X��f���PL�A�R#WAj���SD�A���A+r|��UMM3Y9d�F�10d�&�d��J�<��}1PR�w 
3�POS���J�= �$�V$�q �LB~�>���ܠK�?�����CJ�@����EN5E�@T��A���_�RECOR��B�H 5 O�@7=$LA�>$~�r2��R��`�q�b`�_DLu��0RO�@�aT[� Q��b������! }О��PAUS���dE�TURN��MR�U�  CRp�E�WM�b�AGNAL:s2$LA�!�?$PX�@$P�y A �Ax�1C0 #ܠDO�`X��k�W�v�q�GO_A7WAY��MO�ae����]�CSS_C�CSCB C �8'N��CERI����J`u�QA0�}���@�GAG� R �0�`��{`��{`OF�q�5��#kMA��X��X&���LL�D� �$���sU�D)E%!�`���OVR10�W�,�OR|�'�$�ESC_$`�eDSGBIOQ��l �\�B�VIB&� �c�,�����f�=pSS�W���f!VL��P�L���ARMLO�
��`����d7%SC �bALspH�MPCh �Ch �#h �#h 5�UU���C �'�C�'�#�$'�d�#AC\4�$�pH��Ou�0�!Y��!�SB�� �`k$4�C�P3Wұ~46$VOLT37#$$`�*�^1�0�$`O1*�$o��0�RQY��2b4�0DH_THE����0xSЯ4�7ALPH�4�`���7�@ �0�qb7�rR�5�88� �×���"��Fn�MӁVHBPFUBAFLQ"D�s�`�THR��i2dB�����G(��PVP�����(������1�J2�B�E�C�E�CPSu�Y@� �Fb3���H�(V�H:U �G�
X0��FkQw�[��Na�'B���C IN{HBcFILT�� �$��W�2�T1�[� ��$���H Y6АAF�sDO��Y �Rp� fg�Q�+�c�5h�Q�iSh�QPL��Wqi�QTMOU �#c�i�Q\��X�gmb���vi�h�bAi�fI��aHIG��ca	xO���ܰ��W�"vAN�-u!��	#AV�H!Pa8$P�ד#p��R_:�A�a��B��N0�X�MCN`���f1[1�qVE�p��Z2;&f�I�QO�uh�rx�wGldDN{G|d��aF>!�9�r�aM:�U�FWA�:�Ml���X�Lu��$ !����!l�ZO�����0%O�lF�s�13�D	I�W�@��Q����_��!CURV�A԰0rCR41ͰZ �C<�r�H�v���<�`0��<�(�f�CH�QR 3�S���t���Xp�VCS_�`�ד�F��rژ�����NSTCY_ 'E L����1�t��1��U��24�2B�N�I O7������DE�VI|� F���$5�RBTxSPeIB�P���BYX䱠��T��HND}G��G H tn���L��Q�C�迁5��Lo0 H0��閻�FBP�{tFE{�5�t��T���I�DO���uPMCS�v>�f>�t�"�HOTSW�`s��?ELE��J T����e�2��25�� O� ��HA7�E��344��0	?��A�K �� MDL� 2J~PE��	A��s��tːÈ�s�JÆG!�rD"�ó�����\�T�O��W�	��/��S�LAV�L  �0INPڐ���`%��_CFd�Mw� $��ENU��OG��b�ϑ]զP�0�`ҕ�]�IDMaA�Sa��\�WR�#���"]�VE�$a�SKI�STs��sk$��	2u���J�������p	��Q���_SVh�EXCLUMqJ2M!'ONL��D�Y��|r�PE ղI_V��APPLYZP��HcID-@Y�r�_M�2=��VRFY�0��xr�1�cIOC_f�D�� 1������O���u�LS���R$D_UMMY3�!��z�S� L_TP/B�v�"���AӞ�ّ �N ���RT_\u�� >G&r�[�O D��P_B�A�`�3x�!IF ��_5���H������� �� P� $�KwARGI���� q�2O ��SGNZ�Q �8~P/�/PIGNs�l�$�^ sQANNUN�@�T<0�U/�ߴ�LAzp]	`Z�d~�EFwP}I�@ R @��F?IT�	$TOTA%��d���j�!�M�NIY�CS+���E�A[��
DAYS\�AD�x�@��	� �E�FF_AXI?�T�I��0zCOJA ��ADJ_RTRQ��Up��<P�1D �r5̀Ll�T�0? ]P�"p��m8tpd��V 0w��G��������SK��SU� ��CTR�L_CA�� W>�TRANS�6PIDLE_PW����!��A�V��V_��l�V �DI�AGS���X� �/$2�_SE�#TAC���t!�!0z*L@��RR��vPA��4�p ; SW�!�! �  ��ol�U��o3OH��PP� ��sIR�r��BRK'#��"A_Ak���x 2 x�9ϐZs2��%l��W�0t*�x%RQD�W�%MSx�t5AX��'�"��LIFEC�AL���10��N �1{"�5Z�3{"dp5�xZU`}�MOTN°9Y$@FLA�cZgOVC@p�5HE	>��SUPPOQ�ݑ�Aq� Lj (C�1_�X6�IEYRJZRJW�RJ�0TH�!UC��6�X�Z_AR�p��Y2��HCOQ��Sf6A�N��w$�ICT�E�Y `��CACHE�C9�M��PLAN��UFFIQ@�Ф0<�1�	��6��MSW��EZ 8�KEY�IM�p��TM~�S�wQq�wQ#���TRO�CVIE� �[ A�BGL��/�}�G?� N�?��D\p�mذST��!�R � �T� �T� �T	��PEMAIf�ҁо�_FAUL�]$�Rц�1�U�КR��DTRE�^�< $Rc�uS��% IT��BUF�W}�W��N_� SUB~d��C|��Sb�q�bSAV�e�bu @�B��� �gX�^P�d�u+p�$�_~`�e�p�%yOTT����sP¯�M��OtT�LwAX� � ��X~`9#�c_uG�3
�YN_1��_�D��1 ��2M���T�F���H@ g�`�� 0p��Gb-sC_R�AIK���r��t�RoQ�u7h�qD�SPq��rP��A�I�M�c6�\����s2�U��@�A�sM*`IP����s�!D��6�TH��@n�)�OT�!6�H�SDI3�ABSC���@ Vy��� ��_D�CONV�I�G���@3�~`F��!�pd��psqSqCZ"���sMERk���qFB��k��pET����aeRFU:@D�Ur`����x�CD�,���@p;cHR�A!��bp�ՔՔ+�PSԕC���C���pTQғSp�c/H *�LX�:c d�Rqa�| ����W�� U��U��U�	�U�OQ*U�7R�8R�9R��0TT�^�1k�1x�1��U1��1��1��1���1ƪ2Ԫ2^�k�2�x�2��2��2��2���2��2ƪ3Ԫ3^�3k�x�3���o����3��3��3ƪ46Ԣ�HXTk!0�d <� 7h�p�6�p�O��p����NaFDR^Z$eT^`V��Gr����䂴2REMr� Fj��BOVM�z�A�TROVٳDT�`-�MX<�I�N��0,�W!IND�KЗ
w�׀�p$DG~q36��P�5�!9D�6�RIV���2��BGEAR�IO�%K�¾DN�p��J��82�PB@�CZ_MCCM�@�1��@U���1�f ,②a?� ���PI�!K?I�E��Q�
��H�`m���g� _0Pfq�g RI9ej�k!UP2_ h � �cTD�p���! a�t�����BAC�r�i T�P�b�`�) OG��%���p��IFI�!�pm�>���	�PT�"��M�R2��j  ��Ɛ+"����\�����@���$�B`x%��_ԡ��ޭ_���� M�������DGCLF��%DGDY%LDa��5�6�ߺ4@��U�k��� T�sFS#p�Tl P���e�qP�p$EX_���1M2��2j� 3�5��G ����m ��Ѝ�SW��eOe6DEBUG����%GR���pUn�#BKU_�O1'�7 �@PO�I�5�5MS��OYOfswSM��E�b��@�0�0_E �n �0�CH__�TERM�o��Ɛ�ORI+�p<�N��SM_���b��q�m�T�A�r�P�UP>�Rs� -�1�2�n$�' o$S�EG,*> ELTO���$USE�pNFIAU"4�e1��|�#$p$UFR����0ؐO!�0����OT��'�TAƀU�#N;ST�PAT��P��"PTHJ����Ep�P rF�V"ART�`�`%B`�abU!REL<:�aSHFT��V!\�!�(_SH+@M$�D��� ��@N8r�����OVRq��rSH�I%0��UN� �aAGYLO����qIl�����!�@��@ERV ]��1�?:�¦'�2`��%��5�%�RCq��EASYM�q�EV!#WJi'��}�E���!I�2��U@D��q�%Ba��
5Po��0�p6�OR�MY� `GR��t2b5n� � p��UPa�Uu Ԭ"�)���TOCO!S�1POP ��`�p(C�������Oѥ`KREPR3��aO�P,�b�"ePR�%WU�.X1��e$PWRf��IMIU�2R_	S��$VIS��#(AUqD���Dv" v���$H���P_AD+DR��H�G�"�Q��Q�QБR~pDp1�w H� SZ�a��e`�ex�e��SE�l�r��HS��MNv?x ���%Ŕ��OL���p<Px��-��ACROlP<_!QND_C��גx�1�T �ROUPT���B_�VpQ�A1 Q�v��c_��i���iр�hx��i���i��v�AMCk�IOU��D�g�fsu^d�y $|�P_D��VB`boPRM_�b�A�TTP_אHaz{ (��OBJEr�l�P��$��LE�#��s`{ � \��u�AB_x�T~��S�@�DBGL�V��KRL�YHIoTCOU�BGY �LO a�TEM���e�>�+P'�,PSS�|�P�JQUERY�_FLA�b�HW(��\!a|`u@�3PU�b�PIO��"��]�ӂ/dԁ=dԁ�� _�IOLN��}�����CXa$SL�Z�$INPUTM_g�$IP#�P��L'���SLvpa~���!�\�W�C-�B$�I�O�pF_ASv��$L ��w �F1"G�U�B0m!���0HY��ڑ����UOPs� ` ������[�ʔ[�і"�[PP�SIP�<�іI��2���P_MEMBܿ�i`� X��IP�P�b{�_N�`�����R�����bS�P��p$FOCUgSBG�a��UJ�Ə� �  � o7JsOG�'�DIS[�J7�cx�J8�7�� Im!�)�7_L�AB�!�@�A��A7PHIb�Q�]�D� J7J\���� �_KEYt� {�KՀLMONa=���$XR��ɀ��WAT���3��&�EL��}Sy����&s� �Ю!V�g� �CTR3򲓥��;LG�D� �R���I�
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�G� �I�F�%SO���q �ƀ����v��ƴ��K�S ���w�k�N����E��\���D'�*�U�s5��@L>�n4�DAUZ�EA�p0Հ�Dp�f�GH�B��BOO���3 C���PIT����� ��REC��SCRN����D_p�aMARGf�`��:� ��T�L���S�s���W�Ԣ�Iԭ�JGM�O�MNCH�c��F�N��R�Kx�PRG�v�UF��p0��FW�D��HL��STP���V��+���Є�RES��H�@�몖Cr4@��?B��� +�O�U�q���*�a28����Gh�0PO��������M8�Ģ��EX��TKUIv�I��(� 4�@�t�x�J0J� ~�P��J0��N�a�#�ANA��O"�0VA�IA��dCLEAR~�6DCS_HI"��/c�O�O�S�I��S��IGAN_�vpq�uᛀT�dn� DEV-�LLAL �°BUW`��x0T<$U�E�M��Ł��s��0�A
�R��x0�σ�a��@OS1�2�3���� `� ��ࠜh�AN%-���-�IKDX�DP�2MRO�X�Գ!�ST��Rq��Y{b! �$E&C+��p.&A&q
���`� L���ȟ%Pݘ��T\Q�UE�`�Ua��_ � �@(��`�����# �MB_PN@ �R`r��R�w�TRIqN��P��BASS\�a	6IRQ6Ϡ{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?��?RIAt,1ID`�D�� d1��RQQp�rpDSTB
`� 1�F�HAXD2��|�G�LEXCES?R��ёBMhPa�͠D�BD4�E�q`�`�F_A�J�C[�Ot�H� K��� \��d�bTf$� ��LI�q��SREQUIRE��#MO�\�a�XDESBU��,1L� M�� �p���P�c�DAA$RN��
Q�q�/Ҙ&���-cDC��B�I9N�a?�RSM�Gh�� N#B��N�iPS}T9� � 4��7LOC�RI���;EX�fANG��A^,1ODAQ䵗�@c$��9�ZMF�� ���f��"��%u#��VSUP�' �F�X�@IGGo�� �rq�"��1��#B��$���p%#by��rx����vbPDATA�K�pE;����R��M܋�*� t�`MD
�qI��)�v� �t�A��wH�`��tDIA<E��sANSW��t(h���uD��)�bԣ�(@$`� PCU�_�V6�ʠ�d�PLODr�$`�R���B��B�p�����,1RR}2�E�  ���V�A/A d$C'ALI�@��G~��2��!V��<$R��SW0^D"��A�BC�hD_J2SqE�Q�@�q_J3M�
G�1SP�,��@	PG�n�3m�u�3p�@���JkC���2'AO�)IMk@{BCSKAP^:ܔ9�wܔJy�{BQܜ�����`�_AZ.B��?�ELx��YAOCMP�c|A)��RT�j���c1�ﰈ��@1���t����Z��SMG��pԕ� ER!����INҠACk�@p����b�n _��������D�/R�f�DIU��CDH�@t
�#a�q$V�lFc�$x�$�� �`@���b��̂�E��H �$BE�LP����!ACCE�L���kA°IR�C_R�p@p�T<!�$PS�@B2L�����W3�طx9� ٶPATH���.�γ.�3���p�A_@��_�e�-B�`C�_MG�$D�D��ٰ��$FW��@�p����γ����D}E��PPABN�ROTSPEEu�����O0��DEF�>Q����$USE)_��JPQPC��J�Y����-A 6qYN��@A�L�̐�L�M�OU�NG��|�O9L�y�INCU��a��¢ĻB��ӑ�AENCS���q�B�����D�IN�I�����p�zC�VE�����2�3_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��rPRC����MOS� �gTMOpp�@-GPE�RCH  M�OVӤ �����!3�yD�!e�]�6�<�� ʓA����LIʓdWɗ��p:p3�.�I�TRKӥ�AY����?Q^����m�b��`p�CQ�� MOM�B?R�0u��D����y�0Â��D�UҐZ�S_BCKLSH_C����o� n��TӀ���
c��CLALJ��A8��/PKCHKO0��Su�RTY� �q���M�1�q_
#c�_�UMCP�	C���SsCL���LMTj��_L�0X����E �� �� ���m�`h���6��PC��B��H� �P�ŞCN@�"XT����CN_b��N^C�kCSF����V6����ϡj����nCAT�SH s�����ָ1���֙�0��������PA���_P���_P0� e�`��O1u�$xJG� �P{#�OG���TORQU(�p�a�~�����Ry������"_W ��^�����4t�
5z��
5I;I ;Iz�F��`�!��_8�1��VC"��0�D�B�21�>	P8�?�B�5JRK�<�2��6i�DBL_SMt�Q&BMD`_DLt�&BGRV4
Dt�
Dz��1H_���31�8J�COSEKr�EHLN �0hK�5oDt�jI��jI <1�J�LZ1�5Zc@y���1MYqA�HQBTH|WMYTHET09�NK23z�/Rn�r@[CB4VCBn�CqPASfaYR<4gQt�gQ�4VSBt��R?UGT	S���Cq��a��P#x���Z�C$DUu  ��R䂥э2�Vӑ��9Q�r�f$NE�+p!Is@�|� �$R�#Q�A'UPeYg7EBHBALCPHEE.b�.bS�E �c�E�c�E.b�F�c�j�FR�VrhVghd��lUV�jV�kV�kV�kUV�kV�kV�iHrh@�f�r�m!�x�kH�kUH�kH�kH�kH�i�OclOrhO��nO��jO�kO�kO�kO*�kO�kO�FF.bTQ𰉔E��egSPBA�LANCE��RLmE�PH_'USP���F��F��FPFULC�3��3��E��{1�l�UTO_p ��%T1T2t���2NW�����ǡ��5�P`�擳�T�OU�|��� INSEG���R�REV��R���D3IFH��1���F�1�;�OB��;C���2� �b�4LC�HWAR��i�AB�W!��$MECH`]Q�@k�q��AXk��P��IgU�i�� �
���!����ROBƃ�CR��ͥ�� �C��_s"T �� x $W�EIGHh�9�$�cc�� Ih�.�IF� ќ�LAGK�8S�K��K�BIL?�O1D��U��STŰ�P�; �����������
�Ы�L�� � 2�`�"�DEB�U.�L&�n��PM'MY9��NA#δ�9�$D&���$���� Q   ��DO_�A��� <	���~��L�IBX�P�N��+�_7��L�t�OH  �� %��T���Ѽ�T�����TICK,/�C�T1��%����B��N��c�Ã�R �L�S���S�����PR�OMPh�E� $IR� X�~ ���!�MAI�0��j���_9����t�l�R�0COD��F9U`�+�ID_" =������G_SUFF<0 3�O����DO��ِ��R� �Ǔن�S����!{���ꗰ�	�H)�_FIv��9��ORDX�3 ����36��4X�����GR9�S�.�ZDTD���v��ŧ4 *�L�_NA4���K��DEF_I[�K���g� ��_���i��Ɠ�š���IS`i �萚�D���e����4��0i�Dg����D�� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{ԓ�{� ��{����}��v�� ���g������^�� ��K�Փ����!w�N�P'���^���,`��W\�[R�b��T�EFĨ �O?ULOMB_u��0�VISPIT�Y�A�!OY�A_�FRId��(�SI���R������)3���W�W��0��0_,�EAS %��!�& "����4p�G;� h ���7ƵCOEFF_Om���m�/��G!%�S.�߲CA�5����u�GR` � � $R�4�� �X]�TME�$`R�s�Z�/,)�ER�qT;�:䗰�  ]��LL��S�_S�V�($~�����@���� "SwETU��MEA���Z�x0�u������ g� � �� ȰID�"���!*��&P���*�F�'�� ��)3��#���"��5;`*��REC����!$O�MS�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I��|��MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��|�����zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X17ࡐMO�R�� H	�CU �A3�z�1Q�
��3���$��FVL��2��BbG��� � $SI�@ G�0VO B`נ�OBJE&�!FAD�JU�#EELAYh' ���SD�WOU��p�E1PY���=0Q�T i�0�W�DI�R$ba�pےʠD#YNբHeT�@���R�^�X����OP�WORK}1�,>�SYSBU@p 1�SOP�aR�!�jUĔk�PR��2�ePA`�0�!�cu� 1OP��EUJ��a'�D�Q/IMAG�A	��`fi�IMACrIN,��bsRGOVRD=a�b�0�aP�`sʠ�� �^uz�LP�B��@��!PMC_E(,�Q��N@�M�rǱb��1Ų7�=qSL&��~0���$OVSAL\G*E��*E2y�Ȑ�_=p�w��>p�s ���s	�����B�t�#�}1� @�@;���O&E�RI#A��
N�ЈX�s�f�{��PL�}1�,RTv�m�AT�USRBTRC_T(qR��B �����$� �Ʊ��,�~0� D��`-CSALl`�SA0���]1gqXE���%���C��J�
���cUP(4����PX���؆�q��3�w� ��PG�5� $SUB�������t�JMPWAITXO��s��LOyCFt�!D=�CVF	ь�y�⻑R`�0��CC_�CTR�Q�	�IG�NR_PLt�DB�TBm�P��z�BW�)����0U@���IG��a��Iy�TNLND��Z�R]aK� N��`B�0�PE�s���r���f�SPD}1� L�	�A�`gఠ�S��U!N�{���]�R!�`B�DLY�2����7�PH_PK�E�~�2RETRIEt���2�b���FI�B�� ����8� 2}��0DBGLV�?LOGSIZ$C�KKTؑUy#u�D7�f_�_T1@�EM�@!C\1aA����R��D>�FCHECKK�RS�P�0����@&�f(bLEc�" PA9�QT���P�C߰PN�����ARh�0����Ӯ�PO�BORMATTnaF�f1h�`��2�S��UXy`�	��LB��4� � rEITCH���'7�9PL)�AL_ � $���XPB�q� C,2Dx�!��+2�J3D���� T�pPDCK�yp��oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYL�OA��m�_1t�2<t���J3AR�����դ֏�laTIA4��5��6,2MOM�CP�����������0BϐAD��������PUBk`R��;����;���q��z4�` I$PI\Ds�o�@�1yՕ�w�2�w�Z��I��I��I���p� ���n���y�e`��9S)bT�SPEED� G��(�Е��/��� Е�`/�e�>��M�<�ЕSAMP�6V0��/���ЕMO�@ 2@�A��QP���C�� n�����������LRf`�kb�ІE9h�EIN 09��7S.В9
�yPy�GAMM�%S���D$GE�T)bP�cD]��2
��IB�q�I�G$HI(0;A��LR�EXPA8)LWVM8z)���g���C5�CHKhKp]�0�I_�� h`eT��n�q���eT,���� ��$�� 1�iPI>� RCH_D�313\��30LE�1�1\��o(Y�7 �t�MSW�FL �M��SCRc�7�@�&��%n�f�;SV���PB``�'�!�B�sS_SAaV&0ct5B3NO]�C\�C2^�0�mߗ� uٍa��u���u:e;��1���8��D�P��� ������)��b9���e�GE�3��V��e�Ml�� � F�YL��QNQSRlbfqXG�P�RR�#dCQp� �S:AW70�B�B[�CgR:AMxP�KCL�H���W$�r�(1n�g�M�!o��� �F�P@}t$WP�u�P r��P5� R<�RC�R��%�6@�`��� ��qsr X��	OD�qZ�Ug�ڐ>D�� ��OM# w�J?\?n?�?�?��9��b"�e�]�_��� |��X0��bf�Ӏqf��q`�ڏgzf��E�ڐ��Ec�"�5�t��FdPB��PM��QU�� � 8�L�QCOU!5�Q�THI�HOQBpH�YSY�ES��qU�E�`�"�O��� � �P�@\�UN����Cf�O�� P��Vu��!����OOGRAƁcB2�O�tVuITe �q:p/INFO�����{��qcB�e�OI�r�{ (�@SLEQS� �q��p�vgqS����� 4L�ENA�BDRZ�PTION�t�����Q���)�GCuF��G�$J�,q^r�� R���pU�g�����_ED��N��� �F��PK��j��E'NU߇�وAUT$1܅CO�PY�����n�00M�N���PRU�T8R �Nx�OU���$G[rf�|���PRGADJ���f*�X_:@բ$��(���P��W��P��} ���)�}�EX�YmCDR}�NS.�9�F@r�LGO�#��NYQ_FREQ�R�W� �#�h�TsL�Ae#����ӄ �CcRE� s�IF�ᶕsNA��%a�_}Ge#STATUI`<e#MAIL������q t�������EwLEM�� �/0><�FEASI?�B ��n�ڢ�vA�]� � I�p��Y!q]�Lt#A�ABM���E�pr<�VΡY�BASR҈Z��S�UZ��0�$q���RMS_TR;�qb ���SY��	�ǡ��$���>C��Q`	� 2� _�TM������̲��@ �A��)ǅ�i$D�OU�s]$Nj���P�R+@3���rGRIyD�qM�BARS �sTY@�|�OTO�Rp��� Hp_}�!����d�O�P/�� �s �p�`POR�s���}���SRV��),����DI&0T��Ѡ�� #�	�#�4!�5*!�6!�7!�8�e��F�2��Ep$VALUt��%��ֱ��>/��� ;�1ėq�����(_�AN��#�ғ�Rɀ(���T�OTAL��S��P�W�Il��REG#EN�1�cX��ks0(��a���`TR��R��_S� ��1ଃV �����⹂Z�E��p��q��Vr���V_Hƍ�DA�S����S_�Y,1�R4�S� AR��P2� ^�IG�_SE	s����å_�Zp��C_�Ƃ�EN�HANC�a� T ;�������GINT�.��@FPs^İ_OVRsP�`@p�`��Lv��o��7�p}��Z�@�SLG�
AA�~�25�	��Dd��S�BĤDE�1U�����TE�P���� !Y��
��J��$2�IL_M`C�x r#_��`TQ�`���q���'�BV�CF�P_� 0�M�	[V1�
V1�2�U2�3�3�4�4�
�!���� � m�A�2IN~VIB�P���1�2�2��3�3�4�4��A@-�C2���=p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KEEP_HNADD!�!`$^�j)C�Q�� �$��"	��#O�a_$�A�!�0�#i��#REM�"�$��½%�!��(U}�e�$HPW�D  `#SBWMSK|)G�qU�2:�P	�COLLAB� �!K5�B�� 4��g��pITI1{�9p#>D� ,�@F�LAP��$SYNT �<M�`C6���UP_DLYAA�ErDELA�0ᐢ�Y�`AD�Qz�QSwKIP=E� ���XpOfPNTv�A�0P_Xp�rG�p�RU@ ,G��:I+�:IB1:IG� 9JT�9Ja�9Jn�9J{к9J9<��RA=s� X���4�%1�Q}B� NFLIC�s��@J�U�H�LwNO�_H�0�"?��RIT�g��@_PA�pG��Q� ��^�U�W��LV�d�NGRLT�0_q��O�  p" ��OS��T_JvA� V	�APPR_W�EIGH�sJ4CH?pvTOR��vT���LOO��]�+�tVJ�е�ғA�Q�U�S�X�OB'�'���J2TP���7�X�T� <a43DP=`Ԡ\"<a�q�\!��RDC��L�+ �рR��R�`� ��RV��jr�b�R�GE��*��cN�FL�G�a�Z���SPC��s�UM_<`^2�TH2NH��P.a �1� m`EFv11��� lQ `�!#� <�p3AT�  g�S�&�Vr�p�tMq�Lr���HOME(wry�t2'r�-?�Qcu��w3'r逪������w4'r�'�9�K�]�o���
�w5'r뤏��ȏڏ(����w6'r�!�3��E�W�i�{���7'r퀞���ԟ�����8'r��-�?�Q�c�u�R��S$0�q�p��� sF��`�1�"`P������`/���-�I�O[M�I֠�Ћ�qPOWE�� ��0Za�0p��� �5��$DS=B GNAL���0�Cp��m`S232N3�� �~`��� �/ ICEQP��PE�p��5PIT����O�PBx0��FLOW�@TRvP��!U����CU�M��UXT��A��w�ERFACt�� U��ɲ;CH��� tQ  1_��>�Q$����SOM��A�`T�P.#UPD7 A�ct�T��UEX@�ȟÎU EFA: X"�1RsSPT�����T 
��PPA�0o񩩕`EXP�IOS���)ԭ�_���%��C�#WR�A��ѩD�ag���`ԦFRIEND�saC2UF7P����TwOOL��MYH �C2LENGTH_VTE��I��Ӆ�$SE����UFOINV_����RGI�{QITI�5B��Xv��-�G2-�G17�w�SG�X�"��_��UQQD=#�� �AS��d~C�`��|q�� �$$C/�=S�`�����S0�S0 ��VERsSI� �����5��I��������AAVM_Y�2� � �0  �5���C�O�@�r� r�	 ����S0�!����������������
?QY�B�S���1��� <-�� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O�OiCC�@XLM�T&����  ���DIN�O�A�Dq�EKXE�HPV_���ATQz
��LA�RMRECOV ��RgLMD/G *�5�O�LM_IF *��`d�O�_�_�_�_�j�_'o9oKo]onm, 
��odb��o��o�o�o^��$� <z, A   2D{��PPINFO u[ �Vw��������`�� �����*��&�`�@J���n�����DQ� ���
��.�@�R�d��v���������a
PP�LICAT��?��P��`�Handling�Tool 
� �
V8.30P/�40Cpɔ_LI�
883��ɕ$?ME
F0G�4��-
398��ɘ�%�z�
7DC3�ɜ
��NoneɘVr�|��ɞ@6d�� Vq_ACTI�VU��C죴�M�ODP���C�I��HGAPON���n��OUP�1*�� i�m����Қ�_����1*�  �@�������� Q���Կ�@�
������ ����5�Hʵl�K�?HTTHKY_�� /�M�SϹ�������� �%�7ߑ�[�m�ߝ� �ߵ����������!� 3��W�i�{���� ����������/��� S�e�w����������� ����+�Oa s������� '�K]o� �������/ #/}/G/Y/k/�/�/�/ �/�/�/�/�/??y? C?U?g?�?�?�?�?�? �?�?�?	OOuO?OQO cO�O�O�O�O�O�O�O �O__q_;_M___}_ �_�_�_�_�_�_kŭ��TOp��
�DO_CLEAN9��pc_NM  !{血�o�o�o�o�o��D?SPDRYRwo��HI��m@�or� ��������p&�8�J���MAXݐ Wdak�H�h�XWd��d���PLUGGpW�Xgd��PRC)pB�`�kaS��Oǂ2DtSEGF0�K� �+��o�or�����������%�LAPOb�x�� �2�D� V�h�z�������¯ԯ|�+�TOTAL��|��+�USENUO��\� e�A�k­�R�GDISPMMC�.���C6�z�@@$Dr\�OMpo�:�X��_STRING �1	(�
��M!�S�
��_�ITEM1Ƕ  n������+�=� O�a�sυϗϩϻ����������'�9��I/O SIGN�AL��Try�out Mode�ȵInpy�Simulateḏ�Out��O�VERRLp = �100˲In �cycl�̱P�rog Abor���̱u�Stat�usʳ	Hear�tbeatƷM?H Faul	��Aler�L�:�L� ^�p��������� ScûSaտ�� -�?�Q�c�u������� ��������);pM_q��WOR.� û������ +=Oas�� �����//'.PO����M �6/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~?��?�?�?�?H"DEV P.�0d/�?O*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_PALT	��Q� o_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o��o�o�o�_GRI m�û9q�_as� �������� '�9�K�]�o�������'�R	�݁Q��� �)�;�M�_�q����� ����˟ݟ���%�x7�I�ˏPREG�^ ����[�����ͯ߯� ��'�9�K�]�o����������ɿۿ�O���$ARG_� D �?	���0���  w	$O�	[D��]D��O�e�#�SB�N_CONFIG� 
0˃����}�CII_SAV/E  O������#�TCELLSE�TUP 0�%�  OME_IO�O�O�%MOV_qH������REP���J��UTOBAC�K�����FRA:\o� �Q�o���'`���o���� �� f�o�����*�!�83�`�Ԉ��f�� ���������o�{�� &�8�J�\�n������ ������������"4 FXj|�������끁  ���_i�_\ATB�CKCTL.TM�P 6.VD GIF ��BN`r<�o�N�R��fЗINI�P�Օ�~c�MESSAG�����8��ODE_!D����z��O�0��c�PAUSM!!�~0� (73�U/g+(Od/�/x/ �/�/�/�/�/�/??�?P?>?t?1�0$: TSK  @-��Tߞf�UPDT��d��0
&XWZD_�ENB����6ST�A�0��5"�XIS~��UNT 20���� � 	 �� $� 1����q�TŵӀ��$Gİ2�H����zF��Oo�}Cw�g�^����.�O�O�O��O/_2FMET߀2�CMPTAA Q�@ԑ�A���@���@���@���rK5���5�(d5��P�5�r�5F*�5�338]SCR�DCFG 1�6/�Ь�Ź�_�_oo(o:oLo��o�Q���_�o�o�o �o�o�o]o�o>P bt���o9�iуGR<@M/�s/N5A�/�	i��v�_ED�1�Y� 
 �%-5�EDT-�'�G?ETDATAU�o��9�u?�j�H�o��f�\��A��  ���2�&�!�E���:IB���~�ŏ׏m����3��&۔� �D��ߟJ�����9�ǟ�4���ϯ�(�����]�o�����5 N������(�w��)�;�ѿ_��6ϊ�g� ��(�CϮ���ϝ�+��7��V�3�z�(��@z�����i����8��&���~�]���F����5����9~������]����Y�k�����CR�!ߖ��� W�q���#�5���Y��p~$�NO_DEL���rGE_UNUS�E��tIGALL_OW 1���(*SYST�EM*S	$S?ERV_GR�Vܖ : REG�$8�\� NUM�
���PMUB U�LAYNP\?PMPAL��CYC10#6x $\ULSU0�8:!�Lr��BOXORI�C�UR_��PM�CNV�1�0L�T4DLI�0��	����BN/ `/r/�/�/�/�/�/����pLAL_OUT� �;���qWD_ABOR=f�q�;0ITR_RTN��7�o	;0NONS�0�6 
HCCF�S_UTIL 9#<�5CC_@6Aw 2#; h ?��?�?O#O6]CE_�OPTIOc8�qF@RIA_I�c f5Y@�2�0FF�Q�=2q&}�Ao_LIM�2.�� ��P�]B�T�KX�P
�P�2O��Q��B�r�qF�PQ5T1)TR�H��_:JF_PARAMGP 1�<g^&S�_�_�_�_~�VC�  C�dE�`�o!o`�`U�`�`�Cd��T@ii:a:e>eBa�Gg�C�`� D� kD	�`�w?��2{HE ONFI� �E?�aG_P�1#; ���o�1CUgy�aKoPAUS�1�yC ,����� ����	�C�-�g� Q�w���������я���rO�A�O�H��LLECT_�B�IPV6�EN. QF�n3�NDE>� �G��71234?567890��sB�TR����%
 H�/%)������� W���0�B���f�x��� 㯮���ү+����� s�>�P�b��������� �ο��K��(�:�Г�^�|��B!F� ��I|�IO #��<U%e6�'�9�lK���TR�P2$���(9X�t�Y޼`%��̓ڥH��_MOR֮3&�=��@XB��a��A�$� �H�6�l�~���~S��'�=�r_A?�a�a`D��@K��R�dP��y)F�ha�-�_�'�9�%
�k��G�� ��%Z�%���`�@c.�PDB�+���cpmidbg��	�`�:�  2-' .�QU��p��N g ��@�0i/����]܌0���0�Az<�^�*�@x�@ywg�$V��`@�wf�l�q��ud1�:��:J��DEFg *ۈ��)��c�buf.tx�t����_L64FIX ,�� ����l/[Y/�/}/�/ �/�/�/
?�/.?@?? d?v?U?�?�?�?�?�?��?,/>#_E -���<2ODOVOhOzO��O6&IM��.o�YU>���d�
�I�MC��2/����dXU�C��20�M�QT|:Uw�Cz  B��i�A���A����Au�gB3��*CG�B<��=w�i�B.��B����B��5B��$�D�%B���ezVC�q��C�v�D����D-lE\D�n �hw��29"6��22o�D|���U�� ���C5�C����
��h�D4cdv`D��`/�`v`s]E�D� D�` E4��F*� Ec���FC��u[F����E��fE���fFކ3FY_�F�P3�Z��@��33 ;��>�L���Aw�n,a@:��@e�5Y���a����`A��w�=�`<#���
��?�ozJ�RSMOFST c(�,bIT1��eD @3��
д���,�a��;��bw�?���<�M^�NTEST�1O��CR@�4��>VCF5`A�w�Ia�a�ORI`CTPB�U�C��`4���r��:Sd����qI?�5���qT_�PRO'G ��
�%$/ˏ��t��NUSER � �U������KE�Y_TBL  �����#a��	
��� !"#$%�&'()*+,-�./��:;<=>�?@ABC�GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~��������������������������������������������������������������������������������͓���������������������������������耇��������������������������LCK��
����STAT�/��s_AUTO_�DO �	�c�INDT_ENBP�b��Rpqn�`�T2�����STOr`���X�C�� 26���8�
SONY XOC-56�"b�����@��F( ����HR50�w���>�P�7b�t�A�ff����ֿ�  Ŀ����C�U�0�y� ��fϯ��Ϝ������ϸ�-ߜ�TRL��L�ETEͦ ��T�_SCREEN ���kcs����U�MMEN�U 17�� <ܹ���w������ ����K�"�4��X� j������������ 5���k�B�T�z��� ������������ .g>P�t�� ����Q( :�^p���� /��;//$/J/�/ Z/l/�/�/�/�/�/�/ �/7?? ?m?D?V?�? z?�?�?�?�?�?!O�? 
OWO.O@OfO�OvO�O��O(y��REG 18�y����`�M�����_MANUAL��k�DBCO��R�IGY�9�DBG_oERRL��9��q��_�_�_ >^QNUMLI�pϡ��pd
�
^QPXWORK 1:���_5oGoYoko}oӍ�DBTB_N� �;������ADB_AWAYzfS�qGCP 
�9=�p�f_AL�pR���bbRY�[�
�WX_��P 1<{y�n�,��%oc�P��h_MM��ISO��k@L���sONTIMX�M�
���vy
���2sMOTNEND��1tRECORDw 1B�� ���sG�O�]�K��{ �b��������V�Ǐ� ]����6�H�Z��� ������#�؟���� ��2���V�şz����� ���ԯC���g��.� @�R���v�寚�	��� п���c�χ�#ϫ� `�rτϖ�Ϻ�)ϳ� M���&�8ߧ�\�G�8Uߒ��8����߀��K� �����6��%RC7�n���ߤ��8�����A�4����$���H�3�A�~��;�������9���]�8�����|�B#Z�l���zTOLER3EN\�rB�'r�`�L��^PCSS_�CCSCB 3C>y�`IP��}�~� <�_`r�K������/�{� �5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O��O_�~�LL� D���fFY C[C��PZP^�r_ A� p� ��sp��Q �\	� A�p�Q�_�[?� �_�[oU�p1�P�pSB�V�c �(a�PWoio{h+�o��X�o�oY��[	r�hLP����ޮ?�����:�3߮|��c��aD@�VB��|�G����+��K� �otGhXGr��So����eB   =��Ͷa�>�tYB�� �pC(�p�q�aA"�H�S�Q -��q���ud�v���|��AfP ` 0����D^P��p@�a
�QX��\� aW>� �a9P� �b�e:�L�^�h�Hc�́PQ�R�Q�PU�z �֟�o\^��-�?���c�u����zCz�ů�b2�Щ�_ ����S̡0��]�0� .�����.a��F� X�ѿUҁп�VS���NSTCY 1	E��]�@rIϫ� K�]�oρϓϥϷ��� �������#�5�G�Y��k�}ߏߒ��DEV�ICE 1F5� E_����	� ��?�6�c��V|㰟�����_HNDGD �G5�VP���R�LS 2H�ݠ��/��A�S�e�w����� ZPARAM I��FgHe�RBT [2K��8р<�߬WPpC�{��,`¢�P�Z�z��%>{�C*  �2�j�MTv�,`"nPB , s��M� }�gT�g��
B��!�bcy�[2Dch z����/���/gT#I%D��CǓ` b!�R��A���A,��Bd���A�;���_C14kP�!2�C��$Ɓ��]�ffA�À���B�� �| �0��/�/�T (��5 4a5�}%/7/d?/ M?_?q?�?�?�?�?�? O�?OO%O7OIO�O mOO�O�O�O�O�O�O �OJ_!_3_�_�_3�_ �_�_�_�_o�_(oo Lo^oЁ=?k_IoS_�o �o�o�o�o�o�o #5G�k}�� �����H��1� ~�U�g�y�ƏAo�Տ ���2�D�/�h�S��� go����ԟ����ϟ� ��R�)�;���_�q� ���������ݯ�<� �%�7�I�[�m����� ����}�&��J�5� n�YϒϤϏ��ϣ�ѿ ������F��/�A� ��e�w��ߛ߭����� ����B��+�x�O�a� �����������,� ��%�b�M���q����� ����������L #5�Yk}�� � ��61 CUg����� ���	//h/���/ w/�/�/�/�/�/
?�/ .?@?I/[/1/_?q? �?�?�?�?�?�?�?O O%OrOIO[O�OO�O �O�O�O�O&_�O_\_ 3_E_W_�_?�_�_�_ �_�_"ooFo1ojoE? s_�_�om_�o�o�o�o �o0f=Oa �������� ��b�9�K���o��� Ώ��[o��(��L��7�I���m������$�DCSS_SLA�VE L��}�ё���_4D  љ�~�CFG Mѕ���������FRA:\ĐL�-�%04d.CS�V��  }�� ����A i�CHq�z������|�����"������Ρޯ̩硞Ґ-��*����_�CRC_OUT �N������_�FSI ?њ ����k�}� ������ſ׿ ���� �H�C�U�gϐϋϝ� ���������� ��-� ?�h�c�u߇߽߰߫� ��������@�;�M� _����������� ����%�7�`�[�m� ��������������� 83EW�{� ����� /XSew��� ����/0/+/=/ O/x/s/�/�/�/�/�/ �/???'?P?K?]? o?�?�?�?�?�?�?�? �?(O#O5OGOpOkO}O �O�O�O�O�O _�O_ _H_C_U_g_�_�_�_ �_�_�_�_�_ oo-o ?ohocouo�o�o�o�o �o�o�o@;M _������� ���%�7�`�[�m� �������Ǐ����� �8�3�E�W���{��� ��ȟß՟���� /�X�S�e�w������� �������0�+�=� O�x�s���������Ϳ ߿���'�P�K�]� oϘϓϥϷ������� ��(�#�5�G�p�k�}� �߸߳����� ���� �H�C�U�g���� ���������� ��-� ?�h�c�u��������� ������@;M _������� �%7`[m ������� /8/3/E/W/�/{/�/ �/�/�/�/�/??? /?X?S?e?w?�?�?�? �?�?�?�?O0O+O=O OOxOsO�O�O�O�O�C��$DCS_C_�FSO ?�����A P �O�O_?_ :_L_^_�_�_�_�_�_ �_�_�_oo$o6o_o Zolo~o�o�o�o�o�o �o�o72DV z������� 
��.�W�R�d�v��� ����������/� *�<�N�w�r������� ��̟ޟ���&�O� J�\�n���������߯ گ���'�"�4�F�o� j�|�������Ŀֿ�������G�B�T��OC/_RPI�N_j� �����ς��O����1�XZ�U��NSL��@&� h߱���������"�� /�A�j�e�w���� ����������B�=� O�a������������� ����'9b] o������� �:5GY�} ������// /1/Z/U/g/y/�/�/ �/�/�/�/�/	?2?-? ??Q?z?u?��ߤ߆? �?�?�?OO@O;OMO _O�O�O�O�O�O�O�O �O__%_7_`_[_m_ _�_�_�_�_�_�_�_ o8o3oEoWo�o{o�o �o�o�o�o�o /XSew��� �����0�+�=� O�x�s���������͏ ߏ���'�P�K�]��o����� �PRE_?CHK P۪��A ��,8��2��� 	 18�9�K���+�q� ��a�������ݯ�ͯ �%��I�[�9���� o���ǿ��׿���)� 3�E��i�{�Yϟϱ� ������������-� S�1�c߉�g�y߿��� �����!�+�=���a� s�Q�������� ������K�]�;��� ��q������������� #5�Ak{� ����� CU3y�i�� ����/-/G/ c/u/S/�/�/�/�/�/ �/??�/;?M?+?q? �?a?�?�?�?�?�?�? �?%O?/Q/[OmOO�O �O�O�O�O�O�O_�O 3_E_#_U_{_Y_�_�_ �_�_�_�_�_o/oo SoeoGO�o�o=o�o�o �o�o�o=- s�c����� ��'��K�]�woi� ��5���ɏ������� �5�G�%�k�}�[��� ����ן�ǟ���� C�U�o�A�����{��� ӯ����	��-�?�� c�u�S�������Ͽ� ������'�M�+�=� �ϕ�w�����m���� ��%�7��[�m�K�}� �߁߳��߷����!� ��E�W�5�{��ϱ� ��e�������	�/�� ?�e�C�U��������� ������=O- s����]�� ��'9]oM �������/ �5/G/%/k/}/[/�/ �/��/�/�/�/?1? ?U?g?E?�?�?{?�? �?�?�?	O�?O?OO OOuOSOeO�O�O�/�O �O�O_)__M___=_ �_�_s_�_�_�_�_o �_�_7oIo'omoo]o �o�o�O�o�o�o! �o1W5g�k} ������/�A� �e�w�U�������я ��o����	�O�a� ?�����u���͟��� ��'�9��]�o�M� ��������ۯ��ǯ� #�ůG�Y�7�}���m� ��ſ�����ٿ�1� �A�g�E�wϝ�{ύ� ������	�߽�?�Q� /�u߇�e߽߫ߛ��� �����)���_�q� O���������� ���7�I���Y��]� ��������������! 3WiG��} ����%�A �1w�g��� ���/+/	/O/a/ ?/�/�/u/�/�/�/�/ ?�/9?K?�/o?�? _?�?�?�?�?�?�?O #OOGOYO7OiO�OmO �O�O�O�O�O_�O1_ C_%?g_y__�_�_�_ �_�_�_�_o�_+oQo /oAo�o�owo�o�o�o �o�o);U__q ������� �%��I�[�9���� o���Ǐ�����ۏ!� 3�M?�i��Y����� ��՟�ş����A� S�1�w���g�����������ӯ�+�=��$�DCS_SGN �QK�c��7m�� 16-M�AY-19 10?:20   O�l��4-JANt�08�:38}�����? N.DѤ�����������M4�o���Im��P��Z�q��  O�V�ERSION �[�V3.5�.13�EFLO�GIC 1RK���  	���P�?�P�N�!��PROG_ENB  ��6Ù�o�ULSE  T����!�_ACCL{IM���������WRSTJN�T��c��K�EM�Ox̘��� ���INIT S.�G�Z����OPT_SL �?	,��
 	�R575��Y�7�4^�6_�7_�50
��1��2_�@ȭ��><�TO  Hݷ�t��V�DEX���dc����PAT�H A[�A\��g�y��HCP_�CLNTID ?<��6� @ȸ�����IAG_GR�P 2XK�? ,`��� � �9�$�]�H������123456�7890����S�� |�������!�� ��H���;� dC�S���6� ����.�R v�f��H� �//�</N/�"/ p/�/t/�/�/V/h/�/ ?&??J?\?�/l?B? �?�?�?�?�?v?O�? 4OFO$OjO|OOE� �Oy��O�O_�O2_��@_T_y_d_�_,
�B^ 4�_�_~_`Oo �O&oLo^oI��Tjo�o .o�o�o�o�o �O' �_K6H�l�� �����#��G��2�k�V���B]�?g��?����>�����*��{��V>h)>���ž4	��d��D��?��?ihD=P���� �����(��L�B\ډ�C*����U{���>���:������ߟʟܟ���CT�_CONFIG �Y��Ӛ��egU���STB_F_TTS��
�ɠb����Û�u�O�M�AU��|��MSW�_CF6�Z��  ��OCVIEWf��[ɭ����� �-�?�Q�c�u�G�	� ����¿Կ������ .�@�R�d�v�ϚϬ� ��������ߕ�*�<� N�`�r߄�ߨߺ��� ������&�8�J�\� n���!�������� �����4�F�X�j�|�,���RC£\�e��!*�B^�������C2g{�SBL_�FAULT ]���ި�GPMSK�k��*�TDIAG' ^:�աI���UD1: 6�78901234!5�G�BSP�- ?Qcu���� ���//)/;/M/tJ��
@q��/>$�TRECP��

��/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOi/�{/xO�/UMP_OPTIONk���A�TR¢l��	�EP�MEj��OY_TE�M�È�3B��J�P�AP�DU�NI��m�Q��YN_BRK _ɩ��EMGDI_S�TA"U�aQK�XPN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 J�#q��,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;��������� ��!� ��~��������[F�EATURE �fj5��JQ�Handling�Tool � "�
PEng�lish Dictionary��def.4Dw St�ard��  
! h�Analog I�/OI�  !
�IX�gle Sh�iftI�d�X�u�to Softw�are Update  rt s����matic B�ackup�3\�st��gro�und Edit���fd
�Camera`�F�d�e��CnrRn�dIm���3�C�ommon ca�lib UI�� /Ethe�n��"�Monitor�oLOAD8�tr�?Reliaby�O��ENS�Data ?Acquis>���m.fdp�iag�nos��]�i�Do�cument V�ieweJ��87�0p�ual C�heck Saf7ety*� cy� ��hanced U�s��Fr����C� �xt. DIOm :�fi�� m8����end��Err�I�L��S������s�  t Pa�r�[�� ���J94�4FCTN /Menu��ve�M�� J9l�TP I�nT�fac{�  �744��G��p �Mask Excz��g�� R85��T��Proxy �Sv��  15 �J�igh-Sp�e��Ski
� R�738Г��mm�unic��ons��S R7��ur8r�T�d�022��a����connect� 2� J5��I�ncr��stru�,Қ�2 RK�AREL Cmd�. L��ua��R�860hRun-�Ti��EnvL�o�a��KU�el +:��s��S/Wѹ��7�License����rodu� o�gBook(Sy�stem)�AD� pMACR�Os,��/Off�s��2�NDs�MH��� ����MM�RC�?��ORDE�� echStopr��t? � 84fcMi$�|� 13d�x��]е�׏���M�odz�witchBI�VP��?��.� sv��2Opt�m�8�2��filз�I ��2g 4� !+ulti-�T�����;�P?CM funY��Po|���4$�b&R�egi� r �P�ri��FK+7���g� Num Sel�W  F�#�� �Adju���60q.��%|� fe�ў�&tatu�!$6����%��  9 J�6RDM R�obot)�sco{ve2� 561��RemU�n@� �8 (S�F3Ser�vo�ҩ�)SNPX b��I�\dcs�0}�L�ibr1��H�� �5� f�0��5�8��So� tr�s�sag4%G 91E�p ��&0����p/I��  (i~g TMILIB(M<Ӌ�Firm�����gd7���s�Accd����0�XATXN�Heln��*LR"1x��Spac�A�rquz�imul�aH��� Q���To�u�Pa��I��T���c��&��ev.� f.svU�SB po��"�iuP�a��  r"1�Unexcept���`0i$/����H5-9� VC&�r��[6���P{��RcJP�RIN�V�; d �T@�TSP CS�UI�� r�[XC���#Web Pl6�%d -c�1�R�@4d�����I�R�66?0FV�L�!FVG�ridK1play C�lh@����5R�iR�R.@���R-�35iA���Ascii���"���� 51f�cUpl�� � (T����S���@rityAv�oidM �`��C�E��rk�CoYl%�@�GuF� 5P��j}P����
 B�L�t� 120C C�� o�І!J��P��yH��� o=q�b @oDCS b ./��c��O��q��`�; ����qckpaboE4�DH@�OTШ�?main N��19.�H��an.��A:> aB!FRLM����!i ���MI D�ev�  (�1� #h8j��spiJP�� � �@��Ae1/�r����!hP� M-2 � i��߂^0i�p�6�PC��  i�A/'�Passw�o�qT�ROS �4����qeda�SN��Cli����Gr6x Ar�� 47�!t���5s�DER��.�Tsup>Rt�I��7 (M�a�T2D�V�
�3D Tr�i-���&��_8t;�
�A�@Def?�����Ba: deRe p 4t0�Пe�+�V�st64MB DRAM��h86΢FRO�֫0�Arc� vi�sI�ԙ�n��7| �), �b�Hea�l�wJ�\h��Ce�ll`��p� �sAh[��� Kqw�c�G - �v���p	V,Cv�tyy�s�"�/�6�ut��v�m���xs ���T�D_0��J�m�` 2���a[�>R tsi��MAILYk�/�F2�h��ࠛ 90C H��F02]�q�P5'���T1C��5��F��FC��U�F9�OGigEH�S�t�0/A� if�!2���boF�dri=c ^�OLF�S�����" H5k�OP3T ��49f8���cro6��@ꊠl�ApA�Syn�.(RSS) 1�L�\1y�rH�L� (`2x5�5�d�pCVx9\����est�$SРl��> \pϐSSF��e$�tex�D o@���A�	� BP����a�(R00�Qirt��:���2)�D��1��e�VKb@l B�ui, n��WAP!Lf��0��Va�kTF�XCGM��D��L����[CRG&a�YBU��YKfL��p�f��k�\sm�ZT�Af�@�О�Bf2��и��V#�s���� r���CB���
f(���WE��!��
����T�p��DT��&4 Y�V�`��EaH����
�61Z���
�R=2�
�E (Np��F�V�PK�B��D�#��Gf1`?G����H�р?I�e �����LD�L��N��7\s@���`�z��M��dela<,���2�M�� "L[P��`?��_�%������S��-F�T�SO�W�J57η�VGF�|�VP2֥ 5\b�`0&@�cV:���T;T� ܨ<�ce,?VP�D��$T;F���DI)�<I�a\so<��a-�6Jc6As6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P�
� ����`��Im'g PH�[l���I/A  VP�S��U�Ow��!%S�S>kastdpn)ǲt��� SWIMES5T�BFe�00��-Q�� �_�PB�_�Ru#ed�_�T�!�_�Sx ��_bH573ob2c2��-oNbJ5N�HIojb)�Cdo�cxE� �o�_�lp��o�TdP�o �c�B�or�2.rٱ`(Jsp�EfrSEop�f1�}�r3 RGoNeELS��sL�� ��s�����B	��S�\ $�F�ryz�ft	l�o~�g�o�����@����?�����P  �n�&�"�l ��T�@�<�^��Y��e�u8<Z���alib��Γ���ɟ3���埿�\v� ��e\c�6�Z�f8�T�v�R VW���98S��UJ91�����i�ů[c91+o�w8<���847�:� �A4�j��Q��t6�m���vrc.����HR���ot�0ݿ��'  ��8ޯ�3460�>eS0L��97���U�ЄϦ�60.� g�н�+��'��ܠ�Ϻ�8co��DM�߱U"�����ߕpì߲T! ��na;�� ���u%�����I��loR�d��1a59gϱŭ���95�ϔ�R����1 ��?��o�#��1A�/�d��vt{�UWeǟ����ￇ73[���7��ρ�C W��6I2K�=fR���8��@������d����2��ڔ����@�@"< "http������t7 �� v R7��78����p4�� ��TTPT�p#	��ePCV4/dv߀�j�Q�Fa7�b�$N�0�/2�rIO�p)/;/M/6.sv3��64i�oS�l? to�rah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��O�B4c.K?�g'�)�294g?�� (B�Ofd�\iOA5sb�?U_�?vi�/i��/�/BWn��`�o%�Fo��4l�$of��oXF sI)xo�cmp\7f��mp���duC��0lh����o(A�_Bt� �o]6P��m�I?�w��@���naO��4*O0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե1�1?o��DMs�B	C��7J�\���(�952�XFa AP�ڟ�<�v�`/şaqs8����/Of��I1�9�VRK�0��ph�քH5+�=�sIN/¤SkiW�/�IF��_�%�F�fs�I�O�l����"<𜿚$�`�����\jԿz5bO�vro�uς�3(�ΤH (DϮ��?sG��|��F �Ou�������D)O��*�3P$�FӅ�k���ϻ���럴� �PLx��ʿ��pbox��f�ebo���Sh �>�R.�0wT{����fx6��P��D��03��#_I\m;YE	e�OԆM�hxW�=E�te,���dct\���O$kR�����2�Xm*���ro3��D�l�j9��V<'�  FC����|@�ք f?6KA�RE0�_�~ (Kh��.cf���WcpoO�_K�up���a���H/j#- E�qd/�84���$qu�o��/ o2o?Vo"<�7C�)�s�NJԆx�|?�3l\sy�?0�40�?Τwio�u�]?�w58�?,F�0$OJ�
?Ԇ"io�!��V��u&A��PR��ߩ5, s��v1\�  H5352B�Q21p0�R78P51�0.R0  ne�l J614�Ҡ/WAT�UP��d8P545�*�H8R6��9�VCAM�q97PC�RImP\1tPUIF��C8Q28  in�gsQy0��4P P63rP @P PSCH��?DOCVڀD ��PCSU���08Q0�=PqpVEIO�Cr��� P54Pu;pd�PR69aP����PSET�pt\h�PQ`Qt�8P7`Q�!�MASK��(P�PRXY���R7�B#POCO  \pppb36���PR �Q��b1Pd60Q$c/J539.eHsb��?vLCH-`(��OPLGq\�bPQ0]`��P(`H�CR��4`S�au;nd�PMCSIP`e)0aPle5=Ps�p(`DSW� �  qPb0`0�aPa��(`PRQ`Tq0�RE`(Poa601P<cgPCM�PHcR0@q\j23b�V�`E`8�S`UPvisP`�E` c�`UPcPRS�	a�bJ69E`sF�RDmPsRMCN�:eH931PHcSNsBARa�rHLB�U�SM�qc�Pg52΁fHTCIP0cTMCIL�e"P�`eJ ��PA�PdSTPTXv6p967PTEL�p@��P�`�`
Q8P8$Q�48>a"PPX�8P915�P`[�95qqbwUEC-`F
PGUFRmPfahQCmP;90ZQVCO�`@�PVIP%�537nsQSUIzVSX�P��SWEBIP�SHT�TIPthrQ62�aP�!tPG���cIGt؁�`c�PGS�e�IRC%��cH76D�P�e Q�Q|�Ror��R51P s:P�P&,t53=P8u8=Py�C�Q6]`�b�PI��q52]`sJ56`E`s���PDsCL�q�Pt5�\rd�q7�5UP cR8���u5P sR55]`,s�  P8s��P�`CP�PP��SJ77P0\o��6��cRPP�cR�6�ap�`�QtaT�7�9P`�64�Pd87]`�d90P0c���=P,���5�9ta�T91P� ��1P(S��n�Qpai�P06=PW- C�PF�T	�0��!aLP PTS�pL��CAB%�I БI�Q` ;�H�UPPai-ntPMS�Pa��D��IP|�STY%�t\patPTO�b�P��PLSR76�`�5ؐQ��WaNN�Pai�c�qNNE`�OR�S�`�cR681Pi;nt'�FCB�P(��6x�-W`M�r��!�(`OBQ`plug��`L�aot �`O#PI-���PSPZ��PPG�Q7�`73nΒPRQadRL��(Sp�PSⳲn�@�E`��� �PTS-�� 8W��P�`apw�`���P`cFVR�PlcVs3D%�l�PBVI��SAPL�Pcycn+PAPV1�pa_��CCGIP - U���L�Prog+PC�CR�`�ԁB�P 4�PԁK=�"L�P��$p��(h�<�P��h��̱�@g�Bـ
TqX�%���CTC�p�tp��2��P927�"0ҝPs2�Qb��T�C-�rmt;�	`#�1ΒTC9`HcCT�E�Perj�EIPp.p/�E�P�c��I��use��Fـvr2v�F%���TG�P� �CP��%�d -h�H�-�Tra�PCTI��p��TL� TRS���p�@נ��IP�PuTh�M%�lexsQ{TMQ`ver, �p�SC:���F��Pv�\e�PF�IPSV"`+�H�$cj�ـtr�a�CTW-���CPVG�F-��SVP2mPv'\fx���pc�b���e��bVP4�fx_qm��-��SVPD-���SVPF�P_moҟ`V� cV��t\z��LmPove4��\-�sVPR�\|�tPV�Qe5.W`V 6�*u"��P}�o`���`N��CVK��N�IIP��CV����IPN9�Gene���D�@�D�R�D����  ��yf谔�pos.��/inal��n��D"eR���`��d�P��somB���on,��иR�D�R��\��TXpf��D$b��omp��G "N��P��m����! ��=C-f8����=FXU�����g F��(��Dt� II��r�D��u��� "����Cx_�ui X������fa2��h	Crl2��D,r9ui�Ԣ�� it2c�0c�o��e"�����ާ(.)� ��{�� ��� �IQnQ �I�[ ��_= wwo��,bD� ���|GG�� �����4� �e� v�ʷ� ��&�� 2��Z uz������� �w�TW&q~q �5�׷&�o?� ;0��  �{2� �y� ����W&���� ?�3� A���e�/> �{\�3&T��� �77߸ ��ֽ� ���� �{���&��8 ��l1��S�)� ���d *{J� F's �~��� 6:0�� ��,��s�- Q�v� ���� �,�T� �ZBLx6����6 ��6���N�Par ��s>�tE��j�6dsq��F  �������ЁDhel�����ti-S�� �Ob��Dbcf�O�����+t OFT��P<A� _�V�ZI��D��V�\�qWS��= dt�le�Ean�(bz=d��titv�Zҥz�Ez XWO �H6�6���5 H^�6H691�E4܀�TofkstF� Y6�82�4�`�f80M4�E91�g�`30oBkmon_�E��e�ݱ�� qlm��0� J�fh��B�_ / ZDTfL0�fw(P7�EcklKV0� �6|��D85��ّ�m\b����xo�kn�ktq��g2.g����yLbkLVtms��IF�bk��x����Id I/f���GR� �han�L��Vy��%��%ecre�����io��w ac�- A�qn�h���cuACl�_�^ir��)�g�2�	.�@�& G��R630���p v�p`�&H�f��un���R57v�OJavpG�`Y��owc��-ASF��O��7���SM�����v
af��raf�La�vl�\F c�w a���?VXpoV �{30��NT "L�FFM��=����yh	�a�G-�w�� �m�2.�,�t��̹�g6ԯ��sd_�#MC'V����D����fslm�isc�.  Hg5522��21&d�c.pR78�����0�708�J614Vip ATUu�@�OL�545ҴI�NTL�6�t8 (�VCA���sseCRI���ȑ��UI���rt\�rL�28g��NRmE��.f,�63!���,�SCH�d Ek�DOCV���p���C,�<�L�0Q�isp��EIO��xE,У54����9��2w\sl,�SETĸ��lр�lt2�J�7�ՌMAS�K��̀PRX�Y҇��7���OC-O��J6l�3�l�� (SVl�A�H�pL�@Օ��539R�sv���#1��L�CH���OPLG.f�outl�0��D��HCR
svgb��S@�h��CSaԌ!�{�50��D�l�5�!�lQ��DSW��S0����̀��OP����M7��PR���L�Ҟ��(Sgd���P�CM���R0 \Es��5P՝���0��X��n�q� AJ�1��tN�q�2��PRSa����69�� (AuFRD�Խ���RMCN���93�A�ɐCSNBuA�F9� HLB���� M��4���h�2vA�95z�HTCa�ވ�TMIL6�j9y5,��857.,�PA1�ito��T�PTXҴ JK�T�EL��piL�� 4XpL�80�I)��.и!��P;�J95��s� "N���H�UE�C��7\cs�F�R��<Q��C��57\{VCOa�,����IP1jH��SU�I�	CSX1�A�WEBa��HT�Ta�8�R62��md`��GP%�IG %�tutKIPGS�j�| RC1_meN�H76��7P��ws_+�?x�R51�\iw�N��ԦH�53!��wL�8!�h�R66��H����Ԡ���@;J5�6��1���N0��9�j2��L���R5`%�AJ|�5q�r�`,�8 5���{165!��@�"5l��H84!�29��Ⱦ0��PJ���n �B[�J77!Ԩ�RA6�5h3n���y36P��3R6��-`;о Ը�@��exeKJs87��#J90!��stu+�~@!䬵��k90�kop �B����@!�p�@|B�A�g*�n@!��Q��06!�@[�F�FaP��6��́,�TS� �NC[�CAB$i4Ͱl1I��R7��@�q�y�CMS1�r�og+QM�� �� T�Y$x�CTOa�n�v\+��1�(�,�6��con�~0��1]5��JNN�%e:�8�P��9ORS%xк��8A�815[�FCBaUnZQ�P!��p�{��CMOB��"�G��OL��x�OP]I�$\lr[�SŠ��T	D7�U��CPRMQR9RL���S�V��~`���K�ETS �$1��0���3�Ԯ��FVR1�LZQVc3D$ ���BVa��SAPL1�CLN�[�PV��	rCCG�aԙ��CL�3C{CRA�n "W!�B�H�CSKQn�\0�p��)�0CTPn�ЌQe��p!$bCt�aT0U�pGCTC�yЋRC1��1 (�s��trl�,�r��
TX��T�Caerrm�r�M�C"�s��#CTE���nrr�REa�XqPj�^��rmc�$^�a"�P�QF!$�\��$p "�rG1䖈tTG$c8��QHܑ$SCTI�! �s��CTLqdAC�K�Rp)��rLa�R82��M��YPk�.���OF��.���e�{��CN���^�1�"M �^�a�С�Q`US��T!$��M�QW�$m��VGF�$R MHv��P2�� H5� �ΐq��ΐ�$(MH[�VP�uoY����$�)��D��hg��V{PF��"MHG̑�`e!�+�V/vpcm��N��ՙ�N��$�VcPRqd)��CV�x�V� "�X�,�1�(${TIa�t\mh��K��etpK�A%bY�VP%ɠ�!PN����GeneB�ri�p����8��e�xtt���Y�m �"�(��HB�� �)��x������x�Ȣ�res.�yA�ɠn�����*���p�@M�_�NĀ6L���Ș�yAvL�Xr�Ȉ2��s"R;�Ƚ\ra���	P�� h86��Gau+ʸ�Ͽ�SeL��m�9�69�P�Ȩr`�Ȩ2�ɹ1��n2��h� �0L�XR}�RIB{�e� L�x���c�Ș���N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1��/�k�@���A���ruk�ʘ L�so1p��H�}�ts{���ĺ��s��9��j965��Sc��h��O5 J9�{�
�P�L�J	een��ts I[
x�com��9Fh�L�4 J�v�fo��DIF+��6�Q����rati�|��p��1�0�
R8l߾�M�����P��!8� �j�mK�X� HZ����N��oڠ��3�q��vi̋��80�~�l aSl�yQ��tpk�xb�j�.�@�R�d�������,/n(�8�8 �0���
:�O8�<�LQ}�CO���PT��O (��.�Xp|��~H���?�v f�wv��8�22�p�m���722��j�7�^�@ƙ���cf��=Yvr���vcu���O�O�O�O_�#_5_7�3Y_��wv�4{_�_w�ʈ�u�st_�_�cus �_�Z��oo,o>oPo8�io��nge��(p�Ly747�jWel�ʨHM47ZKEq� {���[m�MFH�?�(wsK�8J��n���o��fhl�;��wmf���? �:�}(4	<g J�{��II)̏މw��X�774kﭏ/7�ntˏ݊e+���se�/�aw��8�ɐR��EX \�!+: �p,��~�00��nh�,:�Mo+�xO��1 "YK�O��\a��#0 ��.8���{h�L?�j+N�mon�:��t�/&�st�?-�w�:� ��)�;��(=h�;
�d Pۻ�{:  ��� �J0���re����S�TD�!treLANG���81�\tqd�������rch.��ռ���htwv�WxWָ� R79���"Lo�51 (��I�W�h�Ո�4�aSww� �vy ��623c�h a?�cti�֘!�X��iؠ�t ��n@,�։����j��"AJP@�3p�Svr{�H�6��!��o- SeT� E3ּ) G�J934��L=oW�4 (S����p��� <���91 ��8!4�j9�所+��ٲy�
��	�btN�ite{�R ��I@� ������P�������p	 ����Z�vol���X ��9�<�I�p���l�d*���F�864{��?��K�	�k�����֘1�wmsk���M�q�Xa�e ����p��0�RBT�1ks.OPTN�qf�Uz$ RTCamT ��y��U��y��U��UlU6L�T�1 Tx����SFq�U�e�6T��USP W�b DT�qT2h�T�!/&+��TX�U\j6&�Up U�UsfdO&��&ȁT���66�2DPN�b0i��%�Q�%62V��$����%�� �#(�(6T=o6e St�%���#5y�$�)5(T�o�%tT0�%5�W6Tp���%�#�#orc���#I���#���%ccat�6ؑ?�4\W6�965"p6}"�#\j536���4�"�?GkruO O,Im?Np�C �?t�0<O�;�e �%���?
;{gcJ7 "AV�?�;avsf�O__�&_8WtpD_V_0GT��F|_:UcK6�_�_r��O�3e\s�O2^y\`O:�migxGvgW'! m�%��!�%T�$E A{6�po6�f�#37N�)5R5_�2E���$0���$Ada�Vd���V�?;Tz78�_�e7DDTF9���#8�`�%��4y�?ted Z@�A}�@�}�04N�}�}���}�dc& }���	�u 6�v��v1�u1\b�u$2}���}� R83�u�"}�<�"}�valg���Nrh�&�8�J�Y��o�ue��� j70��v=1��MIG�uerfa��{q���E�qN�ء��EYE�ce A���񁏯p V�e�A!���2Յ�Q�%��u1�e�i�@��H� e����J0� '��bx��T��E In��B�  W�|��53q7g����(MI��t�Ԇr��ݟ�a!m���nеv!g�U -�v J߆8⹖F���P�y�ac���2���Rɏ jo��2��� djd�8r}� Gog\k�0��g��wmf�Fro�/� Eq'�4"}�3� J8��oni�[��ᅩ}Ĵ�� !o� ��ʛ��m@�RΉe��{n�Д�V�o������  �����⣆"PO�S\����ͯ me�nϖ�⑥OMo�4q3��� �(Coc� An[�t���"e��a\�vp��.��c7flx$�le��8ٰhr�tr�NT� �CF+�x E/�t0	qi�M�ӓxc��p��f�lx����Z�cxb��
0 h��h8��3mo��=� H����)� (�vSER,����g�0߆0\r��vX�= ��I � -� �ti��H��V]C�828�5���L"�RC��n G�/���w�P�y�\v�vm "o�lϚ�x`а�=e�ߠ-�R-�3?������vM [�A�X/2�)�S�rxel�v#�0��h8߷^=� RAX�A�����9�H�E/R�צ����h߶"RXdk��F�˦85���2L/�xB885t_�q�Ro�0iA��5\rO�9�K��v�����8���.�n� "�v��88��8 s�i ?�9 ��/p�$�y O�MS"�x��&�9R H74&�`�745�	p��8p��ycr0C�c�)hP0� j�-�a%?�o��6D950R7tr�l��ctlO�AcPC���j�ui"��L���  ����^%ࣆ!�A��qH��z�&-^7���w ��616C��q�794h���� qM�ƔI��99����(��$FE�AT_ADD ?_	���Q%P?  	�H._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n ���������TDEMO �fY    WM_���� ����//%/R/ I/[/�//�/�/�/�/ �/�/�/?!?N?E?W? �?{?�?�?�?�?�?�? �?OOJOAOSO�OwO �O�O�O�O�O�O�O_ _F_=_O_|_s_�_�_ �_�_�_�_�_ooBo 9oKoxooo�o�o�o�o �o�o�o>5G tk}����� ���:�1�C�p�g� y�������܏ӏ��� 	�6�-�?�l�c�u��� ����؟ϟ����2� )�;�h�_�q������� ԯ˯ݯ���.�%�7� d�[�m�������пǿ ٿ���*�!�3�`�W� iϖύϟ��������� ��&��/�\�S�eߒ� �ߛ��߿�������"� �+�X�O�a���� �����������'� T�K�]����������� ������#PG Y�}����� �LCU� y������/ 	//H/?/Q/~/u/�/ �/�/�/�/�/??? D?;?M?z?q?�?�?�? �?�?�?
OOO@O7O IOvOmOO�O�O�O�O �O_�O_<_3_E_r_ i_{_�_�_�_�_�_o �_o8o/oAonoeowo �o�o�o�o�o�o�o 4+=jas�� ������0�'� 9�f�]�o��������� ɏ�����,�#�5�b� Y�k���������ş� ���(��1�^�U�g� �������������� $��-�Z�Q�c����� ��������� �� )�V�M�_όσϕϯ� ����������%�R� I�[߈�ߑ߫ߵ��� ������!�N�E�W� ��{���������� ���J�A�S���w� ������������ F=O|s�� ����B 9Kxo���� ��/�/>/5/G/ t/k/}/�/�/�/�/�/ ?�/?:?1?C?p?g? y?�?�?�?�?�? O�? 	O6O-O?OlOcOuO�O �O�O�O�O�O�O_2_ )_;_h___q_�_�_�_ �_�_�_�_o.o%o7o do[omo�o�o�o�o�o �o�o�o*!3`W i������� �&��/�\�S�e�� ������������"� �+�X�O�a�{����� �����ߟ���'� T�K�]�w��������� �ۯ���#�P�G� Y�s�}��������׿ ����L�C�U�o� yϦϝϯ�������� 	��H�?�Q�k�uߢ� �߫���������� D�;�M�g�q���� ������
���@�7� I�c�m����������� ����<3E_ i������ �8/A[e� �������/ 4/+/=/W/a/�/�/�/ �/�/�/�/�/?0?'? 9?S?]?�?�?�?�?�? �?�?�?�?,O#O5OOO YO�O}O�O�O�O�O�O �O�O(__1_K_U_�_ y_�_�_�_�_�_�_�_ $oo-oGoQo~ouo�o �o�o�o�o�o�o  )CMzq��� ������%�?� I�v�m����������ُ���;�  2�Q�c�u����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�9� K�]�o����������� ������#5GY k}������ �1CUgy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o�o�o�o +=Oas��� ������'�9� K�]�o���������ɏ ۏ����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������ +=Oas��� ����'9  :>U gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����� ����/�A�S�e� w���������я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{�����@��/=C6Yk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/AS ew������ �+=Oas �������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�� ������!�3� E�W�i�{�������Ï�Տ�����/�A���$FEAT_DEMOIN  E���q��>�Y�I�NDEXf�u���Y�ILECOMP g������t�T���SETUP2 h������  N� ܑ��_AP2B�CK 1i�� � �)B���%�C�>���1�n�E� ���)���M�˯���� ���<�N�ݯr���� ��7�̿[��ϑ�&� ��J�ٿWπ�Ϥ�3� ����i��ύ�"�4��� X���|ߎ�߲�A��� e�����0��T�f� �ߊ�����O���s� ����>���b���o� ��'���K������� ��:L��p���� 5�Y�}�$� H�l~�1� �g�� /2/�V/ �z/	/�/�/?/�/c/ �/
?�/.?�/R?d?�/ �??�?�?M?�?q?O��?O<O���P�� 2�*.VRCO�O�0*�O�O�30�O�O�5w@PC�O_>�0FR6:�O=^�Oa_�KT���_�_�&U�_�\h�R_�_�6G*.FzOo�1	(S�oEl�_io�[STM �b�o�^+P�o�m��0iPend�ant Pane	l�o�[H�o �gp�oYor�ZGIF|���e�Oa��ZJPG �*��e����z��JJS�����0�@���X�%
JavaScriptُ�CSʏ1��f�ۏ� %Casca�ding Sty�le Sheet�s]��0
ARGN?AME.DT���<�`\��^���Д����АDISP* ן���`$�d��V�e���CLLB.Z�I��=�/`:\��\������Coll�abo鯕�	PA�NEL1[�C�%@�`,�l��o�o�2a��ǿV���r����$�3 �K�V�9���ϝ�$�4i���V���zό�!����TPEINS.gXML(�@�:\<�����Custom� Toolbar�}��PASSWO�RD���>FRS�:\��� %P�assword ?Config��? J���C��"O��3��� ��i����"�4���X� ��|�����A���e� ����0��Tf�� ���O�s ��>�b�[� '�K���/� :/L/�p/��/#/5/ �/Y/�/}/�/$?�/H? �/l?~??�?1?�?�? g?�?�? O�?�?VO�? zO	OsO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_;_M_�_q_o�_ �_<o�_`o�_�o�o%o �oIo�o�oo�o8 �o�on�o�!�� W�{�"��F�� j�|����/�ďS�e� ��������T��x� �����=�ҟa���� ��,���P�ߟ񟆯� ��9����o����(� :�ɯ^�����#��� G�ܿk�}�ϡ�6�ſ /�l�����ϴ���U� ��y�� ߯�D���h� ��	ߞ�-���Q߻�������,��$FIL�E_DGBCK �1i������ ( ��)
SUMMA�RY.DG,����MD:`�����Diag Sum�mary���
C?ONSLOG��y������$���Con�sole log�%���	TPACC�N��%g������TP Accou�ntinF���F�R6:IPKDM�P.ZIP����
���)����Exception-�����MEMCHECKК����8�Me�mory Dat�a��LN�)�RIPE����0�%� Packet LE����$Sn�ST�AT*#� �%LStat�us�i	FTP��/�/�:�m�ment TBD�=/� >)E?THERNE�/�o�/�/��Eth�ernU<�fig�uraL��'!DCSVRF1//)/B?��0 veri?fy allE?��M(5DIF�F:? ?2?�?F\8d�iff�?}7o0CHGD1�?�?�?LO� �?sO~3&��
I2BO)O;O�O qbO�O�OGD3�O8�O�OT_ �O{_�
VUPDATE�S.�P�_��FR�S:\�_�]��U�pdates L�ist�_��PSRBWLD.CMo����Ro�_9�PS�_ROBOWEL<^/�/:GIG��o�>_�o�GigE� ��nostic�W�N�>�)>�aHADOW�o�o��ob�Shad�ow Changye��8+"rNOTI?=O���Notifi�c�"��O�A�PMIO�o���h��f/��o�^U�*�UI3�E�W��{�UI������B��� f��_�������O�� �������>�P�ߟt� �����9�ί]�򯁯 �(���L�ۯp���� ��5�ʿܿk� Ϗ�$� 6�ſZ��~��wϴ� C���g���ߝ�2��� V�h��ό�߰���Q� ��u�
���@���d� �߈��)��M����� �����<�N���r�� ��%�����[���� &��J��n�� 3��i��"� X�|��A �e�/�0/�T/ f/��//�/=/�/�/��$�$FILE_��PPR�P���� �����(MDONLY �1i5�  
 �z/Q?�/u?�/�? �?t/�?^?�?O�?)O �?MO_O�?�OO�O�O HO�OlO_�O_7_�O [_�O_�_ _�_D_�_ �_z_o�_3oEo�_io �_�oo�o�oRo�ovo �oA�oew �*��`����&�O��*VISB�CK,81;3*.�VDV����FR�:\o�ION\DOATA\��/���Vision VD filȅ ��&�<�J�4�n��� ���3�ȟW������ "���F�՟�|���� ��m�֯e������0� ��T��x������=� ҿa�s�ϗ�,�>��� b���ϗϼ�K��� o��ߥ�:���^�����ϔ��*MR2_G�RP 1j;�C4  B�}Ї	 71������E��� E�  F@ F�5U�������L���M���Jk�L�zp�JP��F�g�f�?�  �S����9�Y9�}�9��8�j
�6��6��;��A�  l���BH��B���B���$��������������@UUU#�����Y�D�}�h� ���������������
C��_CFG {k;T M����]�NO �:
F0� �� \�RM_CHK�TYP  0��}�000��OM�_MIN	x����50X� S�SBdl5:0��bx�Y����%TP_DEF_�OW0x�9�I�RCOM��$�GENOVRD_�DO*62�TH�R* d%d�_�ENB� �R�AVC��mK�� ��՚�/3�/�q�/�/�� �M!kOUW s��}���ؾ��8��g�;?�/7?Y?[?  C��0����(7�?6�<B�?B����2p��*9�N SMTT#�t[)��X�4�$HoOSTCd1ux����?�� M5Cx��;zOx�  27.0�@=1�O  e�O�O 	__-_;Z�O^_p_�_�_�LN_HS	ano?nymous�_�_�_oo1o yO��FhFk�O�_�o�O�o�o �o�oJ_'9K] �o�_����� 4o�XojoG�~�o^� ������ŏ���� �1�T���y����� ������,�>�@�-� t�Q�c�u��������� ϯ���(�^��M� _�q�����ܟ� �ݿ ��H�%�7�I�[Ϣ� ϑϣϵ����l�2� �!�3�E�Wߞ���¿ Կ����
������� /�v�S�e�w���� ���������+�r� �ߖ�s�����߻��� �������'9K] ��������� 4�F�X�j�l>��} ������/ /1/T��y/�/�/�/�/.D\AENT {1v
; P!J/.?  ��/3? "?W??{?>?�?b?�? �?�?�?�?O�?AOO eO(O�OLO^O�O�O�O �O_�O+_�O _a_$_ �_H_�_l_�_�_�_o �_'o�_Koooo2o{o Vo�o�o�o�o�o�o 5�oY.�R��v��zQUIC�C0���3��t1 4��"����t2��`��r�ӏ!ROUT�ERԏ��#�!�PCJOG$����!192.16?8.0.10��s?CAMPRTt�P��!d�1m�����R�T폟�����$NA�ME !�*!�ROBO���S_�CFG 1u�)� �Au�to-start{edFTP&��=?/֯s��� �0�B��f�x����� ����S������,� ��������ϼ�ޯ�� �������ʿ'�9�K� ]�oߒ�ߥ߷�����p����SM% y�{�U�ό����� �����
��.�@�c���v������������z�%�7�I�K�8� \n���k��� ��3�FXj |����a��7/M*/</N/ `/r/9�/�/�/�/� �/�/?&?8?J?\?� m?���?�//�?�? O"O4O�/XOjO|O�O �O�?EO�O�O�O__ 0_w?�?�?�?�O�_�? �_�_�_�_o�O,o>o Poboto�_o�o�o�o �o�oK_]_o_L�o �_�o�����o�  ��$�6�Y�Y�~��������ƏZ�_ER�R w3�я�P�DUSIZ  jg�^�p���>�?WRD ?r�Cq��  guestb�Q�c�u��������`�SCDMNGRP 2xr�w���H��g�\�b�K� 	�P01.00 8~`�   � ��   B � ��� ����H���L���L��L�����O�8�����l�����a�4�  �Ȥ� �V8���\���)�5`�;��������d�.�@�R�ɛ_�GROUېy������	ӑ���Q?UPD  ?u��Y��İTYg�����TTP_AU�TH 1z�� �<!iPend�an��-�l����!KAREL:q*-�6�H�KC]��m��U�VISI?ON SET������!�����R�0� �H�Bߏ�f�x��ߜ������CTRL �{����g�
&�FFF9E3���AtFRS:DE�FAULT;��FANUC We�b Server ;�)����9�K��ܭ�����������߄WR�_CONFIG ;|ߛ ;���IDL_CPU_kPCZ�g�B�I��y� BH_�MIN�j�)�}�GNR_I�O��g���a�NPT_SIM_D_������STAL_oSCRN�� ����TPMODNTOqL������RTY��0y���� �ENO����Ѳ]�OLNK 1}��M��������eMAS�TE��ɾeSLAVE ~��c�O_CFGٱB�UO�O@CYC�LEn>T�_AS�G 1ߗ+�
 ����//+/ =/O/a/s/�/�/�/�/\��NUM��=
@IPCH�^RTRY_CNZ�����@������b�� @kI�+�E�z?E�a�P_ME�MBERS 2��ߙ� $���2����ݰ7�?�9a�SD�T_ISOLC � ����$J2/3_DSM+�3JOBPROCNn��JOG��1�+��d8�#?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSR�EQO��KANJI�_���a[�MO�N ����b�y N_goyo�o�o�o�Y�`3�<� ��e�_ִ���_L���"?`EYLOGGINL�E�������$�LANGUAGE� ��<T� ,{q�LGa2�	�b�마g�xP��  U��g�'���b���>�MC�:\RSCH\0�0\<�XpN_DISP �+G�H�8�O�O߃LOCp��Dz���AsOGBOOK �������󑧱����X �����Ϗ����0a�*��	p������!�m��!���=p_BUFF 1�p��2F幟����՟D� Coll�aborativ ǖ���F�=�O�a�s� ������֯ͯ߯����B�9�K���DCS� �z� =���'�f��?ɿۿ���|H@{�IO 1��G ~?9Ø��9� I�[�mρϑϣϵ��� �������!�3�E�Y� i�{ߍߡ߱�������Z�E��TMNd�_ B�T�f�x������ ��������,�>�P��b�t�������L��S�EVD0��TYPN1�$6����QRS"0&��<2F�L 1�"�J0� �������FGTP:pOF�NGNAM1D�mrn�tUPS�GI"5��aO5�_LOA�DN@G %�%�DF_MOTN��y�� MAXUALRM�'���(��'_PR"4F0d��1��B_PNP� V� 2�C	M�DR0771ߕz�BL"8063%�@ �_#?�ߒ|/�C��z�6��/􈃟/Po@P 2���+ �ɖ	~T 	t  ��/ �%W?B?{?�k?�? g?�?�?�?O�?*OO NO`OCO�OoO�O�O�O �O�O_�O&_8__\_ G_�_�_u_�_�_�_�_ �_o�_4ooXojoMo �oyo�o�o�o�o�o �o0B%fQ�u �������� >�)�b�M�����{��� �����Տ��:�%��^�p�S�������D�_LDXDISA�pB�MEMO_{APjE ?C
 �,�(�:��L�^�p������IS�C 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%A �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A?���?IܿI���pW�Q_D��^��PL_NAME �!3%,�!�Default �Personal�ity (fro�m FD) �R�R2� 1�L?6(L?�,0	l d���� ����//(/:/ L/^/p/�/�/�/�/�/�/�/ZX2u?0?B? T?f?x?�?�?�?�?\R<?�?�?O O2ODO�VOhOzO�O�O�OZZK`\R�?�N
�O_\TP�O:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHo_)_~o�o �o�o�o�o�o�o  2DVhz�[omo ����
��.�@� R�d�v���������Џ�� Ef  Fb� F7���   ��!��d��@�R�6�t��� ���l���ʝ����� ݘ���� "�@�F�d���� "�|��ݐA�  ϩ�U[�$n�B��E ��� � @D�  &�?�� �?�@��A@�;f��FH�� ;�	l,�	 '|��j�s�d�/>��� ��� �K(��Kd$2�K ��J7w��KYJ˷�ϜJ�	�ܿ�� @�I���_f�@w�z��f��γ�N��� ���	Xl�����_��S�ĽÔ�}�X�����5�?��  ����A�?oi#�;���A��� ���l� �Ϫ�-���PܛG�G�Ѳ��@�n�@a   ?�  ��ܟ�*�͵	'� �� H�I� ��  �Рn�:��Èl�È=��9̈́�в@�ߚ� �����/������̷NP�  '�,���-�@
�@W���?=�@A����B�  CTj�a�Be�Ci��@�#�Bи�L K ,ee��/^^ȹBР��P����̠�����ADz՟�n�3��C�i��@�R�R�Yщ��  =�@� ��Ż�=��?�ff������n� ɠ#ѱ@y9G
(���I�(�@uP~����t�t����>����;�Cd;���.<߈<��g�<F+<AL�������,�d�|,�̠?fff?���?&&��@���@x��@�N��@���@T� H�ِ�!-�ȹ�| ��
`������ �//</'/`/r/]/�/��eF���/�/ �/�/m?��/J?�(�E��G�#�� FY�T?�?P?�?�? �?�?�?O�?/OO?O eOk���O�IQOG�? �O1?�OmO_0_B_T_"������A_�_@	_�_�_�_ o��A��aAn0 bФ/o C�_pUo�_�Op��؃o��o�o�o���W������oC�E�  q�H�d��؜a@q���e�F�BµWB�]�NB2�(A���@�u\?��D�������b��0�|�uR�Ｃ�
x~������Bu*�C��$�)`��$ ���GC�#���rA�U����1��eG�D�I�m�H�� I:��I�6[F����C�I��J��:\IT�H
~QF�y���p�*J�/ �I8Y�I��KFjʻCe�o�� s�����Џ���ߏ� *��N�9�r�]����� �������۟���8� #�\�G�����}����� گů���"���X� C�|�g�����Ŀ��� ����	�B�-�f�Q� ��uχ��ϫ������ ��,��P�b�M߆�q� �ߕ��߹�������(� �L�7�p�[����������s(���33:����$���3���d�,�4���@�R��񴲚�l�~�wa���ex����wa4 �{�� ����(L:ue%P�P~�A�O�������	����G2W} h������/����O�O7/m/[(d =�s/U/�/�/�/�/�/ ?�/1??U?C?y?�=  2 Ef9g�Fb��77�9fBX)aa)`C9A`�&`w`@-o�?9de�O-O?OQOpn�?�?�O�O��O�O9c?�0�A7hJt4w`w`!w`xn
 �O9_K_ ]_o_�_�_�_�_�_�_��_�_o#ozzQ ���h��G���$�MR_CABLE� 2�h ��a�T� @@��0�Ae��a�a�a���`��0�`C�`�aO�8�tB�n���yA�aE�M�GE�#�o�f�#���0��0�DO���By`��޾�*��bE�E��c,��o�g8 [ ���C�07�dw4
v��d����b��E��Z&�l�`y`
qCܛp�bHE�
v���5D�_)D�SҮz�lҠ`��0��q�p�b0�
u��ԋ��b?]�E;h��u/o�c -��4tH�\�?�9�K� ]�o�ԏϏ��
�ɏۏ�@���?��eo �a���������b����� �����`�	 ����@������% �*�}0�6 ��ݐ�����`���	����@������*,� ,�-�\c�OM �ii���3� ��L~@%% 23�45678901�i�{� f��������ԋ��1����
���`�not �sent3������;�TEST�FECSALGR  egfJ�1iqiqZš
:�� �D�CbS�Q�c�u��� 9�UD1:\ma�intenanc?es.xml��ֿ�q� =���DEFAULT�-��4\bGRP 2�M�  =��a��{p  �%�Force�s�or checkS  ���b�z��p����h5-[ �ϻ�������ϖ�D�%!1s�t cleani�ng of co�nt. v�ilation��}�R��+��[�ߔߦ߸�z��mech�'cal`����p�!�0��h5k�@��R�d�v�����(�rolle_Ƶ����/���(�:�����Basic q�uarterly�������,������0����M��M��:@"GpP�a�b`�4�������#AC���M"��{�Pbt���S�uppq�greaCse���?@/&/8/J/\/��C+ �ge��. batBn�y`/��/h5	/ �/�/�/? ?_�ѷen'�v��/�/��/��?�?�?�?�?ѣG=?O�qp"CrB1O��0�/`OrO�O��O�O�t$��Lf�B�C-m��A�O:�OO@$_6_H_Z_l_�t*�cabl�Om���B�S<m��Q�_:�
_ �_�_oo0oo)(Ӂ/�_�_���_�o�o�o��o�o�O@ha�u1�l�2r xm�<qC:��op������ReplaW�fUȼ2�:�._4�F�X�j�|�m�$%���o�������#� ��
��.�@���d��� ŏ׏����П���� U�*�y�����r����� ����	�q��?�߯c� 8�J�\�n���ϯ���� �ڿ)����"�4�F� ��jϹ�˿������� �����[�0�ϑ�f� �ϊߜ߮�����!��� E�W�,�{�P�b�t�� ���߼�����A�� (�:�L�^�������� ������� $s� H������q��� ��9]o�V hz���U�# �G/./@/R/d/� �/�/��//�/�/? ?*?y/N?�/�/�?�/ �?�?�?�?�???Oc? u?JO�?nO�O�O�O�O+J�r	 H�O�O_ _6M2_@OBE:_p_>_ P_�_�_�_�_�_ o�_ �_oHoo(oZo�o^o po�o�o�o�o�o �o� :z �bA?�w  @�q _ ���Fw�� ��H* �**  @q>v�p2T�f�x�:�p������ҏ��eO ^C7�Տ#�5�G�	�k� }���ُ���c���� �W��C�U�g���ß )�����ӯ���	�� -�w�����9��������m�Ͽ��=�O�E�	A�$MR_HI_ST 2�>uN��� 
 \�$Force� sensor �check  1�23456789�0q�3����ß��N}SB�� -319.8 �hours RU�N 9.�Y�!1�st clean�ing of c�ont. ven�tilation�0ÄϖϨ�-�Y�޹�mech��ca�li�%Ό4��o��DN�t��95���1����rol�leh�+�=�O���Y�Basic �quarterlyߒߤ߶�
O4�F� �(�����b�t� ����������M�_� ���:�����p���:��SKCFMAP � >uQ���r5�������ONREL  .��3���EXC'FEN��:
���QFNCXJJO�GOVLIM8d�Ná ��KEY8z��_PAN7�����������SFSPDTYqPxC��SIG�|:��T1MOT��G��_CE_G�RP 1�>u\�D����� /Ⱥ��/�/U/ /y/0/n/�/f/�/�/ �/	?�/???�/c?? \?�?P?�?�?�?�?�?�O)OOMO,���QZ_EDIT5 )�TCOM_CFG 1���[�O�O��O 
�ASI 	�y3�
__+[!_O_��>O�_~bHT_ARC_U�քT_MN_oMODE5�	UAP_CPL�_�gNOCHECK� ?�� �� o.o@oRodovo �o�o�o�o�o�o�o�*!NO_WA�IT_L4~GiN�T�A���EUwTo_ERRs2���3��ƱJ������>_)��|MO�s���}x:EB�  B�4  �r�x���8�?������ �~�rPARAM��r������r_�:H5�5�G� =  r�b�t�s�X��� ���������֟�0��:G�b�t������SUM_RSPA�CE�����Aѯۤ�$ODRDSP�S�7cOFFSET�_CARt@�_�D�IS��PEN_FILE:�7�AF��PTION_I�O��q�M_PR�G %��%$*�����M�WORK ��yf ���춍���� �� �������	� ������It���RG_DSBOL  ��C�{�u��RIENTT�O7 ��Cn�A� �UT_SIM�_Dy���V~�LCT ��}�{B �٭��_PEX��P=��RAT�W �dc��UP S���`���e߰w�]ߛߩ��$�2�r�L6(L�?���	l d ������&�8�J�\� n��������������"�4�F�X���2 �߈�������������*�<w�Tf x�������8J` �D T��Tz�Pg� �����/"/4/ F/X/j/|/�/�/�/� ��/�/??0?B?T? f?x?�?�?�?�?�?�? �?�/�/,O>OPObOtO �O�O�O�O�O�O�O_�_(_:_��O*��y_�]2ӆ��_�^�_ �_�W^]^]��/ooSog��Hgrohozo�o �o�o�o�oF`�#|>G`A�  9y�����OK�1�k_�����<��EA�~nq @D�  �qh����nq?��C��s��q1� ;�	l>��	 |�Q�sy�r�q>��u�
��qF`H<zH�~�H3k7G�L�zHpG�99l7�k_B�T��F`C4��k�H���Rt��-�:����k������s���  �ሏ����Ee�BVT���dZ>�����ڏ ���q-�Fk�yԵ{FbU���n�@6�  ����z�Fo��;�	'�� � ��I�� �  �<:p܋=���ڟ���@���B��,���B���g�:�N����  '|���g�V�B��p�BӀ�C׏����@  #��Bu�&�e�e�^^މB :p2���>�m�6p�Z���Dz?o}�܏���� ��׿������Ǒ���� f�  � ��M���*�?�ff0�_8�J�ܿ 3p���ñ8�Чϵʖq.���(����P���'���s�tL�>��/�;��Cd;��.<�߈<�g�<F+<L ��^oi��rd@��r6p?ff�f?�?&��;�@���@x��@��N�@���@T싶�Z���ћt މ�u�߈w	�x��ti� >�)�b�M��q��� ����������:�%��^�������W����E��  G�aF�� Fk������� ��1U@yd� �����q��	� �{�A��h������a��ird��A {/w/J/5/n/v�A��A���":t�/ �C^/�/Z/ ލ?Ƀ��/�/1??��ĥW����g��pEC� ~1�?04�0�
1�1@IӀ��B�µWB]�NB�2�(A��@�u\?����������b�0�|��uR����
��>�ؽ���Bu*C��$��)`�? ����GC#������rAU����1�eG����I�mH�� �I:�I�6[�F���C4OI���J�:\I�T�H
~QF�y�Ol@�*�J�/ I8Y��I��KFjʻC��-?�O�O__>_ )_b_M_�_�_�_�_�_ �_�_o�_(oo%o^o Io�omo�o�o�o�o�o  �o$H3lW �{������ �2��V�h�S���w� ����ԏ�������.� �R�=�v�a������� П����ߟ��<�'� `�K�]���������ޯ ɯ��&�8�#�\��3=(J���3:a��s����J�3��c48������������1����ڿ��1����e���14 �{2�2�r�`ϖ�P�ϺϨ��%PR�P���!�h�!�K�6�<o��)����u�|� �ߠ����������3� �W�B�{�f�4���������d�A����!� �1�3�E�{�i��������������  2 wEf�7Fb��7��6B�!�!� C%9� �� �0@�/`�r������#�x��+=�3?�, V�8v��0��0��0�.
 D�����/ /%/7/I/[/m//�/��:� ��ֻ�G����$PARA�M_MENU ?�2�� � DEF�PULSE�+	�WAITTMOU�T�+RCV? �SHELL_�WRK.$CUR�_STYL� �4<OPTJJ?PT�B_?Y2C/?R_DECSN 0�Ű<�? �?�?�?�?OO?O:O LO^O�O�O�O�O�O�!�SSREL_ID�  .�����EU�SE_PROG �%�*%�O0_�CC�CR0�B���#CW_HOST !�*#!HT�_=ZT��O_��Sh_zQ�S�_<[_�TIME
2�FXU~� GDEBUG�@��+�CGINP_F�LMSKo5iTR\Do5gPGAb` %l��tkCHCo4hTWYPE�,� �O �O�o#0Bkf x������� ��C�>�P�b����� ����ӏΏ����� (�:�c�^�p�����7eWORD ?	�+
 	RSc`^��PNS��C4��JOv1��TE<�P�COL�է��2��gLP 3������OjTRACE�CTL 1�2���! ��c �Қ�q�D/T Q�2�Ǡ���D � ��7:�ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖπ�Ϻ��������� �6�H�Z�l�~ߐߢ� $߶���������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~������� Щ*<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6Fl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�x�N�߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�?�?�?�?�9�$PG�TRACELEN�  �1  �_��0��6�_UP ��K��A@�1�����1_CFG M�E�3�1
@�<D�0<DZO<C��0uO$BDEFSP/D �/L�1�0���0H_CON?FIG �E�3W �0�0d�DM��2 �1�APpD�sA�A�0��0IN~'@TRL �/M�OA8pEQPE�E��G�A<D�A�ILID(C�/M	~bTGRP 1ýI� l�1B�  �����1A��33FC� F�8� E�� @eN	�A�AsA�Y�Y�A~�@� 	 vO8�Fg�_ ´8cokB;`baBo,o>oxo�bo�o�1>о�?�B/�o�o~�o �=%<�� 
C@yd���"������  Dz@�I�@A0�q�  �������ˏ���ڏ ���7�"�4�m�X����|���Ú)ґ
V�7.10beta�1HF @��=��Aq��Q�  �?� �B�ܠP�p �C���&�B�EQA� ��Q�P�Q�� ß[�m����<CA��0�b��@���f�������ҡ�R�ܣ�Rљ����1�i�������t<B!CeQKNOW_M  lE|7FbTSV ĽJ�BoC_�b�t��� ����������1�]aSuM�SŽK ����	NB�0����ĿK���-�bb��A�RP�����0�Ŗ��bQMR
�S��T�iN���d����V]ST�Q1 {1�K
 4MU�iǨj� K�]�o� �ߓߥ߷�������2� �#�h�G�Y��}�� �����
������,��27�I��1�<t�H��P3^�p������,�4��������,�5 (:,�6Wi{�,�7�����,�8�!3,�M�AD�6 F,�O�VLD  K�D�xO.�PARNUM  �MC/%�WSCH� E
9'p!G)�3Y%UPD/���E�/P�_CMPa_��0@�0'7E~�$ER_CHK�%a5H�&�/�+RS���bQ_MO�+?=5�_'?O�_RES_G6��:�I�o�?�? �?�?O�?O7O*O[O NOOrO�O�O�{4]��<�?�Oz5���O_ _|3 #_B_G_|3V  b_�_�_|3� �_�_�_ |3� �_�_o|3Oox>oCo|2V 1�:�|k1!�@c?�=2THR_INRc0�i!}�o5d�fMASmS�o Z�gMN�o��cMON_QUEUE �:�"�j0���O�N� U1N8v�+DpENDFqd?�`yEXEo`u� B�EnpPAsOPTI�OMwm;DpPROG�RAM %$z%�Cp}o(/BrTAS�K_I��~OCFG �$��K��DATA��T�	��j12/ď֏� �����+�=�O�a�����������͟��IN+FO�͘��3t�� !�3�E�W�i�{����� ��ïկ�����/��A�S�e�w������� '��FJ�a K_�N��T��˶EN!Bg ڽw1��2���GN�2�ڻ P�(O�=��]ϸ�@���v� ��u�uɡdƷ_EDIT �T������G�WERFL��x�c)�RGADJ� Ҷ�A�  $�?j00��a�Dqձ�ӆ5�?I��ʨ�<u�)%e`������FӨ�2�R�V�	H;pl�G�b�_�>�pAod�t$��*�/� **:�j0�$�@킆5Y�T���^��q �߈b~�L��\�n�� ������������ ��4�F�t�j�|����� ��������bL BT�x���� :��$,�P b���/��� �/~/(/:/h/^/p/ �/�/�/�/�/�/V? ? ?@?6?H?�?l?~?�? �?�?.O�?�?OO O �ODOVO�OzO�O_�O �O�O�O�Or__._\_ R_d_�_�_�_�_�_�_�f	g�io�pWo�o{d �o�~o�ozo�B�PREF ��Rږp�p
�IOORITY�w[���MPDSP�q��pw�UT6����ODU[CT3���v��OG��_TG���8��ʯrTOENT� 1׶� (!AF_INE�p�,�7�!tcp|7�_�!udN�~��!icmv���ޯrXYK�ض���q)� ,�����p��&�	��R� 9�v�]�o�����П�������*��N�`�*�sK��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b��t����u�w�HANCE �R��:�Bwd��连�2s�9�Ks��PORT_WNUM�s�p����_CARTR�EP{p�Ω�SKS�TA�w d�LGmS)�ݶ��t���pUnothing�������{��TEMP ޾y���'e��_a_seiban�o\��o lߒ�}߶ߡ������� ��"���X�C�|�g� ������������� 	�B�-�f�Q���u��� ����������, <bM�q��� ����(LٟVERSIyp�w�} disa�bledWSAV�E ߾z	2600H768S	?�!ؿ�����/ 	5(�r)og+^/y�e{/�/�/�/�/"�*�,/? �p����_�p 1�Ћ�� ������Wh?z?�W*pURG�E��B�p}vgu,�W�F�0DO�vƲ�vW�%��4(�C�WRUP�_DELAY ��\κ5R_HOT %Nf�q׿GO�5�R_NORMAL�&H�r6O�OZGSEM�IjO�O�O(qQSKKIPF3��W3x= _98_J_\_]�_�_ {_�_�_�_�_�_�_	o /oAoSoowoeo�o�o �o�o�o�o�o+= aOq���� ����'��7�]��K�������)E�$R�A{���K/�zĀ~Á_PARAM�A�3��K @.�s@`�61�2C<�5�y��C�6$�=BÀBTIF�4`�RCVTMOUu��c��ÀDCR�F3��I ��+Q5
=ޅ5�{�3�1.mU_�  �e�W�{B��1�\�k_�-_�yS;�Cd;���.<߈<��g�<F+<L���Ѱ��d�u�L�������ϯ����)�;�M�_���R�DIO_TYPE�  M=U�k�EFPOS1 1�\�'
 x4/���� �+�$/<��$υ�p� ��D���h��ό��'� �����o�
ߓ�.ߤ� Rߌ�������5��� Y���i��*�<�v��� r���������U�@� y����8���\����� ������?��c����/2 1�KԿ�X�T�x��3 1����nY|�S4 1�'�9K�/�'/�S5 1���/�/�/�/:/S6 1�Q/c/u/�/-??Q?>�/S7 1��/�/�
?D?�?�?�?d?S8 1�{?�?�?�?WO�BO{O�?SMASK 1L��O�D�GXNO���F&�^��MOTEZ�Ż��Q_ǁ�%]pA݂��PL_RANG!Q�]�_QOWER ��ŵ�P1VSM_�DRYPRG �%ź%"O�_�UTA�RT �^�ZU?ME_PRO�_�_�4o��_EXEC_?ENB  J�e�GSPD`O`WhՅ�jbTDBro�jRM��o�hINGVERSION Ź�#o�)I_AIoRPURhP �O\(�MMT_�@T�P�#_ÀOBOT__ISOLC�NTV�@A'qhuNAME��l��o�JOB_O�RD_NUM ?��X#qH�768  j1Z�c@�r�rV��s��r�?�r?�r�pÀPC_TIMEu�za�xÀS232>R�1�� L�TEACH PE�NDANw�:GX��!O Mai�ntenance_ Consj2���"��No UseB�׏�������1�C�y�V�NPO��P@�YQ�c�S�CH_L`��%^ �	ő��!OUD1:럒�R�@�VAIL�q@�Ӏ��J�QSPACE1w 2�ż ��@YRs�i�@Ct�YRԀ�'{��8�?� �˯����"���7� 2�c�u�����G���߯ ѿ򿵿�(��u�A C�c�u�����Ͻ�߿ ���ϵ��(��=�_� qσϕ�C߹������� ���$��9�[�m�� �ߣ�Q������߭���  ���	�W�i�{��� M�������5���. S�e�w�����I�� �����*? as��E��� ��/&//;/]o ������/2/�/ ?"?�/7?Y/k/}/�/ �/O?�/�/�?�?�?O�0OOKA��*S�YPpM*�8.3�0261 yB5/�21/2018 �A �WPfG|��H�_TX`� !�$COMME��$USAp� $ENABL{EDԀ$INN`�QpIOR�B�@RY~�E_SIGN_�`��AP�AIT�C�BW�RK�BD<�_TYyP�CRINDXSp�@W�@%VFRI{��_GRPԀ$U�FRAM�rSRTO�OL\VMYHOL��A$LENGT�H_VTEBTIR�ST�T  $�SECLP�XUFI�NV_POS�@$MARGI�A?$WAIT�`�Z�X2�\�VG2�GG1�AI�@�S�Q	g�`�_WR�BNO_US�E_DI�BuQ_R�EQ�BC�C]S$?CUR_TCQP�R�"a^f �GP_S�TATUS�A @ �A3`�BLk�H�$zc1�h�P@����@_�FX ��@E_MLT_C�T�CH_�J�`CO��@OL�E�CGQQ�$W�@w�b#tDEADLOCKu�DELAY_CNaT�a3qGt�a$wf� 2 R1R[1$X<�2[2�{3[3$Zwy�q%Y�y��q%V�@�c�@�b$V4�`�RV�UV3oh>b>�@ � �d�0NarMSKJ�LgWa�Z�C`NRK�PS_R7ATE�0$���S�
`�Q�TAC��PR�D���e�S*��a4�A�0�DG�A 08�P�flp bquS�2ppI�#`
`�P� 
�S\` � �A�R_ENB�Q �$RUNNER_AXI��<`ALPL�Q�RU�T�HICQ$FL�IP7��DTFER�EN��R�IF_C	HSU�IW��%V)�CG1����$PřA�Q��Pݖ_JF�P�R_P�	�RV_�DATA�A � $�ETIM|���$VALU$��	�OP_  � �A  2� �SC*��	� �$IT�P_!�SQ]PNPOU�}�o�TOTL�o�D�SP��JOGLI�b��PE_PKpc�O�f�i��PX]PTA�S�$KEPT_GMIR��¤"`M�b&�APq�aE�@��y�q�g@١c�q�PG�BRK6�x���L�I��  ?�SJ��q�P�ADEz�ܠB�SOCz�MOTN�v�DUMMY16�Ӂ$SV�`DE�_OP��SFSP�D_OVR
��f�@LD����OR��[TP8�LE��F��l����OV��SF��F����bF�d�ƣ&c�)�fQc�LCHDL}Y��RECOV���`��W�PM��gŢ�#RO������_F�?�� @v�S �NVsER�@�`OFS�PC,�CSWDٱc�ձ����B����TRG�|š�`E_FDO���MB_CM}���B��BLQ�¢	�Q�̄Vza�BUP�g��G
��AM���@`�KՊ�e�_M!�d�A�Mf�Q��T$CAԕ���DF���HB�Kd�v���IOU2��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�y3A��ATIO�0��͠��US����WaAB��R+c�`t��`DؾA��_AUX~w�SUBCPUP���S�`����3Եжc8���3�FLA�B�HW_Cwp"�Ns&��]sAa��$UN�ITS�M�F�AT�TRIz�Z�CY{CL�CNECA����FLTR_2_�FI��TARTU�PJp����A��LPx������_SCT*cF_F�F_P���b��FS��+�K�CHA�/Q��*�d�RS�D��Q����Q���_TH�PROr���հGEMPJ���G�T�� �Q�D�I�@y�RAILAiC/�bMX�LOf�xS��ځ���拁��V��PR#�S`appz�C� 	���FUNC���RI�N`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ngDAQ�B�rkLD�र&q�M�K���TI���j���$�@RIA_[SW��AF��Pñ#��%%�p9r1���MOIQ���DF_l~P(�PD"LM-�{FA�PHRDY�DORG�H; _QP|�s%MULSE~P�z���*�� J��J�ײ��FAN_A�LMLVG��!WR=N�%HARDP���UcO�� K2$SHADOW]�kp�a802��� STOf�+�Y_^�w�AU{`R<��eP_SBR�z5����:F�� �3MPINF?�\�4�λ3REGV/1DG��+cVm �C�CFL4(��?�DAiP���Z`�� �����Z�g	 �P(Q$�A$Z�Q V�@�[��
� ��EG0��o���kAAR�����2�axG��AX�E��ROB��RE%D��W�QD�_�Mh�CSYA��AF��FS�G�WRI�P~F&�ST�R����E�˰EH�H)��D�a\2kPB6P��=V��Dv�OTOr�1)���ARYL�`tR�v�3���FI&�~ͣ$LINKb!�\��Q�_3S��8�E��QXYZ2�Z�5�VOFF���R��R�XxPB��`ds�G�cFI�0�3g�������_J��'�ɲ�S&qR0LT2V[6���aTBja�"2�bC���DU�F]7�TUR� X���e�Q�2XP�ЊgFL�E���x@�`�U9Zy8���� 1	)�%K��Mw��F9���8������ORQj��G;W3���#�Ґd ����uz����1�tOV	E�q_�M��ё?C�u EC�uKB�v'0�x-�w H��t���& `��q ڠ�B�ё�u�q�wh�0ECh����ER��K�	�EP����AT�K�6e9e�W���AXs�'��v� /�R ����!��  ��P��`��`�3p�Yp�1�p�� � � �� (�� 8�� H� � X�� h�� x�� �������DEBU��$%3�I��·RA!B���ٱ�sV��� 
d�J、��@� ����������Q���a ���a��3q��Yq+$�`�%"<�cLAB0b8�u�'�GRO���b<��B_s��"T ҳ*`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Q`θuݸ��PNT0~���SERVE �NZ@ $`EAV�!�PO�����nP!�P@�$!Y@�  $>�TREQ�b
=��BG�K��%"2\��� _ � l��5�D6ESRRVb(�I��V0`�;���TOQ:�7�L��@
�R��e G�%ĩQ�� <�50F� �,�`�z�>�RA~� 2 d!�2����S�  M�`�pxU ����OCu�G�  ��C�OUNT6Q��FZ�N_CFGF� 4#��6��TG4�_�=����(���VC ���M �"��`$6��q ��FA E� &��X�@�����H��A����AP���P@HEL�0��� 5b`B_B;AS��RSR�6E�CSH����1�Ǫ��2��3��4��5*��6��7��8��}�ROO����P�PNLEA�cAB)ë ��ACKu�INO�T��(B$UR0� =��_PU��!0��OU+�Pd�8j��� V���TPFWD_KcAR��� ��RE(�� P�P�>QUE�:RO�p�`r0P1I� x�j�P�f��6�QSEM��0��� �A��STYL�SO j�DIX�&������S!_TMCMA�NRQ��PEND�It$KEYSWITCH���k�HE�`BEATM683PE{@LE��>�]��U��F��S~pDO_HOM# �O�@�EF�pPR�aB�A#PY�C� Ox�!���OV_M|b<<0 IOCM�dnFQ&�h�HKYAG D�Q�7��UF2���M���p�cFO;RC�3WAR�"��OM|@  @�S�#o0U)SP�@1*�2&3&4E���*T�O��L���8OUNLOv�D4K$�EDU1  �S�Y�HDDNF� �M�BLOB  �p�SNPX_;AS�� 0@�0|��81$SIZ�1�$VA{���MU/LTIP-��# �A� � A$��� /4`�BS���0�C���&FRIF�BO�S���3� N=F�ODBUP߰`�%@3;9(űp�S��nZ@ x��SI���TEs�r�cSGL�1T�Rp&�Н3B�<�@�0STMTq�3�Pg@VBW�p�4S�HOW�5@�SV���_G�� 3p$�PCJ�PИ���FBZ�PHSP AW��EP@VD�0WCw� ���A00�� PB XG XG XG$ �XG5VI6VI7VI8*VI9VIAVIBVI� XG�YF�0XGFVH��TXbI1oI1|I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1Y1Y2UIU2bI2oI2|I2�I2�I�`�X�I2p�X�IU2�I2�I2�I2�I�2Y2Y�p�hbI3�oI3|I3�I3�I3��I3�I3�I3�I3��I3�I3�I3�I3�Y3Y4�i4bI4�oI4|I4�I4�I4��I4�I4�I4�I4��I4�I4�I4�I4�Y4Y5�i5bI5�oI5|I5�I5�I5��I5�I5�I5�I5��I5�I5�I5�I5�Y5Y6�i6bI6�oI6|I6�I6�I6��I6�I6�I6�I6��I6�I6�I6�I6�Y6Y7�i7bI7�oI7|I7�I7�I7��I7�I7�I7�I7��I7�I7�I7�I7�Y7U�VP� UFD�y"ՠ��
<AT62��t�R��CMD� ��M5�RXv�]��Q_h�R����e����<�YSL|���  � �% \2��+4�'��W�BVALU��b���'���FH�ID_L,���HI��I����LE_��㴦�$�0C�SAC�! �h �VE_B�LCK��1%�D_CPU5ɧ 5ɛ ������C�� ��R �" � PW�j��#0��LA�1�SBћì���RUN_FLG�Ś�����@� ����������H����Х��TBC}2��# � @ B��e �S�8=�NFTDC����V�0��3d�Q�THF������R�L�ESE�RVE9��F��3��2�E��Н�X ;-$��LEN9��F��f�RA��W"G��W_5�b�1��д2&�MO-�T%S60U�Ik�0�ܱF����[��DEk�21LACE�i0�CCS#0�� _�MA� j��z��T#CV����z�T��� ����.Bi�'A�z�'AIJh�#EM5���J���@@i�V�z���2�Q �0&@o�h��JK��VK9��{����f��J0����JJ��;JJ��AAL����(������4��5�ӕ �N1������.�L�D�_�1* �C�F�"% `�GRCOU���1�AN4��C�#m REQUI9R��EBU�#��n6�$Tk�2$����zя #�& \^�APPR� C� ~0�
$OPEN�OCLOS�St���	i�
��&' 䂟MfЩ���W"-_MG�7CB@�A����BBRK@N�OLD@�0RTMCO_5ӆp1J��P�������������6��1��@ )!�#�(G� �����'<��+#PATH''@!@6#@!�<#� � '��1SCA���6IN��UCJ�[1� -C0@UM�(Y ��# �"�����*���*��� �PAYLOA~J{2LؠR_AN^�3L��91�)1AR_F2LSHg2B4LO4�!F7�#T7>�#ACRL_�%��0�'�$��H��.��$HA�2FLEX���J!�) P �2�D߽߫���0��* :����z� FG]D����z���%�F1]A�E�G4�F�X�j�|���BE���� ��������(��X�T *�A���@�XI�[�m�$\At�T$g�QX<�=� ��2TX���emX���� ���������������+	�J>+ ��-�K]o|�٠AT�F�4�ELFPѪsj�J� *� JEmgCTR�!�ATN���vzHAND_V�B.��1��$, M$8`F2Av����SWu	#-� $$M*0.�]�W�lg��PZ����A@��� 1����:AK��]AkAz��LTN�]DkDzPZ G��C�ST_K�lK�N}DY��� A ����0��<7]A<7W1@�'��d�@g`�P��������" 91B$. M�2D�%"��H����ASYIMj%0�� j&-��-W1�/_�{8� �$ �����/�/�/�/ 3J<�:9�/�89�D_VI�v����V_UNI�ӛ��cD1J����╴�W<�� n5Ŵ�w=4��9��?H�?<�uc�4�3�2%�H���/�j�L�0�DIzuO��q�k�>0 �`
��I��A��#���@�ģ���@���IPl� �1 � /�M�E.Qp��9�ơT}�PT�;pG �+ �Gt� ���'��T��0 $DU�MMY1��$P�S_�@RF�@  tG b�'FLA@ �YP(c|��$GLB_TP�ŗ����9 P�q��2 XX� z!ST9�� �SBRM M21_�V�T$SV_E�R*0O�p����CL�����AGPO��f�G�L~�EW>�3 4\H �$YrZr!W@�x�A1+�A���"t	""�U&�4 8`yNZ�"�$GI�p7}$&� -� �Y�>�5 LH {���}$F�E��NE+AR(PN�CF��%P�TANC�B	!JO�G�@� 6.@?$JOINTwa?p�d�MSET>�7 E x�E��HQtpS{r���up>�8� ��pU.Q?�� LOCK_FOV06���oBGLV�sGLt�TEST_XM� N3�EMP������_�$U&@%�w`#24� Y��5��2�4d��3��CE- ���� $KAR�QM>��TPDRA)�����VECn@��I�U��6��HEf�T�OOL�C2V�DR�E IS3ER6���@ACH� 7b?Ox �Q�29Z��H I�  @$�RAIL_BOX�Ewa�ROBO���?��HOWW�AR�1�_�zROLMj��:qw�jq�� �@ O_Fkp!G d�l>�9��W �R O8B: h�@�c�OU�	;�Һ�3ơ�r�q_�_$PIP��N&`�H�l�@��#@CORDEDd�p >�f�fpO�� < 7D ��OB⁴s d���Kӕ���qwSYS�ADR���f��TCHt� 7= ,8`ENo��1Ak�_{�-$Cq,B�e�VWVA��>� �  &��P�REV_RT��$EDITr&VSHWRkq�֑ &RJ:�v�D��JA�$~�a$HEAD�h6�� �z#KE:�E�CPSPD�&JKMP�L~��0R*PF��?��1%&I��5S�rC�pNE; �q��wTICK�C��M��1<�3HN���@ @� 1Gu�!_�GPp6��0STY'"xLO��:�2l2�?�A t 
m G�3%%$R!{�=��S�`!$��w`��������Pˠp6SQU���E��u�TERC��0��TSUtB ����hw&`gw�Q�)�pO����@IZh��{��^�PR�0kюB1XPU���Eg_DO��, XS�K~�AXI�@���UR�pGS�r� ^0��&��p_) �ET��BPm��o��0Fdo��0A|���R�h���a;�SR�Cl>@P��b_� yUr��Y��yU��yS�� yS���UЇ�U���U�� �U�]��Ul[��Y�bXk�]Cm������YRSC�� D �h�DS~0��Q�S�P���eATހ���A]0,2N�ADDR�ES<B} SHIyF{s��_2CH����I��=q�TV
srI��E"���a�C*e�
��
;�VW�AN��F \��q��0l|\A@�rC�_B"R�{zp�ҩq�TXS�CREE�Gv��1TINA���t�{����A�b?�H T1�ЂB�����I���A��BE�y RRO�������� B��D��UE4I �g�!p�9S��RSM]0�GUNEX(@~Ƴ�j�S_S�ӆ��Á։�ģ��ACY�0� [2H�pUE;�J�¸���@GMT��L�ֱ�A��O	�BB�L_| W8���K ���0s�OM��L1E/r��� TO!�s��RIGH��BRD<
�%qCKGR8л��TEX�@����WIDTH�� �B[�|�Z<��I_��Hi�� L 8K���_�!=r���R:�_���Yґ��O6q�M�g0紐U��h�Rm��LUMh��FpGERVw��P����`�N��&�GEKUR��FP)�)� �LP��(RE%@�a)�ק�a�!��f �5*�6�7�8Ǣ#B@�É@���tP�fW��S@M�USR�&�O <����U8�Qs�FOC)��PRI;Qm� :����TRIP�m�SUN����Pv��0���f%��'���@�0 �Q����AG ��0T� �a>q�OS�%�RPo���8�R/�A�H�L4����	U¡�SU�g��¢�5��OFF���T��}�O�� 1�R�����S�GU�N��6�B_S�UB?���,�SRT�N�`TUg2��mCO9R| D�RAUrPE�yTZ�#'�VCC���	3V AC36�MFB1f$c�PG� �W (#��ASTEM�����0�PE��T3G�X y�\ ��MOVEz�<���AN�� ���|M���LIM_X�� 2��2��7�,�����0ı�
��VF�`EӐ� }��04Y��IQB�7���5S��_Rp� 2��� WİGp+@��}СP��>3�Zx ����3���A�ݠCZ�DRID���ѡVy08�90� De�MY_UBYd���6��@��!��X��GP_S��3��L�K�BM,�$+0DE�Y(#EX`�����U/M_MU� X����ȀUS�� ���G0`PACI���а@ ��:��:,�:����CRE/�3qL�+���:[��TARG"��P�r��R<��\ d`��A��$�	4��AR��SW2 ��-��@Oz�%qA(7p�yREU�U�01�Z,�HK�2]g0��qP� N� �E9AM0GWOR��ާMRCV3�^ U���O�0M�C�s�	���|�REF _���x(�+T� �� �������3_RCH4(a�P�Ѐ��hrj�NA�5��0�_ ��2����L@��n�@@OU~7w6���Z��a2[��R1E�p�@;0\�c�a�'2K�@SUL��]2��C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��PQ5I�]7q�}�Tg`�4D`�0.`0�APg_HUC�5SA��CMPz�F�6�5�5
�0_�aR��a�1Ir\!X�9|"GFS��_ad ��M��0p�UF_x��B� �ʼ,RO��Q��'��6��UR�3GR�`.��3IDp���)�D`�;��A��~�IN��H{D���V@AJ���S͓UWmi=�0����TYLO*�5�����bt m+�cPA� �cCACH�vR�UvQ���Y��p�#CF�I0sFR�XT���Vn+'$HO����P!A 3�XBf�(1 ���$��`VPy� ^b_S�Z313he6K3he1�2J�eh chG�chW�A�UMP�j��IM5G9uPAD�ii�IMRE�$�b_SIZ�$P����0 ��ASYNBUF��VRTD)u5tqΓ?OLE_2DJ�Qu�5R��C��U��vPQ�uECCUlV�EMV �U�r�WVIsRC�aIuVTPG����rv1s��5qMPL�Aqa��v�V0�c���� CKLAS��	�Q�"��d  ��ѧ%ӑӠ@}¾�$8�Q���Ue |�0!�rSr�T�#0! 񕠄r�iI��m�vK�B�G��VE�Z�PK�= �v�Q�&�_HO|�0��f � >��3�@Sp�SLOW�>�RO��ACCaE���!� 9�VR�#0���p:���AD���F��PAV�j�� D����M_B"���^�'JMPG ��g:�#E$SSC��x&�HvPq��hݲvQS�`rqVN��LEXc�Gi T`�sӂ��Qn�FLD �DEsFI�3�02���:��VP2�Vj�� �A��V�4[`MV_PIs��t�0��A�@��FI��|�Z��Ȥ�����A���A���~�GAߥ1 LO9O��1 JCB����Xc��^`�#PLANE��R��1F�c�����pr�M� [`�噴��S����f����Af� �R�Aw�״tU��p�RKE��d�VAN�C�A���� k���ϲ�BR_AA� l��2� ��p8�#��m h�@��BO K�$������kЦ�0OU&A�"A�
�p�pSK�TM@FV{IEM 2l �8�P=���n <<���dK�UMMYK1�P��`D�Ȧ��CU��#AU��wo $��TITᱟ$PR����O�P���VSHIyF�r�p`J�`�Qsԙ�fOxE$� _R�`U�#����s ��q������G�"G��޵'�T�$�SCO{D7�CNTQ i�l� >a�-�a�;�a�H�a�V���1�+�2u1���D����  .� SMO�Uq�Ӳa�JQ�����a_��R[�r�n�*@L�IQ�AA/`�XVR���s�n�TL���Z7ABC�t�t�tc�
L�ZIP��Yu���LVbcLn"z���MPCFx�Mv:�$�� ���?DMY_LN����8���@y�w Ђ(a\�u� MCM�@Cbc�CART_�DP~N� $J71D��=NGg0S�g0�BUXW� ��U�XEUL|B yX���	������x 	���m��YH�Db  y� 80���0EIGH�3n�?(� H��9��$z ���|�,����$B� Kd'���_��L3�RVS�F8`���OVC�2@'�$|�>P&��
q�4��5D�TR�@ �9Vc��SPHX��!�{ ,� *<��$R�B2 2 ����C!�  ��� V+L�b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/ ?�/�/V(7%3@/R/ d/v/�/6?�/�/�?�?@�?O4OOION;4]? o?�?�?�?SO�?�?�O�_�O0_Q_8_f_N;5 zO�O�O�O�Op_�O_ o8o�_MonoUo�oN;6�_�_�_�_�_�oo %o4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8����� Ǐ=�_�n���R���şx��ڟN;G � џ�
�� ��?���W�i�{����� ��ï�.�������A��dW�<�N�|� ������Ŀֿ�ޯ� ��0�B�_�R�d�� �϶������������ �*�L�^��rτ�
� �����������&�p8�J�l�~� `ҟ @�з��������-����&�,� ��9�{�����a��� ������������A 'Y����� ����a#�1�
��N;_MO�DE  ��S ��[�Y�AB���
/\/*	|/��/R4CWORK_{AD�	�T1/R  ���� ��/� _INTVA�L�+$��R_O�PTION6 ��q@V_DAT�A_GRP 2,7���D��P�/~? �/�?�9��?�?�?�? OO;O)OKOMO_O�O �O�O�O�O�O_�O_ 7_%_[_I__m_�_�_ �_�_�_�_�_!ooEo 3oioWoyo�o�o�o�o �o�o�o/e S�w����� ��+��O�=�s�a� ������͏���ߏ� �9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_T�IM����� SC�R ��Ƙ_��5�;#U!P"�1!��� �?E�W�i�{����� .�ïկ�����'(+~�T"2F��"�dR�I�Y��2�o+@a얿����)�u�� k0ϴ��_; ��  T� �� �2�D�)�T D��Q�zόϞϰ��� ������
��.�@�R߀d�v߈ߚ�/V凷�����߽���R�;�o ��W�p��
�t���Diz$� �0 � �T"1!�� ����������� ����*�<�N�`�r� �������������� &8J\n�� ������"4FX ��࿁� ������/` 4�=/O/a/s/�/�/�/@�/�/�/�!!/ �0޲ k�ݵu�0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ ok$o6oHo Zolo~o�o�o�o�o1/ �o�o 2DVh z�/5?����� ���&�8�J�\�n� ��������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	���-�?�Q�c�u��� ���`Ò�ϯ��� �)�;�M�_�q�����@����˿ݿ� �����3� ���&2�,��	1234�5678v�h!�B!��2�C
h���0�ϵ��� �������!�3�9ѻ� \�n߀ߒߤ߶����� �����"�4�F�X�j� |�h�K߰��������� 
��.�@�R�d�v��� ����������� *<N`r��� ����&�� J\n����� ���/"/4/F/X/ j/|/;�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�/�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ �?L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o=_�o�o�o�o �o�o 2DVh�z�����h� �����u�o.�@�R����Cz  B���   ���2�&� � _�
~���  	�_��2�Տ����_�%p������ďi� {�������ß՟��� ��/�A�S�e�w��� ������N������ +�=�O�a�s������� ��Ϳ߿���'�9�DK�_������<v��_��$SCR_G�RP 1
�� �� t{ ��� ���	 �����������������_������)�a�����&�DE� �DW8���l�&�G��CR-35iA� 9012345�67890��M�-20��8��C�R35 ��:�
������������� ��:֦�Ӧ�G���&������	��]�o������:���#H���>�����������&���ݯ:� �j����g������B�t����������9A����  @�`���@� ( ?��=��Ht�P
��F?@ F�`z� y������ � $H��Gs^p��B��7� �/�0//-/f/Q/ �/u/�/�/�/8���P�� 7%?����"?W?x-2?<���]?� H�1�?t�ȭ7��������?-4A , �&E@�<�@G�	B-1 3OZOlO-:�HA�H�O�O|O P�B(�B�O�O_���EL_DEFAU�LT  �����`SHOTSTR#]JA7R�MIPOWERFOL  i�/UYToWFDO$V /U�RRVENT 1�����NU �L!DUM_E�IP_-8�j!?AF_INE#P�_�-4!FT�_->��_;o!��`o ��*o�o!RPC_OMAIN�ojh�vo��o�cVIS�oii���o!TPpP�U�Ydk!
�PMON_PROXYl�VeZ�2r��]f��!R?DM_SRV��Y9g�O�!R��k���Xh>���!
�`M���\i���!R�LSYNC�-9�8֏3�!ROS̽_-<�4"��!
�CE4pMTCOMd���Vkn�˟!	��OCONS̟�Wl����!��WASR�C��Vm�c�!N��USBd��XnR� ��Noӯ�������!���E��i�0���WR�VICE_KL �?%�[ (%SVCPRG1��D-:Ƶ2ܿ�˰3�D	�˰4,�1�˰5T�DY�˰6|ρ�˰7�� ��˰�����9����ȴf�!�˱οI�˱ ��q�˱ϙ�˱F��� ˱n���˱���˱�� 9�˱��a�˱߉�� 7߱��_������ ��)����Q���� y��'���O���� w������� ��˰��İd�c�� ����=( as^����� �/�/9/$/]/H/ �/l/�/�/�/�/�/�/ �/#??G?2?k?V?}? �?�?�?�?�?�?O�? 1OCO.OgORO�OvO�O �O�O�O�O	_�O-_��_DEV �Y��MC:5X��`GTGRP �2SVK ��bx 	� 
 ,�PK 5_�_�T�_�_ �_o�_'o9o o]oDo �ohozo�o�o�o�o�o �o5{�_g� �������� �?�&�c�u�\����� ��Ϗ���J\)��� M�4�q���j�����˟ ݟğ��%���[� B��f������ٯ�� �����3��W�i�P� ��t���ÿ���ο� ��A�(�e�L�ί�� RϿ��ϸ������ � �O�6�s�Zߗߩߐ� �ߴ������'�~ϐ� ]���h������ �������5��Y�@� R���v���������@� 	��?&cu\ ������� �;M4qX�� �����/�%// I/[/B//f/�/�/�/ �/�/�/�/�/3??W? �L?�?D?�?�?�?�? �?O�?/OAO(OeOLO �O�O�O�O�O�O�O�O�_"Ud �NLy�6 * 		S=>��+c"_�VU@Tn_Y_B����B�2�J�j�~Q´~_g_�_�Q%�JOGGING��_�^7T(?VjZ��Rf��Y��A�/e�_%o7e�Tt�] /o�o{m�_�o�m?Qi �o�o;)Kq%��o�}os�� ����9�{`�� )���%���ɏ���ۏ �S�8�w��k�Y��� }���ş���+��O� ٟC�1�g�U���y��� ����'����	�?� -�c�Q���ɯ����w� ��s����;�)�_� ����ſOϹϧ����� ����7�y�^ߝ�'� ��ߵߣ�������� Q�6�u���i�W��{� ������=��M��� A�/�e�S���w����� �������=+ aO������u� ��9']� ��M����� �/5/w\/�%/�/ }/�/�/�/�/�/=/"? 4?�/?�/U?�?y?�? �?�??�?9?�?-OO =O?OQO�OuO�O�?�O O�O_�O)__9_;_ M_�_�O�_�Os_�_�_ o�_%oo5o�_�_�o �_[o�o�o�o�o�o�o !coH�o{� �����; �_ �S�A�w�e������� я���7���+��O� =�s�a������П� ����'��K�9�o� ������_���[�ɯ�� �#��G���n���7� ��������ſ���� a�Fυ��y�gϝϋ� �ϯ�����9��]��� Q�?�u�cߙ߇ߩ��� %���5���)��M�;� q�_���߼��߅��� ����%��I�7�m��� ����]����������� !E��l��5� ������_ D�we��� ��%
//��� =/s/a/�/�/�/��/ !/�/??%?'?9?o? ]?�?�/�?�/�?�?�? O�?!O#O5OkO�?�O �?[O�O�O�O�O_�O _sO�Oj_�OC_�_�_ �_�_�_�_	oK_0oo_ �_co�_so�o�o�o�o �o#oGo�o;)_ Mo����o� ���7�%�[�I�k� ���������ُ� ��3�!�W���~���G� i�C����՟���/� q�V������w����� ���ѯ�I�.�m��� a�O���s�������߿ !��E�Ͽ9�'�]�K� ��oϑ�����Ϸ� ���5�#�Y�G�}߿� ����m���i������ 1��U��|��E�� ��������	���-�o� T������u������� ����G�,k���_ M�q���� ���%[I m���	��� //!/W/E/{/��/ �k/�/�/�/�/	?? ?S?�/z?�/C?�?�? �?�?�?�?O[?�?RO �?+O�OsO�O�O�O�O �O3O_WO�OK_�O[_ �_o_�_�_�__�_/_ �_#ooGo5oWo}oko �o�_�oo�o�o�o C1Sy�o��o i�����	�?� �f�x�/�Q�+���Ϗ �����Y�>�}�� q�_�������˟��� 1��U�ߟI�7�m�[� }����ǯ	��-��� !��E�3�i�W�y�ϯ ��ƿ�������� A�/�eϧ���˿UϿ� Q���������=�� dߣ�-ߗ߅߻ߩ��� �����W�<�{��o� ]���������/� �S���G�5�k�Y��� }��������������� C1gU���� ��{����	? -c���S�� ����/;/}b/ �+/�/�/�/�/�/�/ �/C/i/:?y/?m?[? �??�?�?�?? O?? �?3O�?COiOWO�O{O �O�?�OO�O_�O/_ _?_e_S_�_�O�_�O y_�_�_o�_+oo;o ao�_�o�_Qo�o�o�o �o�o'ioN` 9������ A&�e�Y�G�i�k� }�����׏���=�Ǐ 1��U�C�e�g�y��� �֟���	���-�� Q�?�a���ݟ��퟇� �ϯ��)��M��� t���=���9���ݿ˿ ��%�g�Lϋ��� mϣϑϳ�������?� $�c���W�E�{�iߟ� �߯������;���/� �S�A�w�e������ �������+��O� =�s������c����� ������'K��r ��;������ �#eJ�}k �����+Q"/ a�U/C/y/g/�/�/ �//�/'/�/?�/+? Q???u?c?�?�/�?�/ �?�?�?OO'OMO;O qO�?�O�?aO�O�O�O �O__#_I_�Op_�O 9_�_�_�_�_�_�_o Q_6oHo�_!o�_io�o �o�o�o�o)oMo�o A/QSe�����%{,p�$S�ERV_MAILW  +u!��+q~�OUTPUT��$�@�RV� 2�v  $�� (�q�}��SA�VE7�(�TOP1�0 2W� d? 6 *_�π(_������#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u����������Ͽݷ��Y�P��'�FZN_C�FG �u�$�~����GR�P 2�D� ?,B   A[�+q�D;� B\���  B4~�R�B21��HELL���u��j�k��2�����%RSR �������
�C�.�g� Rߋ�v߈��߬������	���-�?�Q��  �_�%Q���(_���,p��⦼�ޖ�g�2,pd�����HK 1�� ��E�@�R� d��������������� ��*<e`r����OMM ������FTOV_�ENB�_���HO�W_REG_UI��(�IMIOFW�DL� �^�)WAIT���$V�1�^�NTIMn���VA�|_)_UNIT����LCTRY�B�
�MB_H�DDN 2W� 2�:%0 �pQ/ �qL/^/�/�/�/�/�/��/�/�"!ON_ALIAS ?e�	f�he�A?S?e? w?�:/?�?�?�?�?�? OO&O8OJO�?nO�O �O�O�OaO�O�O�O_ "_�OF_X_j_|_'_�_ �_�_�_�_�_oo0o BoTo�_xo�o�o�o�o ko�o�o,�oP bt�1���� ���(�:�L�^�	� ��������ʏu�� � �$�Ϗ5�Z�l�~��� ;���Ɵ؟����� � 2�D�V�h�������� ¯ԯ���
��.�ٯ R�d�v�����E���п ���ϱ�*�<�N�`� r�ϖϨϺ���w��� ��&�8���\�n߀� �ߤ�O���������� ��4�F�X�j�|�'�� �����������0� B���f�x�������Y� ��������>P bt����� �(:L�p ����c�� / /$/�H/Z/l/~/)/ �/�/�/�/�/�/? ?�2?D?V?]3�$SM�ON_DEFPR�O ����1 �*SYSTEM*�0m6RECAL�L ?}9 (� �}4xcop�y fr:\*.�* virt:\tmpback�1�=>147.87�.149.40:�17680 �29{8 �65172]?,O+M}5�5a�?�?`�6�?O�O�O}9�4�s:orderf?il.datML_O�uO�O_*_}0�2mdb:JO�O�1�O_ �_�_8C�?QO^_t_�_ o)o<O�_�_rOo�o �o�O�OU_p_�o% 8_J_�on_ ���_ Io[o�_~�!�4oFo �jo������o�oM �oz���0Bݏf ��������S��v� �����>�ϟ�t�� ������ΏW�r���� '�:�կ������� ��K�]���#�6� ǿٿl����ϡϴ�Ư O��|���2�D��� h��ϋߝ߰�¿U�� x�	��.�@���d������,�<��N�ou�tput\tes�t_serverw.pcC�: o��� _�62791424:3597y� 
��������a�w�+� ��-�?�Z�c�u��� *��P������� ;�L^q�&9� K���o������� d��/"/5�� k��/�/��V/� {/??���������/ �?�?/AS�/�/�? O���?��?O�O �O=/�/]Os/�O_(_ �/�O�O�/_�_�_92�B??Q8_writ�e\?n;�_o%o83A<�_�Yread�_n; o�o�o�?�?RO�Iyo 
/OAO�oeO�o+���}�$SNPX�_ASG 2�����q�� P 0 '�%R[1]@g1.1��y?��s%�!��E�(�:�{� ^�������Տ��ʏ� ��A�$�e�H�Z��� ~���џ����؟�+� �5�a�D���h�z��� ��ů�ԯ���
�K� .�U���d�������ۿ ������5��*�k� N�uϡτ��ϨϺ��� ���1��U�8�Jߋ� nߕ��ߤ�������� ��%�Q�4�u�X�j�� ������������;� �E�q�T���x����� ������%[ >e�t���� ��!E(:{ ^������/ �/A/$/e/H/Z/�/ ~/�/�/�/�/�/�/+? ?5?a?D?�?h?z?�? �?�?�?�?O�?
OKO .OUO�OdO�O�O�O�O �O�O_�O5__*_k_ N_u_�_�_�_�_�_�_ �_o1ooUo8oJo�o�no�o�o�d�tPAR�AM �u��q �	��jP��d9p�ht���pOFT_KB_?CFG  �c�u��sOPIN_SI/M  �{vn���p�pRVQS�TP_DSBW~�r"t�HtSR �Zy � & �ROB195_?SERV M����vTOP_O�N_ERR  �uCy8�PTN �Zuk�A�4�RING_PR��D��`VCNT?_GP 2Zuq�!px 	r��ɍ`���׏��wVD���RP 1�i p �y��K�]�o����� ����ɟ۟����#� 5�G�Y���}������� ůׯ�����F�C� U�g�y���������ӿ ��	��-�?�Q�c� uχϙϫ��������� ��)�;�M�_�qߘ� �ߧ߹��������� %�7�^�[�m���� ����������$�!�3� E�W�i�{��������� ������/AS ew������ �+=Ovs �������/ /</9/K/]/o/�/�/ �/�/�/�/?�/?#? 5?G?Y?k?}?�?�?�?��?�?�?�?OO)�P�RG_COUNT�8v�k�GuKBEN�B��FEMpC:t}O_�UPD 1�{T  
4Or�O�O �O__!_3_\_W_i_ {_�_�_�_�_�_�_�_ o4o/oAoSo|owo�o �o�o�o�o�o +TOas��� �����,�'�9� K�t�o���������ɏ ۏ����#�L�G�Y� k���������ܟן� ��$��1�C�l�g�y� ��������ӯ����	� �D�?�Q�c������� ��ԿϿ����)��;�d�_�q�=L_IN�FO 1�E[�@ �2@����������� ��B��  B4 �4�*�@HYSDEBU)GU@�@���d�If�SP_PASSUE�B?x�LOG � ���C���Qؑ�  ��A��?UD1:\��U���_MPC�ݵE&�$8�A��V� �A�?SAV !��������X���SV�Z�TEM_TIM�E 1"���@k 01@<X��X���E�����$T1S�VGUNS�@VE'��E��ASK_?OPTIONU@�Et�A�A+�_DI���qOG�BC2_GRP 2#�I�����?@�  C���<K~o�CFG %z�Ɠ� �����` ��	�.>dO� s������� *N9r]�� �����/�8/#/\/n/v$Y,�/Z/ �/�/H/�/?�/'?? K?]�k?=�@0s?�?�? �?�?�?�?O�?OO )O_OMO�OqO�O�O�O �O�O_�O%__I_7_ m_[_}__�_�_�X�  �_�_oo/o�_SoAo co�owo�o�o�o�o�o �o=+MOa �������� �9�'�]�K���o��� ������ɏ���#��_ ;�M�k�}�������� ß�ן��1���U� C�y�g����������� ����	�?�-�c�Q� s����������Ͽ� ���)�_�Mσ�9� �ϭ�������m��� #�I�7�m�ߑ�_ߵ� ������������!� W�E�{�i������ ��������A�/�e� S�u�w����������� ��+=O��sa ������� 9']Kmo� ������#// 3/Y/G/}/k/�/�/�/ �/�/�/�/??C?�� [?m?�?�?�?-?�?�? �?	O�?-O?OQOOuO cO�O�O�O�O�O�O�O __;_)___M_�_q_ �_�_�_�_�_o�_%o o5o7oIoomo�oY? �o�o�o�o�o3! CiW���� �����-�/�A� w�e����������я ���=�+�a�O��� s�������ߟ͟��o �-�K�]�o�ퟓ������ɯ���צ��$�TBCSG_GR�P 2&ץ��  �� 
 ?�  6� H�2�l�V���z���ƿ��������(�_d�E+�?��	 HC���>Ǚ��G����C��  A�.�e�q�C;��>ǳ33��SƑ/]϶�Y��=Ȑ� ?C\  Bȹ��{B���>����,P���B�Y�z��L�H�0�$����J�\�n�����@�Ҿ�� �������=�Z�%�7���?3������	V3.00~.�	cr35��	*����
��������� 3��4��   {�CT��v�}��J2�)�������CFG [+ץ'� *�V�����I����.<
� <bM�q��� ����(L7 p[����� �/�6/!/Z/E/W/ �/{/�/�/�/�/.�H� �/??�/L?7?\?�? m?�?�?�?�?�? OO $O�?HO3OlOWO|O�O ����Oӯ�O�O�O!_ _E_3_i_W_�_{_�_ �_�_�_�_o�_/oo ?oAoSo�owo�o�o�o �o�o�o+O= s�E���Y�� ���9�'�]�K�m� ������u�Ǐɏۏ� ��5�G�Y�k�%���}� ����ßşן���1� �U�C�y�g������� ӯ������	�+�-� ?�u�c���������� Ͽ���/�A�S��� ��qϓϕϧ������ ��%�7�I�[���m� �ߑ߳������߷�� 3�!�W�E�{�i��� �����������A� /�e�S�u��������� ������+a O�s��e��� ��'K9o] ������� #//G/5/k/}/�/�/ [/�/�/�/�/�/?? C?1?g?U?�?y?�?�? �?�?�?	O�?-OOQO ?OaO�OuO�O�O�O�O �O�O___M_�e_ w_�_3_�_�_�_�_�_ oo7o%o[omoo�o Oo�o�o�o�o�o! 3�o�oiW�{� ������/�� S�A�w�e�������я �������=�+�M� s�a���������ߟ� �_	���_ן]�K��� o�������ۯɯ��� #���Y�G�}�k��� ��ſ׿������� �U�C�y�gϝϋ��� ���������	�?�-� c�Q�s�u߇߽߫��� �����)��9�_�M� ����/����i���� ��%��I�7�m�[��� ���������������� EWi{5�� ������A /eS�w��� ��/�+//O/=/ _/a/s/�/�/�/�/�/ �/?'?��??Q?c?? �?�?�?�?�?�?�?O �?5OGOYOkO)O�O}Op�O�O�O�N  �@�S V_R��$TBJOP_G�RP 2,�E��  ?��V	-R4S.;\=��@|u0{S~PU >��U�T @�@LR	� �C� �Vf?  C���ULQ�LQ>�33�U�R�����U�Y?�@=��ZC��P�����R��P  Bȸ�W$o/gC��@g��dDb�^�㙚eeao�P&ff~�e=�7LC/kFaB o�o�P��P��efb-C�p�B�^g`�d�o�PL�P�t<�eVC\ � �Q@�'p�`��  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�anaaF`C�;�`L�w��aQoxp�x�p:���XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb����X �	��1��)�W��� c������������ 󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSc7r35QT*�QT��A�� E��'E�i�F�V#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG��G#
�D���E'
E�MKE���E��ɑE�ۘE���E���F���F��F���F(��F�5��FB��F�O��F\��F�i��Fv��F���vF�u�<#�
<t����ٵ=�_��V �R�p�V9�~ ]ESTPARtp��HFP*SHR\�A�BLE 1/;[$%�SG�� �W�
G�G�G� WQG�	G�
G�GȖ�QG�G�G�ܱv�'RDI~�EQ�ϧ� ��������W�O_�q�@{ߍߟ߱���w�S]�CS !ڄ������ ������&�8�J�\� n������������� ] \�`��	��(�:� ����
��.�@�w��NUM  �EUEQ�P	P ۰�ܰw�_CFG �0��)r-PIMEBF_TTb��CSo�,VERڳ-B�,R 11;[' 8��R�@� �@&  ��� ����//)/;/ M/_/q/�/�/�/�/�/ ?�/?J?%?7?M?[? m?>�@�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_��_l_�Y@c�Y�MI_CHAN�8 c cDBGLV��:cX�	`�ETHERAD �?f�\`���?�_uo�oQ�	`RO�UTV!	
!��d�o�lSNMAS�KQhcba255.uߣ'9ߣY��OOLOFS_D�Ib��U;iORQCTRL 2		�Ϸ~T��� ��#�5�G�Y�k�}� ������ŏ׏�����.��R�V�PE_�DETAI/h|zP�GL_CONFI�G 8�	����/cell/$�CID$/grp1V�̟ޟ�������o?�Q�c�u����� (���ϯ������ ;�M�_�q�����$�6� ˿ݿ���%ϴ�I� [�m�ϑϣ�2����� �����!߰���W�i� {ߍߟ߱�%}F��� ����/�A�C�i�H�Eߞ�������� ��?��.�@�R�d�v� ������������� ��*<N`r� ������& 8J\n��!� ����/�4/F/ X/j/|/�//�/�/�/ �/�/??�/B?T?f? x?�?�?+?�?�?�?�? OO�?>OPObOtO�O��O�O���Us�er View ���}}1234567890�O�O�O�_#_5_=T�P��]_���I2�I:O�_�_�_@�_�_�_X_j_�B3�_ GoYoko}o�o�o o�op^46o�o1CU�ovp^5�o������	�h*�p^6 �c�u����������ޏp^7R��)�;�M� _�q�Џ��p^8�˟ ݟ���%���F�L�� lCamera�J���� ����ӯ���E~�� !�3��OM�_�q��������y  e��Yz��� 	��-�?�Q���uχ� ��俽���������>��e�5i��c�u߇� �߽߫�d������P� )�;�M�_�q��*�<� �i���������)� ��M�_�q�������� ��������<�û��= Oas��>��� �*'9K] f�Q������ �/�%/7/I/�m/ /�/�/�/�/n<�� ^/?%?7?I?[?m?/ �?�?�? ?�?�?�?O !O3O�/<׹��?O�O �O�O�O�O�?�O_!_ lOE_W_i_{_�_�_FOXG9+_�_�_oo(o :o�OKopo�o)_�o�o@�o�o�o ��	g�0�oM_q��� No����o�%�7� I�[�m�&l�n�� Ə؏���� ��D� V�h���������ԟ 柍�g�ڻ}�2�D�V� h�z���3���¯ԯ� ��
��.�@�R���3u F�鯞���¿Կ��� ���.�@ϋ�d�vψ� �ϬϾ�e�w���U�
� �.�@�R�d�ψߚ� ������������*� ��w���v���� ����w�����c�<� N�`�r�����=�w�� -�����*<�� `r�������x���  �� 1CUgy��������    -/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_�i_�  
��( � �%( 	 y_�_�_�_�_�_�_ o	o+o-o?ouoco�o�o�o�Z* � Q&�J\n ������o��� 9�(�:�L�^�p�� �������܏� �� $�6�}�Z�l�~�ŏ�� ��Ɵ؟���C�U�2� D�V���z�������¯ ԯ���
��c�@�R� d�v�����᯾�п� )���*�<�N�`ϧ� ���ϨϺ������� �&�8��\�n߀��� �߶���������E�"� 4�F��j�|���� ��������e�B� T�f�x����������� ��+�,>Pb ���������� (o�^p� ������ /G $/6/H/�l/~/�/�/ �/�//�/�/?U/2?�D?V?h?z?�?�/�`@� �2�?�?�?�3��7�P��!frh�:\tpgl\r�obots\m2�0ia\cr35?ia.xml�?;O MO_OqO�O�O�O�O�O�O�O ���O_(_ :_L_^_p_�_�_�_�_ �_�_�O�_o$o6oHo Zolo~o�o�o�o�o�o �_�o 2DVh z������o� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟�ݟ��&�8� J�\�n���������ȯ ߟٯ���"�4�F�X� j�|�������Ŀ־�8�.1 �?@8?8�?�ֻ� ֿ�3�5�G�iϓ�}� ���ϳ��������5߀�A�k�U�wߡ߿���$TPGL_OUTPUT ;�!��! �� ������,�>�P�b� t����������� ��(�:�L�^�p������������2345678901�� �������"�� BTfx��4�@����
}$ L^p��,>� �� //$/�2/Z/ l/~/�/�/:/�/�/�/ �/? ?�/�/V?h?z? �?�?�?H?�?�?�?
O O.O�?<OdOvO�O�O �ODOVO�O�O__*_ <_�OJ_r_�_�_�_�_ R_�_�_oo&o8o�_ �_no�o�o�o�o�o`o �o�o"4F�oT�|����\��} �����0�B�T�e��@������� ( 	 ��Џ��� ���<�*�L�N�`� ��������ޟ̟�� �8�&�\�J���n��� ������ȯ���"�������*�X�j�F��� ��|�¿Կ��C���� ��3�E�#�i�{�忇� ��S����������/� ��S�e�߉ߛ�y߿� ��;�������=�O� -�s���ߩ��]��� �����'����]�o� �����������E��� ��5G%W}�� ����g��� 1�Ug	w�{ ��=O	//�?/ Q///u/�/��/�/_/ �/�/�/�/)?;?�/_? q??�?�?�?�?�?G? �?O�?OIO[O9OO �O�?�O�OiO�O�O�O !_3_�O_i_{__�_�_�_�_�_�R�$T�POFF_LIM� >�op:�y�mqbN_SV`�  l�jP_�MON <6�)dopop2l�a�STRTCHK �=6�f� bVTCOMPAT-h��afVWVAR �>Mm�h1d ��o �oop`b�a_DEFPRO�G %|j%R�OB195_SE�RV	�j_DIS�PLAY`|n"rI�NST_MSK � t| ^zINqUGp�o tLCK�|�}{QUICKMEyN�dtSCRE�p�6��bt_scdt�q��b*��ST�jiRACE_CFG ?Mi��d`	�d
?��u�HNL 2@"|i����k r͏ ߏ���'�9�K�]��w�ITEM 2A��� �%$12�34567890<����  =<��П<��  !���p��=��c��^� ���������.���R� �v�"�H�ί��Я� �����*�ֿ���r� 2ϖ�����4�޿�ϰ� ��&���J�\�n���@� ��d�v��ς������ 4���X��*��@�� ���ߨ������� T���x������l� �������,�>�P��� ����FX��d���� ��:�p" ��o����� F6HZt~�� N/t/�/��// /2/ �/V/?(?:?�/F?�/ �/�/j?�??�?�?R? �?v?�?QO�?lO�?�O �OO�O*O|O_`O _ �O0_V_h_�Ot_�O_ _�_8_�_
oo�_@o �_�_�_Lodo�_�o�o 4o�oXojo3�oN�o r��o��s��S�B���z� 3 h��z ��C�:y
 P�v�]���~�UD1:\������qR_GRP� 1C��� 	 @Cp���@$��H�6�l�Z��|� ����f���˟���ڕ?�  
���<� *�`�N���r������� ޯ̯��&��J�8�Z���	�u�����s�SCB 2D� �����(�:��L�^�pς��|V_C�ONFIG E��� ��~����Ϝ�OUTPUT� F���� ��5�G�Y�k�}ߏߡ� �������������#� 6�H�Z�l�~���� ����������%�9� K�]�o����������� ������"�5GY k}������ �1CUgy �������	/ ,?/Q/c/u/�/�/ �/�/�/�/�/??(/ ;?M?_?q?�?�?�?�? �?�?�?OO$?7OIO [OmOO�O�O�O�O�O �O�O_ O2OE_W_i_ {_�_�_�_�_�_�_�_ oo._AoSoeowo�o �o�o�o�o�o�o ������!�6oew� �������� +�=�0oa�s������� ��͏ߏ���'�9� J�]�o���������ɟ ۟����#�5�F�X� k�}�������ůׯ� ����1�C�T�g�y� ��������ӿ���	� �-�?�P�c�uχϙ� �Ͻ���������)� ;�L�^�q߃ߕߧ߹� ��������%�7�I� Z�m��������� �����!�3�E�V�i� {��������������� /AR�d�w� �������+=O2u���k}gV�Kv� ���////A/S/ e/w/�/�/�/`�/�/ �/�/??1?C?U?g? y?�?�?�?`�?�?�? 	OO-O?OQOcOuO�O �O�O�?�O�O�O__ )_;_M___q_�_�_�_ �O�O�_�_oo%o7o Io[omoo�o�o�o�_ �o�o�o!3EW i{����o�� ���/�A�S�e�w� ������������ �+�=�O�a�s����� ����̏ߟ���'� 9�K�]�o��������� ȟۯ����#�5�G��Y�k�}�������ž��$TX_SCRE�EN 1G�g�}i�pnl/��gen.htmſ�*�<��N�`ϽPan�el setupd�}�dϥϷ����������ω�6�H�Z� l�~ߐ�ߴ�+����� ��� �2�߻�h�z� ������9�g�]�
� �.�@�R�d������ ����������}��� <N`r��; 1��&8� \��������QȾUALRM_�MSG ?��� �Ȫ-/?/p/ c/�/�/�/�/�/�/�/�??6?)?Z?%SEoV  -�6�"ECFG Iv��  ȥ�@�  A�1  w B�Ȥ
 [? ϣ��?OO%O7OIO�[OmOO�O�O�G�1G�RP 2J�; 0Ȧ	 �?�O �I_BBL_NO�TE K�:T?��lϢ��ѡ�0RDEFP�RO %+ (%N?u_Ѡc_�_�_�_ �_�_�_o�_o>o)o�boMo�o\INUSER  R]�O�o�I_MENHIS�T 1L�9  �( _P��'�/SOFTPAR�T/GENLIN�K?curren�t=menupage,69,1�opBTfx �(
~253/������p)�~381,23�L�^�p��	#�71�̏ޏ�����q0��uedi�t(rROB195t0RV��Y�k�}����(�7H�ԟ���
����)q10X�j� |�����/���4H�ܯ � ��5R�`q|oB� T�f�x������1�ƿ ؿ���� ϯ�D�V� h�zόϞ�-������� ��
�߫Ͻ�R�d�v� �ߚ߬�;�������� �*��N�`�r��� ��7�I�������&� 8�#�\�n��������� ��������"4F ��j|����S ��0BT� x�����a� //,/>/P/�t/�/ �/�/�/�/�/o/?? (?:?L?^?I��?�?�? �?�?�?�?�/O$O6O HOZOlO�?�O�O�O�O �O�OyO_ _2_D_V_ h_z_	_�_�_�_�_�_ �_�_o.o@oRodovo o�o�o�o�o�o�o �o*<N`r�o? ������ 8�J�\�n�����!��� ȏڏ��������F� X�j�|�����/�ğ֟ �������B�T�f� x�����+�=�ү��� ��,���P�b�t���������z�$UI_�PANEDATA 1N���ڱ�  	��}/frh/�cgtp/wid�edev.stm� ?_fonts?ize=14��!��3�E�W� )pr�imYς�  } } �itree�� �Ͼ�������[��)� �M�4�q߃�jߧߎ� ���������%�7���[�7��� � {���&���flex���6�e���������J�ual��"��ϧ�X�j�|� ����G����������� BT;x_�@�����i� ݰ ܳ7�-?Qcu ����0���� /!/3/�E/i/P/�/ t/�/�/�/�/�/?? ?A?(?e?w?^?�?  �?�?�?OO+O~? OOaO��O�O�O�O�O �OFO_�O'_9_ _]_ D_�_�_z_�_�_�_�_ �_o�_5o�?�?Eo}o �o�o�o�o�o*o�onO 1CUgy�o� ������	�-� �Q�8�u���n����� Ϗ�Tofo�)�;�M� _�q�ď����˟ݟ ���z�%�I�0�m� T�������ǯ����� �!��E�W�>�{��  ���ÿտ����^� /�Aϴ�e�wωϛϭ� ��&������� �=� $�a�s�Zߗ�~߻ߢ� ��������%�]� o�����
���N� ���#�5�G�Y���}� ��v����������� ��1UgN�r��4�F����"4FX)�}�� l�����/j '//K/2/D/�/h/�/ �/�/�/�/�/�/#?5?�?Y?��C�=��$U�I_POSTYP�E  C�?� 	 e?�?��2QUICKME/N  �;�?�?��0RESTORE� 1OC��  �*default�;�  REEVI�EW:LDUAL��?mmenup�age,107,�1fO�O�O�O�OrD�ozF381,26,22�O_ _2_D_ mF_j_|_�_�_�_ EAL?�_�_G_�_"o4o FoXojoo�o�o�o�o �oyo�o0B�_ Oas�o���� ���,�>�P�b�t� �������Ώ���� �����L�^�p����� 7���ʟܟ� ���$� 6�H�Z�l��!����� ������� �2�կ V�h�z�����A�¿Կ����
��=SCK@N� ?�=uw1sc+@u2K�U3K�4K�5K�6K��7K�8K��2USE1R-�2�D�ksMì�U3��4��5��6���7��8���0NDO_CFG P�;�� ��0PDATE� ���N�one�2��_IN_FO 1QC�@��10%�[���Iߊ� m߮��ߣ�������� ��>�P�3�t��i����<-�OFFSET T�=�ﲳ$@ ������1�^�U�g� ��������������� $-ZQcu����?�
����UFRAME  �����*�RTOL_�ABRT	(�!E�NB*GRP �1UI�1Cz  A��~��~���������0UJ�9MSKG  M@�;N�%8�%��/�2V7CCM��V�ͣ#+RG�#Y�9���/j����D�BH�Yp71C���37f11?�C0�$MRf�2_�*S�Ҵ�	����~XC5G6 *�?�6����1$�5���A@v3C��. ��8�?��OOKOx1�FOsO�5�51���_O�O�� B����A2�DWO�O7O _�O8_#_\_G_�_k_ }_�__�_�_�_�_"op�OFoXo�%TCC�#A`mI1�i������� GFS��2a�Z; �| 2345678901�o �b�����o��!5�a�4BwB�`56 �311:�o=L �Br5v1�1~1�2��}/ ��o�a��#�G Yk}�p����� ��ُ�1�C�U�6� H���5�~���ߏ����	���4�dSELE�C)M!v1b3�VIRTSYNC��� ���%�SIO�NTMOU�������F��#b������(u� FR:\H�\��A\�� ��� MC��LOG���   UD1懦EX����' B@ �����̡m��̡  OB�CL�1�H� ��  =	 1�- n6  -#������[�,S�A��`=��͗���ˢ��TRAIN�⯞b�a1l�
0d�$j�T2cZ; ( aE2ϖ�i��;�)� _�M�g�qσϕϧ���������	��F�ST�AT dm~2@�zߌ�*j$i߾���_GE�#eZ;�M`0�
� 02���HOMIN� f����� ~�(����БC�g�X����JMPERR 2=gZ;
  ��*j l�V�7���������� ����
��2�@�q�d��v�B�_ߠRE� h\Wޠ$LEX��iZ;��a1-e��VMPHASE  5�r�c�!OFF/��F�P2n�j�0R�㜳E1@���0ϒE1!1?s33�����ak/�kxPk䜣!W�m[�䦲 �[����o3;� [i{ ����/� O�?/M/_/q/��/ ��//�/'/9/�/=? 7?I?s?�/�?�/�/�? �??Om?O%O3OEO �?�?�O�?�O�O�?�O �O�O__gO\_�OE_ �O�_�O�O/_�_�_�_ oQ_Fou_�_|o�o�_ �oo�o�o�o�o;oMo ?qof-�oI�� ���7�[P� ��������ˏ� �!�3�(�:�i�[�ŏ�g�}������TD__FILTEW�n��g �ֲ:���@� ��+�=�O�a�s��� ������֯������0�B�T�f�x���S�HIFTMENU� 1o[�<��% ��ֿ����ڿ���� I� �2��V�hώ��π�ϰ�������3�
��	LIVE/SN�AP'�vsflsiv��E����/ION * Ub�h�menu~߃���߰�ߣ���p���a	����E�.�50�s�P�@� ��AVɠB8z�z��}���x�~�P�� � ���MEb�Կ�<�0���MO���q���z�WA�ITDINENDb������OK1N�OUT���SD���TIM����o�G���#���C����b������RELE�ASE������TM��������_AC�T[�����_DA�TA r��%�L����xRDIS�b�E�$XVR��s���$ZAB�C_GRP 1t��Q�,#�0�2\���ZIP�u'��&����[MPCF_G 1v�BQ�0�/� w�<�ɤ� 	�Z/  85�/�/H/�/l$?��+�/�/ �/?�/�/???r?�?  �D0�?�?��?�?�?�;���x��]hYLIND�֑y� ���? ,(  *VOgM�.�SO�OwO�O�M  i?�O�O^PO1_�OU_ <_N_�_�O�_�_�__ �_�_x_-ooQo8o�_0�o�oY&#2z� ���oC�e?@a?>N|�oq����q�A�$DSPHER/E 2{6M��_� ;o���!�io|W� i��_��,��Ï��� Ώ@��/�v���e�؏ ��p����������6ZZ�� �N