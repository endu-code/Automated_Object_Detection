��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�� RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DIS�� /�SMB�	"�BCJ@"CI2�AIP6EXPS�!�PAR�� �Q{CL�
 <(yC�0�SPTM�E�� PWR��X�V<�Ro l5�d�!�"%�7�ICC��%� kfR�0leP�� _DLV��YNo3 <oNbX�_�P~#Z_IND9E
C�`OFF� ~UR�iD��c�   t �!N�`MON�%sD�.&rHOU�#EWA,v�Sq;vSqJvLOCAܗ Y$N�0H_[HE���@I"�/ 3 $ARPhz&�1F�W_\ d�I!F�`;FA�D�k01#�HO_� I�NFO�sEL	%# P K  !k0�WO` $A7CCE� LVZk:�2H#ICE�L��  �$�s# ����k���
��
�`�K`SQi��V �5|�I�0A�Lh�z�'0 ��
�
��F����V �܅w�$� 2ċ��w������� č��!r�Z���4����Ċ!14�7.87.224�.20h�S���9A6����܁܁3�_{p�_  ċ� bfh.ch̟ �1�C�U�g�y�����௯��ӯ^�� _FL�TR  ��π V]� ������n��nxč2n��rSH��PD 1ĉ � P!
robstation֯.՚!k�.�Q� ſ��������޿?� �c�&χ�JϫϽπ� �Ϥ����)���M�� "߃�Fߧ�j��ߎ��� ����%���I��m�0� ��T��x������ ��3���W��{���P� ��t����������� ��Sw:�^� �����= �a$Zׯ$ _L��A1��x!1!.�ğP�1�Q255.%�S���2��E  �//*/<&3F/�@� l/~/�/�/<&4�/��50�/�/??<&5 6?��0\?n?�?�?<&6�?�%@�?�?�?
O�1�?P��MY�� MY���c��� Q�	 �VN<�O�O_�O�+_=_O_"_s_�_NP d_�_�_�_�_�_o!o@3o�_Woio{oVNLo M��o�l�oAo
�.@U}iRC�onnect: �irc\t//alertsE��� �Pu����1��C�UуP_R8�d��H�~�������Ə ؏���� �2�D�V�"S$���8�(p���@�o͟ߟ��QA8��d�A�B4��j��h9�Q+��@DM�_�A+��SMB 	X�8%ğVO�߯���_CLN�T 2
X� 4C�ɯ0��l�c�B� T���x���Ͽ����� �)�;��_�q�Pϕ���MTP_CTR/L ��%���� �dc���ߋ��?�*��c߳l��N���@�{�Vߵ�Ƥ��������ѓC��UST�OM {����}�@ }�DTCWPIPu�{��h\�E�TEL�{�z�A���H!Ta��t�çrobl�olr�  ���!KCL���|F��!CRT���������!CGONS&����n+���