��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�5J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA� R�!R�	� � $TIT�!$I��N �D@d�Dd �Dc@�D5�FU6�F7�F8�F9�G0�G�GJA�E�GbA�E
�G1�G1�G �F�G�2�B!SBN_C�F>"
 8F CN�V_J� ; �"�!_�CMNT�$F�LAGS]�CH�EC�8 � ELL�SETUP ރ $HO30IO��0� %�SMAC{RO�RREPR�X� D+�0��R{�T� UTOBACK�U�0 ��)DEVIC�CT	I*0�� �0�#��`B�S$INTE�RVALO#ISP�_UNI�O`_D�O>f7uiFR_F�0AIN�1���1<c�C_WAkda^�jOFF_O0N�DEL�hL� ?aA�a1b?9a�`C#?��P�1E��#s�ATB�d��MO<� �cE D [�M�c��^qREV��BILrw!XI�� QrR  �� OD�P�q$NO^PM�Wp�t�r/"�w� �u��q�r�0D`S �p E RD_E��pCq$FSSB�n&$CHKBD_[SE^eAG G�"$SLOT_�H�2=�� V�d�%��3���a_ED�Im   � )�"��PS�`(4�%$EP�1�1$�OP�0�2�a�p_�OK�UST1P_�C� ��d��U �PLACI4!�Q�4�<( raCOMM� ,0$D����0�`���EOWB BIGALwLOW� (Kt�"(2�0VARa�Є@�2aI�L�0OUy� ,Kvay��P9S�`�0M_O]�����CCFS_UT~p0 "�1�3�#�ؗ`X"�}R0 � 4F IMCM�`O#S�`��upi �_�p�B}�a����M/ h�pI?MPEE_F�N���N���@O��r�DQ_�~�n�Dy�F�����_�r0 � T� '��'�DI��n0"��p�P��$I���� w�CF�t X� �GRP0��M=qN�FLI�7��0UI�RE��$g"� SW�ITCH5�AX_�N�PSs"CF_L�IM� � �0EED��!��PqP�t�`PJ_dVЦMODEh�.Z`�P|Ӻ�ELBOF�  ������p� ���3���� FB/��0t�>�G� �� �WARNM�`/�p�qP��n�NST� �COR-0bFL{TRh�TRAT�P�T1�� $ACC�1a��N ��r$OcRI�o"V�RT�Ps_S� CHG�0I��rT2��1�I��T�I1��� x i#�Q�.�HDRBJ; C�Q�2L�3L�4L�5�L�6L�7L� N�9�s"��O`S <�F +�=�O��#92��L�LECy�"MULTI�b�"N��1�!t���0T�� �STY�"�R`�=l��)2`����*�`T  |� �&$��۱m�a�P�̱�UTO��:�E��EXT����pÁB���"2� (䈴![0������p<�b+�� "D" ���ŽQ��<煰kc!(�9�#���1��ÂqM�ԽP��" '��3�$ L� E���P<��`A�$JO�Bn�T���R��IG3�% dK��������<���\��+�Y�6�C�O_M��& �t�pFLܐBNG AgTBA� ��� M��
�!��p� �q���0�P[`��O�'[���0tna*����"J��_R���C�DJ��IdJk�D�%C�`�Z���0���P_�P��@ ( @�F RO.��&�t�I9T�c�NOM�
�����Sp�P`T)"w@���Z�P�d���RA�0��2b"�����
$T����MD%3�T��`U31��ʩp(5!HGb�T1�*E�7�c�KAb�pWAb�cA4#YNT��>�PDBGD�� *(��PUt@X���W���AX��a��ewTAI^cBUF���0!+ � l7n�PIW�*5 P�7M�8M�9
0�6}F�7SIMQS@�>KEE�3PAT�n�^�a" 2`#�"�L�64FIX!, !���!d��D�2Bus�=CCI�:FPCH�P:BAD�aHCEhAOGhA]HW�_�0>�0_h@�f�Ak���F�q@\'M`#�"�DE3�- l�p3G��@FSOES]FgHBSU�I�BS9WtB��. `{ ��MARG쀜���FACLp�SLEWx aQe�ӿl�xRMC�/�>\pSM_JBM��� �QYC	g�e��Д�0 ā�CHNv-�MP�$G� �Jg�_� #��1_3FP$�!TCuf!À�#�����d�#a��V`&��r�a;�fJR�о�rSEGFR�PIyO� STRT��N��cPV5���!41�r��
r>İ�b��B�O�2` +�[���,qE`�,q�`y�Ԣ}t��yaSCIZ%���t�vT�s�� �z�y,qRSINF}Oбc���k��`��`�`L�ĸ T`7�gCRCf�ԣCC/��9��`a�uah�ub�MIN��uaDs�#�G�D�YC��C�����e`�q0��� �EV�q�F�_�eF��N@3�s�ah��Xa+p,�5!�#1�!VS�CA?� A��s1�"!3 ��`F/k� �_�U��g��]��C�� �a�s�o�R�4� ����N����5za�R�HANC���$LG��P�f1$f+@NDP�t�AR5@�N^��a�q���c��M�E�18���}0��RAө�AZ 𨵰�%O��FCTK��s`�"�S�PFADIJ�OJ�ʠ�ʠ��� <���Ր��GI�p�BMP�d�p�Dba���AES�@	�K�W_��BAS�� �G�_5  M�I�T��CSX[@@�!6�2�	$X���T9�{sC��N�`�~P?_HEIGHs1;�gWID�0�VT #ACϰ�1A�Pl�<���EXPg���|���CU�0MMENuU��7�TIT,AE�%)�a2���a��8 P� a�E�D�E.`��PDT���REM.��AU�TH_KEY  H������ �b�O	�<��}1ERRLH� ��9 \� �q-�OR�DB�_ID�@l �P�UN_O��Y�$�SYS0��4g�-�I�E�EV�#q'�OPXWO�� �:j�O$SK7!f21&��Td�TRL��; ��'AC�`��ĠI�ND9DJ.D��_Ė�f1��f���PL�A�RWAj���SD�A��!+r|�ПUMMY9d�F�1E0d��'���J�<��v}1PR� 
3��POS��J�= l�$V$�q/ �L~�>���ܠK�?����CJ�@\����ENE�@T���A���_�REC�OR��BH z5 O�@=$LA�>$~�r2�R��`�q�U�`�_Du��0RO�@V�T[�Q�U��������! }У�PAU�S���dETURN,��MRU�  ;CRp�EWM�b�A�GNAL:s2$L�A�!?$P�X�@$P�y A �Ax�C0 #ܠDO�`X�k�W�v�q�GO_AWAY��MO�ae���]�C�SS_CCSCB� C �'N��CERI��гJ`u�QA�0�}��@�GAG� R�0�`��0{`��{`OF�q��5��#MA��Xf���&шLL�?D� �$���s�U�D)E%!`���O�VR10W�,�OR�|�'�$ESC_|$`�eDSBIOQ���l ��B�VIB&� �c,�����f�=pSSW���f!�VL��PL���AORMLO
��`�����d7%SC �bA1LspH�MPCh @�Ch �#h �#h 5�UU���C�'�C�'�#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$4�C��P3Wұ46$V7OLT37$$`�*�^1��$`O1*��$o��0RQY���2b4�0DH_TH�E����0SЯ4�7ALPH�4�`���7�@Q �0�qb7�rR�5�88� ×���"(��Fn�MӁ!VHBPFUAFLQ"Dt�s�`�THR��@i2dB�����G(��PVP�����������Ђ�H2�B�E�C�E�CPSu�Y@��Fb3��� H�(V�H:U�G�
X0��FkQw�[�Na�'B���C INHBcFILT���$��W �2�T1�[ ��$h���H YАAF�sDO��Y�Rp� fg �Q�+�c5h�Q�iSh�QPL���Wqi�QTMOU�#c�i�Q \��X�gmb��vi�h�biAi�fI�aHIG��ca	xO��ܰ��W�"vAN-u!��	#�AV�H!Pa8�$P�ד#p�R_:�A(�a��B�N0�X�MCN���f1[1�qVE�p��Z2;&f��I�QO�u�rx�wGldDN{G|d��a!F>!�9��aM:�U�'FWA�:�Ml��� X�Lu��$!����!l��ZO����0%O�lF��s�13�DI�W� @��Q���_��!�CURVA԰0rC	R41ͰZ�C<�r�H� v���<�`U�<�(�f�CH�QR3�S���t0���Xp�VS_�`�$ד�F��ژ�����҈NSTCY?_ E L����A1�t�1��U��24�2B�NI O7�����އDEVI|� �F��$5�RBT.xSPIB�P���#BYX����T���HNDG��G HC tn���L�@�Q�C���5��Lo0� H��閻�FBP�{tFE{�5�t�h�T��I�DO���uPMCS�v>�f�>�t�"HOTSWt�`s�?ELE��J T���e�2��2d5�� O� ��HA7�E��344�0&?��A�wK �� MDL�/ 2J~PE��	A���s��tːÈ�s�J ÆG!��rD"�ó���L��\�TO��W�	���/��SLAV�wL  �pINPڐp���`%ن_CFd�M� $��ENU��OG��b�ϑ]զP�0`ҕ�]�IDMA�Sa��\��WR�#��"]�VE\�$a�SKI�STs�H�sk$��2u���J�À�����	��Q���_�SVh�EXCLU8MqJ2M!ONL��D�Y��|�PE ղI�_V�APPLYZP��HID-@Y�r��_M�2��VRF�Y�0��r�1�cIO#C_f�� 1����2��O��u�LS���R�$DUMMY3ҏ!���S� L_TP/Bv�"���AӞ�>ّ N ����RT_u�� � ��G&r[�O{ D��P_BA�`g�3x�!F ҁ�_5���H��da�tA�P�� P� $�KwARGI8��� q�2O[���_SGNZ�Q �8~P/�/PIGNs�l�$�^ sQANNUN�@�T<0�U/�ߴ�LAzp]	�Z�d~�EF�wPI�@ R @��F?IT�	$TOTA%��d����!�M�NI�Y�S+���E�A�[�
DAYS\�A�Dx�@��	� �EFF_AXI?�1TI��0zCOJA� �ADJ_RT+RQ��Up��<P$�1D �r5̀Ll�T�p? ]P�"p��pmtpd��V 0w��G��������S�K�SU� ��CT�RL_CA�� }W�TRANS��6PIDLE_PW����!��A�V��V�_�l�V �D�IAGS���X�w /$2�_SE�#TAC���t!�!0�z*@��RR��vPAh���p ; SW�!@�!�  ��ol�U��foOH��PP� ���IR�r��BRK'#��"A_Ak���x  2x�9ϐZs2��%�l�W�pt*�x%RQ�DW�%MSx�t5A�X�'�"��LIFEgCAL���10��N�1{"�5Z�3{"dp�5�ZU`}�MOTNr°Y$@FLA�c�ZOVC@p�5HE|	��SUPPOQ�ݑAq� Lj (C�1S_X6�IEYRJZRJWRJ�0TH�!UC��6�XZ_AR�p��YM2�HCOQ��Sf6�AN��w$�ICT�E�Y `��CACHE�C9�M��PLAN��UFFIQ@�Ф0<�1�	��6
���MS�W�EZ 8�KEgYIM�p��TM~�SwQq�wQ#���貟OCVIE� �[; A�BGL��/�}�?� 	�?��D�\p�ذST��!�R� �T� �T� �T<	��PEMAIf�ҁ���_FAUL��]�Rц�1�U��� �TRE�?^< $Rc�u�S�% IT��BU!FW}�W��N_� 'SUB~d��C|��8Sb�q�bSAV�e�b�u �B��� �gX�^P �d�u+p�$�_~`�e�p%yOTT����s�P��M��OtT�LwAX � ��X~`9#�c�_G�3
�YN_1�_�D��1 �U2M���T��F��H@ g�`� 0p��Gb-s7C_R�AIK���r�t�RoQ�u7h�q'DSPq��rP��A�IM�c6�\����s2��U�@�A�sM*`I�P���s�!D��6�T!H�@n�)�OT�!6��HSDI3�ABSC���@ Vy���� �_D�CONVI�G���@3�~`	F�!�pd��psq�SCZ"���sMER�k��qFB��k��pEiT���aeRFU:@�DUr`����x�CAD,���@p;cHR�	A!��bp�ՔՔV+PSԕC���	C��p��ғSp�_cH *�LX� :cd�Rqa�| ����W� �U��U��U�	�U�TOQU�7R�8R�9R���0T�^�1k�1x�1���1��1��1��1*��1ƪ2Ԫ2^�k�U2x�2��2��2��U2��2��2ƪ3Ԫ%3^�3k�x�3���To���3��3��3ƪ94Ԣ�EXTk!0�d <� 7h�p�6�p�O��p����NaFDR^Z$eT^`V��Gr����䂴2REMr� Fj��BOVM�z�A�TROVٳDT�`-�MX<�I�N��0,�W!IND�KЗ
w�׀�p$DG~q36��P�5�!9D�6�RIV���2��BGEAR�IO�%K�¾DN�p��J��82�PB@�CZ_MCCM�@�1��@U���1�f ,②a?� ���PI�!?I�E��Q���a�m���g� _0Pfq�g RI9ej�k!UP?2_ h � �cTD�p���! a����i�w�C�ri T��P�b�`�) OG���%���p��IF�I�!�pm�>��	�P�T�",���MR2>��j ��Ɛ +"����\��������P$�B`x%��_ԡ��"�_���� M���߾��DGCLF�%D7GDY%LDa��!5�6�ߺ4��M���S�k��� T�sFS#p�Tl P���e�qP�p$EX_���1M2��2j� 3�5��G ����m ��Ѝ�SW��eOe6DEBUG����%GR���pUn�#BKU_�O1'�7 �@PO�I�5�5MS��OYOfswSM��E�b��@�0�0_E �n �p C��T�ERM�o� E�D�ORI+�p~� �SM_���b�q�2O ��TA�r����UP�Rs� 9-�1�2n$�' �o$SEG,*> E�LTO��$US]E�pNFIAU"�4�e1���#$p$UFR���0ؐO!�0��f��OT�'�TAƀ�U�#NST�PA�T��P�"PTHJ�����E�P rF�V"ART�``%B`�abU!�REL:�aSHF�T��V!�!�(_SH"+@M$���� ��@rN8r����OVRq�N�rSHI%0��UN�= �aAYLO�����qIl����!�@��@ERV]��1�?:�� �'�2��%��5�%��RCq��EASYM�q�EV!WJi'��}�AE���!I�2��U@D@��q�%Ba��
5Po�X�0�p6OR�MY�& `GR��t2b5�n� � ��UPa�Uu� Ԭ")���TO�CO!S�1POP@ ��`�pC�������YOѥ`REPR3�b�aO�P�b�"eP�R�%WU.X1��e$7PWR��IMIU�2sR_	S�$VIS���#(AUD���Dv" ;v��$H���P__ADDR��H�AG�"�Q�Q�QБR~p\Dp1�w H� SZ� a��e�ex�e��cSE��r��HS���MNvx ����%Ŕ��OL����p<P��-��AC�ROlP_!QND_�C��ג�1�T �RO�UPT��B_�VpQ�A1Q�v��c_��i ���i��hx��i���il��v�ACk�IOU���D�gfsu^d�gy $|�P_D��xVB`bPRM_�b{e�ATTP_א�Haz (��OBcJEr��P��$���LE�#�s`{ � ��u�AB_�x�T~�S�@�D�BGLV��KRL~�YHITCOU�[BGY LO a�TEM��e�>�+P'��,PSS|�P�JQUERY_FLA�bG�HW��\!a|`�u@�PU�b�PIO��"�]�ӂ/dԁ=d�ԁ�� �IOLN���}����CXa�$SLZ�$INoPUT_g�$IPb#�P��'���SLvpa~��!�\�W�C-��B$�IO�pF_AuSv��$L ��w �F1G�U�B0m!a���0HY���ڑ��RS:��UOPs� `������@[�ʔ[�і"�[PP�S�IP�<�іI�2�da�t�IP_MEM�B��i`� X��I1P�P�b{�_N�`����R�����b�SP��p$FOC�USBG�acs�{UJ�Ƃ �  �� o7JOG�'�D�IS[�J7�cx�J8�7� Im!�)�7_LAB�!�@��A��APHIb��Q�]�D� J7Jx\���� _KEYt�� �KՀLM�ONa���$X�R��ɀ��WATC�H_��3���ELĉ�}Sy~���s� ĮЮ!V�g� �CTaR3򲓥��LG�D�� �R��I�
LG_SIZ���JŰq IƖ�I�FDT�I H�_�jV�GȴI�F� %SO���q �Ɩ���v��ƴ��K�S����w��k�N�����E��\���'�*�UȢs5��@L>�4�DAUZ�EA�pՀ�Dp��f�GH�BiᢐBO}O��� C����PIT���� ��R{EC��SCRN��ⵖD_p�aMARGf�`��:���T�$L���S�s��W�Ԣ��Iԭ�JGMO�MN3CH�c��FN��R��Kx�PRGv�UF���p0��FWD��H]L��STP��V��+���Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*�a2�8����Gh�0P!O��������M8�Ģv��EX��TUIv�	I��(�4�@� t�x�J0J�~�P���J0��N�a�#ANA8��O"�0VAIA��d�CLEAR�6DCS_HI"�/c�5O�O�SI��9S��IGN_�vp�q�uᛀT�d� DE�V-�LLA �°B�UW`��x0T6<$U�EM��ŁR����0�A�R���x0�σ�a�@OSU1�2�3�a�`� �ࠜh�ApN%-���-�IDX�D	P�2MRO��Գ!�+ST��Rq�Y{b!� �$E&C`+��p.&A&,���`� L��ȟ%P ݘ��T\Q�UE�`�U�a��_ � ��@(��`�����# �MB_PN@ R`r�y�R�w�TRIN��P��BASS�a	6gIRQ6�MC(��� ��CLD�P�� ETRQLI`��!D�O9=4FLʡh2�Aq3zD�q7���LDq5[4q5ORG �)�2�8P�R��4�/c�4=b-4�t� ��rp[4*�L4q5S�@T�O0Qt�0*D2FRCLMC@D�?�?RIAtr,1ID`�D� d1���RQQprpDS3TB
`� �FᆻHAXD2���G�LE�XCES?R`�BMhPa���BD4+2��A�q`�`�F_�A�J�C[�O�H� K���� \���bTf$�� ��LI�q�SRE�QUIRE�#MOx�\�a�XDEBU��__N�ML� M�� �p���P�c��AA,1N��
Q�q�0/�&���-cDC��B�sIN�a?�RSM�Gh� N#B��N�ae��bPST9� �� 4��LOC�R�I���EX�fAN�G��A,1ODAQ䵗�@$��9�ZMF�����f��"��p�%u#ЖVSUP�%��aFX�@IGGo�� �rq�"��@1��#B��$���p%#�by��rx���vbPD'ATAK�pE;�������M��*� tV�`MD�qI��)�v� �t�A�wH�`��t�DIAE��sANSAW��th���uD���)�bԣ(@$`� PCU_�V6�ʠ�d&�PLOr�$`�R���B���B�p������RRR2�E��  ��V�A/A ?d$CALI�@��	G~�2��!V��w<$R�SW0^D�"��ABC�hD_�J2SE�Q�@�q_�J3M�
G�1SPH�,��@PG�n�3m�(u�3p�@��JkC��4�2'AO)IMk@{BCSKP^:ܔ9�wܔJy�{BQܜ��8���`_AZ.B���?�EL��YAOC�MP�c|A)��RT�j���1�ﰈ��@�1�������Z��S�MG��pԕ� ER�!���INҠACk�p����b�
n _�������D4�/R��DIU��C�DH�@
�#a�qc$V�Fc�$x�$���`@���b���̂�E�H ��$BELP����!A/CCEL���kA>°IRC_R�pG0��T!�$P)S�@B2L������W3�ط9� ٶPACTH��.�γ.�3���p�A_��_�e�-Br�`C���_MG�$DD��ٰ��$FW�@�p����γ칲��DE��PPA�BN�ROTSPEEu��O0���DEF>Q����$OUSE_��JPQP�C��JY����-A 6qYN�@A�L�̐��L�MOU�NG̭�|�OL�y�INCU��a�¢ĻB��ӑ�AENCS���q�B������D�IN�I`Y����pzC�VE��<���23_U ��b^�LOWL���:�O0��0�Di�B�P�Ҡ� ��PRC����M3OS� gTMOpp�@�-GPERCH  M�OVӤ ����� !3�yD!e�]�6�<�$� ʓAY���LIʓ�dWɗ��:p3�.�I�T3RKӥ�AY���� ?Q^�Y�m�b��`p�CQ�� MOM�B?R �0u��D���y�0�̂��DUҐZ�S_�BCKLSH_C Y���o�n��TӀ����
c��CLAL�J��A��/PKCH�KO0�Su�RTY�� �q��M�1�q_�
#c�_UMCP�	C����SCL���LMTj�_L�0X����E�� �� � ��m�h���6��PC����H� �P��2�CN@�"XT����CN_��N^C�kCSF����V6�����ϡjY��nCAT�SHs�����ָ1����֙���������P�A���_P���_ P0� e���O1u�$x�JG� P{#�OG|���TORQU(� p�a�~����Ry������"_W��^�����4Pt�
5z�
5I;I ;Iz�F�`�!��_8�1��VC��0�D�B�2�1�>	P�?�B�5JR�K�<�2�6i�DBL�_SM�Q&BMD`_sDLt�&BGRV4`
Dt�
Dz��1H_��8�31�8JCOSEKr�EHLN�0hK�5oDt� jI��jI<1�J�LZ1�51Zc@y��1MYqA�H�QBTHWMYTHE{T09�NK23z��/Rn�r@CB4VCBn�CqPASfaYR<40gQt�gQ4VSBt��RN?UGTS���Cq���a��P#���Z�C$DUu ��R䂥э2��Vӑ��Q�r�f$N	E�+pIs@�|� �	$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b��F�c�j�FR�VrhV�ghd��lV�jV�kV��kV�kV�kV�kV�iHrh�f�r�m!�x��kH�kH�kH�kH��kH�iOclOrhOT��nO�jO�kO�kUO�kO�kO�kO�F�F.bTQ���E��egS�PBALANCEl��RLE�PH_'USP衅F��F��FPFULC�3���3��E��1�l�UT�O_p �%T1T2t���2NW������ǡ��5�`�擳�T��OU���� INSsEG��R�REV���R���DIFH��1ٟ��F�1�;�OB��;C��2� �b~�4LCHWAR���;�ABW!��$MECH]Q�@k�q��AXk�P��IgU�i�� 
���!����7ROB��CRY�ͥ�&� �C��_�s"T � x $WEIGHh�F9�$cc�� Ih��.�IF ќ�LAG�K�8SK��K�BI�L?�OD��U��S	TŰ�P�; ���(�������
�Ы�<L��  2�`�"�/DEBU.�L&�n�=�PMMY9��qNA#δ9�$D&�ƪ�$��� Q   �DO_�A��� <	���~�H�L�BX�P�N�Ӣ+�_7�L�t�OH  ��� %��T����ѼT�����TgICK/�C�T1��%������N��c����R L�S���S��ž��PROMPh�E~� $IR� �X�~ ���!�MAI��0��j���_9�����t�l�R�0CO�D��FU`�+�ID�_" =�����G_�SUFF<0 h3�O����DO�� ِ��R��Ǔن�S���P�!{������	�H)��_FI��9��O�RDX� ����3�6��X�����GqR9�S��ZDTD����v�ŧ4 =*�L_NA4���|K��DEF_I[� K���g��_���i���0��š���IS`i  �萚����e��"��4�0i�Dg����D� O��LOCKEA!uӛϭ�0����{�u�UMz�K� {ԓ�{ԡ�{����}� ��v�Ա��g����� ��^���K�Փ����!w�N�P'���^����,`�W\�[R���TEFĨ ��OULOMB�_u�0�VIS�PITY�A�!O>Y�A_FRId��F(�SI���R��H����3���W�!W��0��0_,�EAS%��!�& �"���4p�G;穯 h ��7ƵC?OEFF_Om��H�m�/�G!%�S.��߲CA5����u�G�R` � � �$R� �X]�TME�$R�s�Z�/,)ËER�T;�:䗰��  ]�LL��S��_SV�($�~����@���� �"SETU��MEA��Z�x0�u���>��� � � �� ȰID�"���!�*��&P���*�F�'����)3��#�A��"�5;`*�ЧREC���!7�S�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I���0�MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X17ࡐMO�R�� H	�CU �A3�z�1Q�
��3���$��FV���2�SbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�N�HeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų7�=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	����y��=q�#}1� @�@;���MOE�RI#A��
N��X�s�f�\7���P�L}1�,RTv�m�A�TUSRBTRC_T(qR��B ������$ �Ʊ��,�~0� !D��`-CSALl`�`SA���]1gqXE�� �%���C��J�
�Ʊ�UP(4����PX���؆�q��3�w� ��PG�5� $SUB���������t�JMPWAI�TO��s��LOyCF8t�!D=�CVF	ь��y���R`�0��CC�_CTR�Q�	�I�GNR_PLt�D�BTBm�P��z�B�W)����0U@���I�G�a��Iy�TNL�N��Z�R]aK� N��B�0�PE�s���r܊�f�SPD}1� L	�A�`gఠ�S��CUN�{���]�R!��BDLY�2������PH_PK�E�~�2RETRIEt���2�b����FI��B� ����8� �2��0DBGL�V�LOGSIZ,$C�KTؑUy#u��D7�_�_T1@�E�M�@C\1A����R���D�FCHECKLK�R�P�0����@�&�(bLEc�" PEA9�T���P�C߰iPN�����ARh� 0���Ӯ�PO�B?ORMATTnaF��f1h���2�S��UqXy`	���PLBо�4�  rEI�TCH��{ 8P�L)�AL_ �# $��XPB�q� �C,2D�!��+2�J�3D��� T�pP�DCKyp��oC� _�ALPH���BE0WQo���� ��I��wp � �b@P�AYLOA��m�_�1t�2t���J3A�R��؀դ֏�laTWIA4��5��6,2MOMCP��������4���0BϐAD��������PUBk`R ��;���;�����z4��` I$PI \Ds�oӓ1yՕ�w�2��w�Z��I��I��I ���p����n���y��e`�9S)bT�SPEED� G��(�Е ��/���Е�`/�e��>��M��ЕSAM�P�6V��/���ЕMO�@ 2@�A��QP ���C��n��������� ��LRf`kb�ІE9h��EIN09��7S�.В9
yPy�G�AMM%S���D�$GET)bP�cD4]��2
�IB�q��I�G$HI(0;AH��LREXPA8)LWVM8@z)��g���C5�GCHKKp]�0�I_��h`eT��n�q���eT,���� ��$�� 1��iPI� RCH_�D�313\��30LE@�1�1\�o(Y�7 �t�_MSWFL �M��SCRc�7�@�&��ز%n�f�SV����PB``�'�!�B�sS_SAV&0ct5B3NO]�C\�C2^�0 �mߗ�uٍa��u����u:e;��1���8��D �P��������� )��b9��e�GE�3���V�2�LN m�� 7� �YL��Q
NQSRlbfqXG �P�RR#dCQp� $�S:AW70�B�B[�ȤCgR:AMxP�KCL �H���W�r�(1n�g�9M�!o�� �F�P@}t$WP�u�P r ��P5�R<�RC�R ��%�6�`��� ��qsJr X��OD�qZ�U�g�ڐ>D� ��OM#w�J?\?n?�?��?��9�b"�8�PuL]�_��� |� �X0��bf��qf��q`��ڏgzf��Eڐ� �Z��Fb�"ɐ�t��FdPB��PM��QU�� � 8�L�QCOU!h Q�THI�HOQBpH�YSY�ES��qU�E�`�"�O��� � �P�@\�UN����Cf�O�� P��Vu��!����OOGRAƁcB2�O�tVuITe �q:p/INFO�����{��qcB��OI�r�{ (�@SLEQS� �q��p�vgqS����� 4L�ENA�BDRZ�PTION�t�����Q���)�GCuF��G�$J�,q^r�� R����U�g���OS_ED������ �F��PK���E'NU�߇وAUT$1܅COPY�����n�00�MN���PR�UT8R �Nx�OU��$G[rf�@b_RGADJ���*�3X_:@բ$�����P��W��P��} ���)�}�EX�YCzDR�qRGNS.�9�F@r�LGO�#��NYQ_FREQ�R�W� �#�h�TsL�Ae#����ӄ �CcRE� s�IF�ᶕsNA��%a�_}Ge#STATUI`<e#MAIL������q t�������EwLEM�� �/0><�FEASI?�B ��n�ڢ�1�]� � I�p��Y!q]�Lt#A�ABM���E�pr<�VΡY�BASR҈Z��S�UZ��0�$q���RMS_TR;�qb ���SY��	�ǡ��$���>C��Q`	� 2� _�TM������̲��@ �A��)ǅ�i$D�OU�s]$Nj���P�R+@3���rGRIyD�qM�BARS �sTY@��OTO�Rp��� Hp_}�!����d�O�P/�� �s �p�`POR�s���}���SRV��),����DI&0T��Ѡ�� #�	�#�4!�5*!�6!�7!�8��q�F�2��Ep$VALUt��%��ֱ��>/��� ;�1ėq�����(_�AN��#�ғ�Rɀ(���T�OTAL��S��P�W�Il��REG#EN�1�cX��ks0(��a���`TR��R��_S� ��1ଃV �����⹂Z�E��p��q��Vr���V_Hƍ�DA�S����S_�Y,1�R4�S� AR��P2� ^�IG�_SE	s����å_�Zp��C_�Ƃ�EN�HANC�a� T ;�������GINT�.��@FPs^İ_OVRsP�`@p�`��Lv��o��7�p}��Z�@�SLG�
AA�~�25�	��Dd��S�BĤDE�1U�����TE�P���� !Y��
��J��$2�IL_M`C�x r#_��`TQ�`���q���'�BV�CF�P_� 0�M�	[V1�
V1�2�U2�3�3�4�4�
�!���� � m�A�2IN~VIB�P���1�2�2��3�3�4�4��A@-�C2���=p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KEEP_HNADD!�!`$^�j)C�Q�� �$��"	��#O�a_$�A�!K��#i��#REM�"�$��½%�!��(U}�e�$HPW�D  `#SBWMSK|)G�qU�2:�P	�COLLAB� �!K5�B�� 4��g��pITI1{�9p#>D� ,�@F�LAP��$SYNT �<M�`C6���UP_DLYAA�ErDELA�0ᐢmY�`AD�Q�p�QSKIP=E� i���XpOfPNTv�A�0P_Xp�rG�p �RU@,G��:I+�:IB1 :IG�9JT�9Ja�9Jn��9J{�9J9<��RA=s� X���4��%1�QB� NFLIC�s�@J�U�H�LwNO_H�0�"?��R�ITg��@_PAz�pG�Q� �K�
^�U��W��LV�d�NGRLT�0_q���O�  " ��OS��T_�JvA V	�APPR�_WEIGH�sJg4CH?pvTOR��vT��LOO��]�+�"tVJ�е�ғA�Q�UL�S�XOB'�'�
A`SJ2P���7�X�T�<a43DP=`Ԡ\"p<a�q\!�pRDC�ѮL� �рR��R�`� �RV��jr�b�RGE��*��cNFLG�a�Z���SsPC�s�UM_<`>^2TH2NH��P~.a 1� m`�EF11��� �lQ �!#� <�p3AT� g�S�&�Vr�p�t�Mq�Lr���HO�MEwr�t2'r��-?Qcu� Rt3'r������� tt4'r�'�9�K�]�o���
�5'r뤏��ȏڏ(�����6'r�!�3��E�W�i�{��7'r퀞���ԟ�����8'r��-�?�Q�c�u�R�uS$0�q�p�� sF��`�la�!`P�����`/���-�IO[M�I֠���1�R�pWE�� ���0Za*��� ��5��$DSB� GNAL���0Cxp��m`S2323�'� �~`��� / gICEQP��PEp̤�5PIT����OPyBx0��FLOW�@�TRvP��!U���CuU�M��UXT�A|��w�ERFAC��� U��ȳCHN��� tQ  _���>�Q$����OM���A�`T�P#UKPD7 A�ct�T���UEX@�ȟ�U E�FA: X"�1RSP�T�����T ���PPA�0o񩩕`EXP�IOS���)ԭ��_���%��C�WR�A��ѩD�ag֕`Ԧ?FRIENDsaC2�UF7P����TOO�L��MYH C2L�ENGTH_VT�E��I��Ӆ$�SE����UFIN�V_���RG9I�{QITI5B�ױXv��-�G2-�G�17�w�SG�X��_��UQQD=#���AS��d~C�`��q��_ �$$C/�S�`����� �0��>��VERSI� ��w�0�5���I��������AAV�M_Y�2 �� 0 � �5��C�O�\@�r� r�	 ����� ����������������
?�QY�BS���1���� <-������ 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO�jO|O�O�O�OiCC��@XLMT&��C��  ��DINp�O�A�Dq�EXE�HiPV_��ATQ�z
��LARMRECOV ��RgLMDG �*�5�OLM_�IF *�%�d �O�_�_�_�_j�_'o�9oKo]onm, 
 ��odb��o�o�o�o�^��$� z, A�   2D{�PPINFO u[ �Vw��������`������ �*��&�`�J���n�����DQ����
� �.�@�R�d�v����������a
PPLIC�AT��?�P���`Han�dlingToo�l 
� 
V8.30P/40Cp�ɔ_LI
88�3��ɕ$ME�
F0G�4�-

398�ɘ��%�z�
7D�C3�ɜ
�Non�eɘVr���ɞ@/6d� Vq?_ACTIVU�r�C죴�MODP����C�I��HGAP�ON���OU�P�1*��  i�m����Қ_�����1*�  �@��������Q����Կ�@�
������ ���5��Hʵl�K�HTTHKY_��/�M�S� ����������%�7� ��[�m�ߝߣߵ��� �������!�3��W� i�{���������� ����/���S�e�w� �������������� +�Oas�� �����' �K]o���� ����/#/}/G/ Y/k/�/�/�/�/�/�/ �/�/??y?C?U?g? �?�?�?�?�?�?�?�? 	OOuO?OQOcO�O�O �O�O�O�O�O�O__ q_;_M___}_�_�_�_`�_�_�_kŭ�TOp���
�DO_CLE�AN9��pcNM  !{衮o�o�o��o�o��DSPDgRYRwo��HI��m@�or���� �����&�8�J���MAXݐWdak�H�h�XWd�d���PLUGGW�Xgd���PRC)pB�`"�kaS�Oǂ2^DtSEGF0�K�  �+��o�or�������8���%�LAPOb� x�� �2�D�V�h�z��������¯ԯ�+�T�OTAL����+�U�SENUO�\� �e�A�k­�RGDI_SPMMC.����C6�z�@@Dr\�O�Mpo�:�X�_STRING 1	(��
�M!�S��
��_ITE;M1Ƕ  n�� ����+�=�O�a�s� �ϗϩϻ����������'�9�I/O SIGNAL���Tryout� ModeȵI�npy�Simul�ateḏOu�t��OVER�RLp = 100�˲In cyc�l�̱Prog� Abor��̱~u�Statusʳ�	Heartbe�atƷMH F�aul	��Aler�L�:�L�^�p�����������  ScûSaտ��-�?�Q� c�u������������� ��);M_q��WOR.�û�� ����+= Oas��������//'.PO ����M �6/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�?�?H"DEVP.�0d/ �?O*O<ONO`OrO�O �O�O�O�O�O�O__�&_8_J_\_n_PALT	��Q�o_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o�_GRIm�û9q �_as���� �����'�9�K��]�o�������'�R 	�݁Q����)�;� M�_�q���������˟ ݟ���%�7�I�ˏPREG�^����[� ����ͯ߯���'� 9�K�]�o����������ɿۿ�O��$AR�G_� D ?	����0���  	$�O�	[D�]D���O�e�#�SBN_C�ONFIG 
�0˃���}�CI�I_SAVE  �O�����#�TC�ELLSETUP� 0�%  O�ME_IOO�O�%?MOV_H���ώ��REP��J��U�TOBACK�����FRA;:\o� Q�o���'`��o��ҟ��� ��  f�o�����*�!�3�`��Ԉ��f���� ������o�{��&�8� J�\�n���������� ��������"4FX j|�������끁  ��S�YSUIF.SV� V T.TP �D MP 6.VD GIF PH�D_q��N}qS#��f�INI�P�o���c�MESSAG�����8�>�ODE_D�����z��O�0�c�PA�USM!!�0� �(73�U/g+(Od/�/x/�/�/�/ �/�/�/???P?>?�t?1�0$: TSK � @-��T�f�UP3DT��d�0
&�XWZD_ENB8����6STA�0���5"�XIS��UN�T 20Ž� �� 	 ���z��en�g�-���S�o�U@�	�H����tL�Oo��}Cw�g�^����.�O�O�O�O/_n2FMET߀2CM�PTAA��@��$A-�@����@���@����]5��5��(d5��P5��r�5F*5��338]SCRD�CFG 1�6��Ь�Ź� _�_oo(o:oLo��o�Q���_�o�o�o�o �o�o]o�o>Pb�t���o9�i�G�R<@M/�sUP_kNA�/�	i�n�v_ED�1�Y�� 
 �%-BCKEDT-��'�GETDATAU�o�9��?�j�H�o�f�\��A�^�  ���2�0&�!�E���:IB����~�ŏ׏m����3 ��&۔��D��ߟJ� ����9�ǟ�4��� ϯ�(����]�o�����5N������(��w��)�;�ѿ_��6 ϊ�gϮ�(�CϮ���ϝ�+��7��V�3� z�(��z�����i���B�8��&���~�]����F�ߟ�5����9~������]����`Y�k�����CR� !ߖ���W�q���#�5����Y��p$�NO_D�EL��rGE_U�NUSE��tIG�ALLOW 1z��(**�TEM*S	$SERV_GR��V� : REG�q$�\� NUM�
<��PMUB U�LAYNP\PMPAL�>CYC10#6� $\ULSU`�8:!�Lr~�BOXORI��CUR_��PoMCNV��10L�T4DL!I�0��	����B N/`/r/�/�/�/�/�/����pLAL_OU�T �;���qW?D_ABOR=f��q;0ITR_RT�N�7�o	;0NON�S�0�6 
HCC�FS_UTIL s#<�5CC_@�6A 2#; h� ?�?�?O#O6]CE�_OPTIOc8�qF@RIA_IIc f5Y@�2�0�F�Q�=2q&}ނA_LIM�2�.� ��P�]B���KX�P
�P�,2O�Q��B�r�qF�PQ5T1)TR�H�_:JF_PA�RAMGP 1�<g^&S�_�_�_��_�VC�  C��d�`�o!o`��`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?���2HE ONFI�� E?�aG_P�1#; ���o 1CUgy�a�KPAUS�1�yC ,���� �����	�C�-� g�Q�w���������я4���rO�A�O�H~�LLECT_�B1�IPV6�EN. QF܍3�NDE>� ��G�71234567890���sB�TR����%
 	H�/%)����� ��W���0�B���f�x� ��㯮���ү+���� �s�>�P�b������� ���ο��K��(Ϡ:ϓ�^�|��B!F�� �I|�IO #��<U%e6�'��9�K���TR�P2$���(9X�t�Y޼`�%�̓ڥH��_MO�R�3&�=��@XB��a��A� $��H�6�l�~���~S"��'�=�r_A?�a�a�`��@K��R�dP�)F�ha�- �_�'�9�%
�k���G� ��%Z�%���`�@c.�PD�B��+���cpmidbg��	�`&:�����p��N>  ��@��b.���]ܭ@as<�^��@�sg�$�f�l�q��ud�1:��:J��DE�F *ۈ��)��c�buf.t�xt����_L�64FIX , ������l/[Y/�/}/ �/�/�/�/
?�/.?@? ?d?v?U?�?�?�?�?��?�?,/>#_E -���<2ODOVOhOXzO�O6&IM��.o�=YU>���d�
�6IMC��2/���ñdU�C��20�M��QT:Uw�Cz  B��i�A���A����Au�gB3��*CG�B<�=w�i�B.���B���B��5�B�$�D�%�B���ezVC�q��C�v�D����D-lE\D�n�j��Bl9"��22o�D|������ ���jC�C����
ЙxObi�D4cdv`Dů�`/�`v`s]E��D D�` E�4�F*� Ec���FC��u[F����E��fE���fFކ3F�Y�F�P3�Z���@�33 ;��O>L���Aw�n,au@��@e�5Y��H�a���`A��w�=�`<#�*
��?�oz�JRSMOFST� (�,bIT1���D @3��
д�X'�a��;��b�w?���<��M�NTEST�1O�CR@�4��>V�C5`A�w�Ia+ah�aORI`CTPB�U�3C�`4���r��:d�*�qI?�5���qT_�PROOG ��
�%$/�ˏ�t��NUSER�  �U������K�EY_TBL  �����#a��	
��� !"#$�%&'()*+,�-./��:;<=�>?@ABC�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~��������������������������������������������������������������������������������͓���������������������������������耇��������������������������LC�K�
����STA�T/��s_AUTO/_DO �	�c��INDT_ENB�P���Rpqn�`�T2����STOr`���;XC�� 26�) �8
SONY �XC-56�"b�����@��F( �А�HR5!0w���>�P�7b�t�Aff����ֿ� Ŀ����C�U�0� yϋ�fϯ��Ϝ�����p���-ߜ�TRL��oLETEͦ ���T_SCREEN� ��kc�s���U�MME�NU 17�� <ܹ���w����� ����K�"�4�� X�j���������� ��5���k�B�T�z� �������������� .g>P�t� �����Q (:�^p��� �/��;//$/J/ �/Z/l/�/�/�/�/�/ �/�/7?? ?m?D?V? �?z?�?�?�?�?�?!O �?
OWO.O@OfO�OvO��O�O(y��REG c8�y����`�M��ߎ�_MANUAyL�k�DBCO���RIGY�9�DBG�_ERRL��9��ۉq��_�_�_ }^QNUMLI�p�ϡ�pd
�
^QP�XWORK 1:���_5oGoYoko}o�ӍDBTB_N� S;������ADB_AWA�YfS�qGCP r
�=�p�f_AL�pR��bbRY�[�
�WX]_�P 1<{y�n�,�%oc�P��h�_M��ISO��k@|L��sONTIMXכ�
���vy
���2sMOTNEN�D�1tRECOR�D 1B�� �<��sG�O�]�K� �{�b��������V�Ǐ �]����6�H�Z�� �������#�؟��� ���2���V�şz��� �����ԯC���g�� .�@�R���v�寚�	� ��п���c�χ�#� ��`�rτϖ�Ϻ�)� ��M���&�8ߧ�\� G�Uߒ�߶�����I� �����4�� �p7� n���ߤ������ ���"���F�1���|� �������[�����i� ��BTf���b�TOLERENC��dB�'r�`L���^PCSS_CCS�CB 3C>y�`IP�t}�~� <�_`r�K�� ���/�{��5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_��~�LL� D���&qET�c�a C[C��PZP^�r_ A� p� ��sp��QGPt[	 CA�p�Q�_�[? ��_�[oU�p��P�pSB�V�c��(a�PWoio{h+�o³X�o�oY���[	r�hLW��N�:p����}6ګ�wc��aD@V�B��|�G����+��Kۃ �otGhXGr��So����eB �  =��Ͷa>L�tYB�� �pC�p�q�aA"�H�S�Q-� �q���ud�v������AfP ` 0��c�D^P��p@�a
�QXTHQ����a aW>� �a9P��b�e:�L�^�h�Hc�́PQ�RFQ�PU �z�֟�o\^��-��?��c�u����zC%z�ů�b2�ЩްRD�����l)*����S̡0��]�@0�.��@���EQ�p ��F�X�ѿUҁп��VSȺNSTCY� 1E��]� ڿ��K�]�oρϓϥ� �����������#�5߀G�Y�k�}ߏߒ��D�EVICE 1F5� MZ�۶a���	� ��?�6�c���	�{䰟���_HNDGD G5�VP��|�R�LS 2H�� ���/�A�S�e�w������ ZPARAM �I�FgHe�R�BT 2K��8bр<��WPpC�C��,`¢P�Z�z��U%{�C��2��jMTLU,`"nPB, s��M� }�0gT�g��
B��!�bcy�[2Dc hz����/�x�/gT#I%D���C�` b!�R��A���A,��B_d��A��P��_cC4kP�!2�C��$|Ɓ�]�ffA�À_��B�� �| a���/�/�T (�� 54a5�}%/7/d? /M?_?q?�?�?�?�? �?O�?OO%O7OIO �OmOO�O�O�O�O�O �O�OJ_!_3_�_�_3 �_�_�_�_�_o�_(o oLo^oЁ=?k_IoS_ �o�o�o�o�o�o�o #5G�k}� ������H�� 1�~�U�g�y�ƏAo� Տ���2�D�/�h�S� ��go����ԟ����ϟ ���R�)�;���_� q����������ݯ� <��%�7�I�[�m��� ������}�&��J� 5�n�YϒϤϏ��ϣ� ѿ������F��/� Aߎ�e�w��ߛ߭��� ������B��+�x�O� a����������� ,���%�b�M���q��� ������������ L#5�Yk}� �� ��6 1CUg���� ����	//h/�� �/w/�/�/�/�/�/
? �/.?@?I/[/1/_? q?�?�?�?�?�?�?�? OO%OrOIO[O�OO �O�O�O�O�O&_�O_ \_3_E_W_�_?�_�_ �_�_�_"ooFo1ojo E?s_�_�om_�o�o�o �o�o0f=O a������� ���b�9�K���o� ��Ώ��[o��(���L�7�I���m�������$DCSS_SL�AVE L����ё~��_4D  љ���CFG M�ѕ�������FRA:\Đ�L-�%04d.C�SV��  }�� m���A i�CHq�z������|�����  �����Ρޯx̩ˡҐ-��*�����_CRC_OU/T N�������_FSI ?>њ ���� k�}�������ſ׿ � ����H�C�U�gϐ� �ϝϯ��������� � �-�?�h�c�u߇߰� �߽���������@� ;�M�_������� ��������%�7�`� [�m������������ ����83EW� {������ /XSew� ������/0/ +/=/O/x/s/�/�/�/ �/�/�/???'?P? K?]?o?�?�?�?�?�? �?�?�?(O#O5OGOpO kO}O�O�O�O�O�O _ �O__H_C_U_g_�_ �_�_�_�_�_�_�_ o o-o?ohocouo�o�o �o�o�o�o�o@ ;M_����� �����%�7�`� [�m��������Ǐ�� ����8�3�E�W��� {�����ȟß՟�� ��/�X�S�e�w��� �����������0� +�=�O�x�s������� ��Ϳ߿���'�P� K�]�oϘϓϥϷ��� ������(�#�5�G�p� k�}ߏ߸߳����� � ����H�C�U�g�� ������������ � �-�?�h�c�u����� ����������@ ;M_����� ���%7` [m����� ��/8/3/E/W/�/ {/�/�/�/�/�/�/? ??/?X?S?e?w?�? �?�?�?�?�?�?O0O +O=OOOxOsO�O�O�O��O�C�$DCS_�C_FSO ?�����A? P �O�O _?_:_L_^_�_�_�_ �_�_�_�_�_oo$o 6o_oZolo~o�o�o�o �o�o�o�o72D Vz����� ��
��.�W�R�d� v������������ �/�*�<�N�w�r��� ������̟ޟ��� &�O�J�\�n������� ��߯گ���'�"�4� F�o�j�|�������Ŀ ֿ������G�B�TϾ�OC_RPI�N _jϳ����ς��O��`��1�Z�U��NSL��@&�h߱��������� "��/�A�j�e�w�� ������������ B�=�O�a��������� ��������'9 b]o����� ���:5GY �}������ ///1/Z/U/g/y/ �/�/�/�/�/�/�/	? 2?-???Q?z?u?��� �߆?�?�?�?OO@O ;OMO_O�O�O�O�O�O �O�O�O__%_7_`_ [_m__�_�_�_�_�_ �_�_o8o3oEoWo�o {o�o�o�o�o�o�o /XSew� �������0� +�=�O�x�s������� ��͏ߏ���'�P��K�]�o����� �PR�E_CHK P�۪�A ��,�8�2��� �	 8�9�K��� +�q���a�������ݯ �ͯ�%��I�[�9� ���o���ǿ��׿�� �)�3�E��i�{�Y� �ϱϏ��������� ��-�S�1�c߉�g�y� ���߯����!�+�=� ��a�s�Q����� ���������K�]� ;�����q��������� ����#5�Ak {����� �CU3y�i ������/-/ G/c/u/S/�/�/�/ �/�/�/??�/;?M? +?q?�?a?�?�?�?�? �?�?�?%O?/Q/[OmO O�O�O�O�O�O�O�O _�O3_E_#_U_{_Y_ �_�_�_�_�_�_�_o /ooSoeoGO�o�o=o �o�o�o�o�o= -s�c��� ����'��K�]� woi���5���ɏ���� ����5�G�%�k�}� [�������ן�ǟ� ���C�U�o�A����� {���ӯ����	��-� ?��c�u�S������� Ͽ῿�����'�M� +�=σϕ�w�����m� �����%�7��[�m� K�}ߣ߁߳��߷��� �!���E�W�5�{�� �ϱ���e�������	� /��?�e�C�U����� ����������= O-s����] ����'9] oM������ �/�5/G/%/k/}/ [/�/�/��/�/�/�/ ?1??U?g?E?�?�? {?�?�?�?�?	O�?O ?OOOOuOSOeO�O�O �/�O�O�O_)__M_ __=_�_�_s_�_�_�_ �_o�_�_7oIo'omo o]o�o�o�O�o�o�o !�o1W5g� k}������ /�A��e�w�U����� ��я��o����	� O�a�?�����u���͟ �����'�9��]� o�M���������ۯ�� ǯ�#�ůG�Y�7�}� ��m���ſ�����ٿ �1��A�g�E�wϝ� {ύ�������	�߽� ?�Q�/�u߇�e߽߫� ���������)��� _�q�O�������� ������7�I���Y� �]������������� ��!3WiG� �}����%� A�1w�g� �����/+/	/ O/a/?/�/�/u/�/�/ �/�/?�/9?K?�/ o?�?_?�?�?�?�?�? �?O#OOGOYO7OiO �OmO�O�O�O�O�O_ �O1_C_%?g_y__�_ �_�_�_�_�_�_o�_ +oQo/oAo�o�owo�o �o�o�o�o);U_ _q����� ���%��I�[�9� ���o���Ǐ����� ۏ!�3�M?�i��Y� ������՟�ş�� ��A�S�1�w���g��� �������ӯ�+�=���$DCS_SG�N QK�c���7m� 09�-MAY-19 �14:33   �O�14-JA}Nt�08:38}������ N.DѤ���������h��x,rWf*�o��^M��  O��VERSION �[�V3.�5.13�EFLOGIC 1RK���  	���P�?�P�N��!�PROG_EN/B  ��6Ù��o�ULSE  �TŇ�!�_ACC�LIM�����Ö��WRSTJ�NT��c��K�E�MOx̘��� ���I?NIT S.�G��Z���OPT_SL� ?	,��
 ?	R575��YЫ74^�6_�7_�50��1��2_�@ȭ�|�<�TO  H�跿��V�DEXҚ�dc����PA�TH A[�A�\�g�y��HCP�_CLNTID y?��6� @�������IAG_G�RP 2XK� ,`� ��� �9�$�]�H������1234567890����S�� |�������!�� ��H���@;�dC�S���6 �����.� Rv�f��H ��//�</N/� "/p/�/t/�/�/V/h/ �/?&??J?\?�/l? B?�?�?�?�?�?v?O �?4OFO$OjO|OOE� �Oy��O�O_�O2_���_T_y_d_�_,
�B^ 4�_�_~_`O o�O&oLo^oI��Tjo �o.o�o�o�o�o �O '�_K6H�l� ������#�� G�2�k�V���B]��� Ǐُ�������(���L�B\Drx�@���PC����4�  79֐�$��>���:�����ߟ�ʟܟ���CT_C�ONFIG Y���Ӛ�e�gU���STBF_TTS��
��b����Û�u�O�MAU���|��MSW_CuF6�Z��  伿OCVIEW��[ɭ������-� ?�Q�c�u�G�	����� ¿Կ������.�@� R�d�v�ϚϬϾ��� ����ߕ�*�<�N�`� r߄�ߨߺ������� ��&�8�J�\�n�� ��!����������� ��4�F�X�j�|����KRC£\�e��!*� B^������C2�g{�SBL_FA?ULT ]��ި>�GPMSKk���*�TDIAG �^:�աI���UD1: 6789012345�G�BSP�-?Q cu��������//)/;/M/� �
@q��/$��TRECP��

 ��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOi/{/�xO�/UMP_OP�TIONk���AT�R¢l��	�EPM�Ej��OY_TEM�P  È�33B�J�P�AP�D�UNI��m�Q��Y�N_BRK _�ɩ�EMGDI_�STA"U�aQSUN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 J�#�{�,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;��A����O ���� � I ߵ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$
T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����裆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7����; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  D�C����(7�?�<B�?B����2�ٸ*9�N SMTT#t�[)��X}�C�f�HoOSTCd1ux����?�� M5Cx��;zOx�  27.0�@=1�O  e�O�O 	__-_;Z�O^_p_�_�_�LN_HS	ano?nymous�_�_�_oo1o yO��FhFk�O�_�o�O�o�o �o�oJ_'9K] �o�_����� 4o�XojoG�~�o^� ������ŏ���� �1�T���y����� ������,�>�@�-� t�Q�c�u��������� ϯ���(�^��M� _�q�����ܟ� �ݿ ��H�%�7�I�[Ϣ� ϑϣϵ����l�2� �!�3�E�Wߞ���¿ Կ����
������� /�v�S�e�w���� ���������+�r� �ߖ�s�����߻��� �������'9K] ��������� 4�F�X�j�l>��} ������/ /1/T��y/�/�/�/�/.D\AENT {1v
; P!J/.?  ��/3? "?W??{?>?�?b?�? �?�?�?�?O�?AOO eO(O�OLO^O�O�O�O �O_�O+_�O _a_$_ �_H_�_l_�_�_�_o �_'o�_Koooo2o{o Vo�o�o�o�o�o�o 5�oY.�R��v��zQUIC�C0���3��t1 4��"����t2��`��r�ӏ!ROUT�ERԏ��#�!�PCJOG$����!192.16?8.0.10��s?CAMPRTt�P��!d�1m�����R�T폟�����$NA�ME !�*!�ROBO���S_�CFG 1u�)� �Au�to-start{edFTP&��=?/֯s��� �0�B��f�x����� ����S������,� ��������ϼ�ޯ�� �������ʿ'�9�K� ]�oߒ�ߥ߷����� ����(:~�k� �Ϗ���������� ��1�C�f���y��� ���������,�>� R�?��cu��`� ����(�$ M_q������  /H%/7/I/[/ m/4�/�/�/�/�/� ~/?!?3?E?W?i?� ���?�/�?/�?O O/O�/�?eOwO�O�O �?�ORO�O�O__+_ r?�?�?�?�O|_�?�_ �_�_�_o�O'o9oKo ]ooo�_o�o�o�o�o �o�oF_X_j_~ok �_������o� ��1�TU��y����������U�)�_ER�R w3�я�P�DUSIZ  jg�^�p���>�?WRD ?r�Cq��  guestb�Q�c�u��������"�SCDMNGRP 2xr�w���Cq�g�\�b�K� 	�P01.00 8~(q   �5p��5pz�5pB � �{ ����H���L���L��L�����O�8�����l�����a�4� x��Ȥ�x��V8���\���)�5`�;��������d�.�@�R�ɛ_�GROUېy������	ӑ���Q?UPD  ?u��Y��İTYg�����TTP_AU�TH 1z�� �<!iPend�an��-�l����!KAREL:q*-�6�H�KC]��m��U�VISI?ON SET���� ��g�G�U������R� 0��H�Bߏ�f�x�����߮���CTRL C{����g�
S��FFF9E3���AtFRS:D�EFAULT;��FANUC W�eb Server;�)����9�K��܀����������߄W�R_CONFIGw |ߛ ;���IDL_CPU�_PCZ�g�B��Dpy� BH_�MI�Nj�)�}�GNR_�IO��g���a�N�PT_SIM_D�_�����STAL�_SCRN�� ����TPMODNT�OL������RTY`��y���� �ENO����Ѳ]�OLNK 1}��M���������eMA�STE��ɾeSL?AVE ~��c>�O_CFGٱ�BUO�O@CY�CLEn>T�_A�SG 1ߗ+�
 ����// +/=/O/a/s/�/�/�/��/��NUM�z�
@IPCH��^RTRY_CN Z���@��������� @kI��+E�z?E�a�P_M�EMBERS 2Y�ߙ� $���2����ݰ7�?�9a�S�DT_ISOLC�  ����$J_23_DSM+��3JOBPROC�N��JOG��1��+�d8G�?��+�O�/?
�LQ�O__/_�O S_e_w_�_`�O H�m@��E#?&BPOS�REQO��KANJ�I_���a[�MON ����b�yN_goyo�o�o�o�$Y�`3�<� ��e�_ִ��_L���"?`�EYLOGGIN�LE��������$LANGUAGgE ��<T�Y {q�LGa2�	��b���g�xP�� � ��g�'Զ�b���>�M�C:\RSCH\�00\<�XpN_D?ISP �+G�pJ��O�O߃LOC�p�Dz���AsO�GBOOK �������󑧱����X�����Ϗ���`�a�*��	p� ����!�m��!���=p�_BUFF 1�p��2F幟����՟D� Col�laborativǖ���F�=�O�a� s�������֯ͯ߯����B�9�K���DC�S �z� =���'�f��?ɿۿ����H@{�IO 1��� ~?9ü�� 9�I�[�mρϑϣϵ� ���������!�3�E� Y�i�{ߍߡ߱����ߴ���E��TMNd �_B�T�f�x���� ����������,�>� P�b�t�������L��SEVD0��TYPN1�$6���QRS"0&��<2�FL 1�"�J0���������GTP:pO>F�NGNAM1D��mr�tUPS�GI�"5�aO5�_LO{ADN@G %��%TI�pZUZ�AUN#�(MAXUALRM�'���(���_PR"4F0�d��1�B_PNP�� V 2�C	�MDR0771�ߕ�BL"806=3%�@ �_#?�hߒ|/�C��z��6��/���/Po@P �2��+ �ɖ	�T 	t  ��/�%W?B?{?� k?�?g?�?�?�?O�? *OONO`OCO�OoO�O �O�O�O�O_�O&_8_ _\_G_�_�_u_�_�_ �_�_�_o�_4ooXo joMo�oyo�o�o�o�o �o�o0B%fQ �u������ ��>�)�b�M����� {��������Տ�� :�%�^�p�S��������D_LDXDI�SApB�MEM�O_APjE ?=C
 �,� (�:�L�^�p�������� 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%� �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A�z�4��~�K��������K:z�j]�Q_D��^��PL_NAME �!3%,�!�Default �Personal�ity (fro�m FD) �R�R2� 1�L?6(L?�,0	l d���� ����//(/:/ L/^/p/�/�/�/�/�/�/�/ZX2u?0?B? T?f?x?�?�?�?�?\R<?�?�?O O2ODO�VOhOzO�O�O�OZZK`\R�?�N
�O_\TP�O:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHo_)_~o�o �o�o�o�o�o�o  2DVhz�[omo ����
��.�@� R�d�v���������Џ�� Ef  Fb� F7���   ��!��d��@�R�6�t��� ���l���ʝ����� ݘ���� "�@�F�d���� "�|��ݐA�  ϩ�U[�$n�B��E ��� � @D�  &�?�� �?�@��A@�;f��FH�� ;�	l,�	 '|��j�s�d�/>��� ��� �K(��Kd$2�K ��J7w��KYJ˷�ϜJ�	�ܿ�� @�I���_f�@w�z��f򿿾γ�N�������	Xl�����_��S�ĽÔ�}�I ����5�?��  ����A�?oi#�;����� ���l� �Ϫ�-���ܛ�G�G�Ѳ��@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=�����в@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj��a�Be�Ci��#��Bи�ee^��^^ȹBР ��P����̠�����ADz՟�n�3��C��i�@�R�R�Y���� { �@� ����  ���?�ff0������n� ɠ #ѱy9G
(���I�	(�@uP~����t��t���>����;�C�d;��.<���<�g�<F+<L�������,��d�,�̠?fff�?��?&&��@���@x��@��N�@���@T�H�ِ�!-�ȹ �|��
`���� ���//</'/`/`r/]/�/��eF�� �/�/�/�/m?��/tJ?�(E��G�#�� FY�T?�?P? �?�?�?�?�?O�?/O O?OeOk��O�IQO G�?�O1?�OmO_0_�B_T_������A _�_	_�_�_�_ o���A��An0 bФ/o �C�_Uo�_�Op���؃o�o�o�o���W������oC�E�� q�H�d�����a@q��e�F�Bµ�WB]�NB2��(A��@�u�\?�D��������b�0�|�u�R����
x~��ؽ��B�u*C��$�)�`�$ ����GC#����rAU�����1�eG�D�I��mH�� I:��I�6[F�﫹C�I���J�:\IT��H
~QF�y���p�*J��/ I8Y�I��KFjʻCe �o��s�����Џ��� ߏ�*��N�9�r�]� �����������۟� ��8�#�\�G�����}� ����گů���"�� �X�C�|�g�����Ŀ �������	�B�-� f�Qϊ�uχ��ϫ��� �����,��P�b�M� ��qߪߕ��߹����� ��(��L�7�p�[��@�������s($�ϳ�3:����$���3���d�,��4��@�R�wa�ǲ��l�~�wa����e����wa4 �{������(L�:ueP�P~�A �O������	����G2 W}h����� �/���O�O7/m/[(d=�s/U/�/�/�/ �/�/?�/1??U?C?�y?�=  2 E�f9gFb��77�b9fB)aa)`C9A`	�&`w`@-o�?w`e�@O)O�?MO�Ow`�?@�?�O�O�O�O9c?�0T�A7ht4w`w`�!w`xn
  �O9_K_]_o_�_�_�_ �_�_�_�_�_o#ozz�Q ��h��G����$MR_CA�BLE 2�hO �a�T� @@�0�Ae��a�a��a��`��0�`C��`�aO8�tB�^n�d��`�aE�4�E�#��o�f�#��0�|�0�DO��By`���Š��bED4E�c,��o�g8  ���Cu�07�d4
v�ے�0 �b���XE�Z&�lȠ`y`
qC�p�bHE݈
v#g�5DͣҮ�qz�lҠ`�p�0�q�p�b0�
v׸%c���b=%	E;h��u/o�c -��4tH�\�?�9�K� ]�o�ԏϏ��
�ɏۏ�@���?��eo �a���������b����� �����`�	 ���������`�� ���퐺@�����ŀ�U�ݐ����������������*,� ,�-�\c�OM �ii���3� �V ���%% 23�45678901�i�{� f��������ԋ��1����
���`�not �sent3������;�TEST�FECSALGRG  e�qiG�1d.�Zš
:�� �D�CbS�Q�c�u��� 9�UD1:\ma�intenanc?es.xml��ֿ�q� =���DEFAULT�-�i4\bGRP 2�M�  =��a����   �%Force��sor chec�k  ���b�z��p����h5-[ �ϻ��������dID�%!1�st clean�ing of c�ont. v�i?lation��}�Rߗ+��[�ߔߦ������mech��cal`����B��0��h5k߀@�R�d�v�����(�rolle_Ƶ�����/���(�:�����Basic �quarterl!y�������,����`������M��M��:C@"GpP�a�b`i4��������#C���M"���{Pbt����Suppq�gre�ase����?/&/8/J/\/��C�+ ge��. ba�tn�y`/��/h5	 /�/�/�/? ?_���en'�v��/�/��/��?�?�?�?�?F�G=?O�qp"CrB1O��0�/`OrO��O�O�O�t$��Lf���C-m��A�O:��OO$_6_H_Z_l_��t*cabl�Om����S<m��Q�_:�
 _�_�_oo0oo)(��/�_�_���_�o�o��o�o�o�O@h�au1�l�2r !xm�<qC:��op�������ReplaW�fUȼ2�:�._4�F�X�j�|�m�$%���o������� #���
��.�@���d� ��ŏ׏����П��� �U�*�y�����r��� ������	�q��?�߯ c�8�J�\�n���ϯ�� ���ڿ)����"�4� Fϕ�jϹ�˿����� �������[�0�ϑ� fߵϊߜ߮�����!� ��E�W�,�{�P�b�t� ����߼�����A� �(�:�L�^������ �������� $ s�H������q�� ���9]o� Vhz���U� #�G/./@/R/d/ ��/�/��//�/�/ ??*?y/N?�/�/�? �/�?�?�?�?�???O c?u?JO�?nO�O�O�O8�O+J�r	 H�O�O __6M2_@OBE:_p_ >_P_�_�_�_�_�_ o �_�_oHoo(oZo�o ^opo�o�o�o�o�o ��o :z �bA?�  @�q  _���Fw��� �H* �** @q>v�p2T�f�x��:�������ҏ�� eO^C7�Տ#�5�G�	� k�}���ُ���c�� ���W��C�U�g��� ß)�����ӯ���	� �-�w�����9����� ��m�Ͽ��=�O�E�	A�$MR_H�IST 2�>u�N�� 
 \�$Forc�e sensor� check  �12345678�90q�3�������N}SB�� -319.8� hours R�UN 9.�Y�!�1st clea�ning of �cont. ve�ntilatio�n0ÄϖϨ�-�� $��mech���cali�%Ό4���o�DN�t&��95��1����rolleh�+�=��O���Bas�ic quarterlyߒߤ߶� 
O4�F��(���� ��b�t���������� �M�_����:������p���:�SKCFM�AP  >u�Q��r5��������ONREL  .�3���?EXCFEN��:q
��QFNCX�JJOGOVLI�M8dNá ��KE�Y8��_PAN7����������SFSP�DTYPxC��S�IG�:��T1M�OT�G��_C�E_GRP 1�>u\�D�� ���/Ⱥ��/ �/U//y/0/n/�/ f/�/�/�/	?�/??? �/c??\?�?P?�?�? �?�?�?O)OOMO,����QZ_EDIT�5 )TCOM_�CFG 1����[�O�O�O 
�ASOI �y3�
__+[_O_���>O�_bHT_AR�C_UքT_MN_MODE5��	UAP_C�PL�_gNOCH�ECK ?�� �� o.o@o Rodovo�o�o�o�o�o��o�o*!NO_WAIT_L4l~GiNT�A���|EUwT_ERRs2���3��ƱJ������>_)��|MO�s��}x:Ov���?8�?������ l��rPARAuM�r������j���5�5�G� =  r�b�t�s�X��� ���������֟�0����b�t������SUM_RSPA�CE�����Aѯۤ�$ODRDSP�S�7cOFFSET�_CARt@�_�D�IS��PEN_FILE:�7�AF��PTION_I�O��q�M_PR�G %��%$*�����M�WORK ��yf �!�춍�����r����	 �������gT��RG_DSBL  ���C�{u��RIE�NTTO7 ��Cٴ A �UT�_SIM_Dy����V�LCT ��}{B �٭�ď_PEX�P=��R[AT�W dc�>�UP ���`���e�w�]ߛߩ���$�2r�L�6(L?���	l d������ &�8�J�\�n���� �����������"�4�F�X���2�߈����� ��������*�<w�Tfx��������J`�ˣG���Tz�Pg���� ��/"/4/F/X/j/ |/�/�/�/���/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?�/�/ ,O>OPObOtO�O�O�O �O�O�O�O__(_:_��O��y_�]2����_�^�_�_�W^]@^]��/ooSog� Hgrohozo�o�o�o�o��oF`�#|`�AG�  9y����OK��1�k�����<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	 '|�Q�s�r�q/>��u �sF`�H<zH~��H3k7GL�z�HpG�9�9l7�k_B�T�F`C4T��k�H���t��-��Ae���k������s���  ��ሏ����EeBVT����dZ��g���ڏ ����q-�Fk�y�{FbZU���n@6�_  ���z��Fo��Be	'� �� ��I� ��  �:p܋=����ڟ웆�@���B�,���B��g�AgN���� � '|���g��B�*��p�BӀC׏�����@  #�B�u�&�ee�^^މB:p2����>�m�6p�Z���Dz ?o}�܏������׿�������Ǒ��� f� � � �M���*�?�ff�_8�Jφܿ 3pϑ�ñ8@�Чϵʖq.·�(����P���'��s�tL��>��/�;�Cd;���.<߈<��g�<F+<AL ��^oiΚrd@�|�r6p?fff?��?&�п�@���@x��@�N��@���@T� ��Z���ћtމ�u�� �w	�x��ti�>�)�b� M��q��������� ����:�%�^��������W���S�E�  �G�aF�� Fk���������1 U@yd���� ��q��	��{�A ��h�����a��ird��A{/w�/J/5/n/vA��A0���":t�/ C^/�/xZ/ ލ?���/��/1??���W���t�g��pE� ~1��?04�0
1�1@�IӀ��BµW�B]�NB2�(�A��@�u\�?����������b�0�|�uR�����
�>��ؽ��Bu�*C��$�)`��? ���G�C#���r�AU����1��eG���I�m�H�� I:��I�6[F����C4OI���J�:\IT��H
~QF�y��Ol@�*J�/� I8Y�I��?KFjʻC��-? �O�O__>_)_b_M_ �_�_�_�_�_�_�_o �_(oo%o^oIo�omo �o�o�o�o�o �o$ H3lW�{� ������2�� V�h�S���w�����ԏ �������.��R�=� v�a�������П���� ߟ��<�'�`�K�]� ��������ޯɯ��&�8�#�\��3(J��g�3:a������J�3��c4�������������1��㚅ڿ��1����e���14 �{ 2�2�r�`ϖτϺϨ�J�%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ��� �������3��W�B� {�f�4���������d�A����!��1�3� E�{�i��������������  2 Efn�7Fb�7��6�B�!�!� C9� �� �0@�/`r������#x��+=�3?, V�8�v��0�0�:�0�.
 D� ����//%/7/�I/[/m//�/�:� ���ֻ�G����$PARAM_M�ENU ?2���  �DEFPUL�SE�+	WAI�TTMOUT�+�RCV? S�HELL_WRK�.$CUR_ST�YL� 4<OP9TJJ?PTB_?Y2�C/?R_DECSN 0�Ű<�?�?�?�? �?OO?O:OLO^O�O��O�O�O�O�!SSR�EL_ID  �.�����EUSE_PROG %�*q%�O0_�CCCR0��B���#CW_HOSoT !�*!HT�_=ZT��O_�Sh_zQ��S�_<[_TIM�E
2�FXU� GD�EBUG�@�+�CG�INP_FLMS�Ko5iTRDo5gP+GAb` %l�tk�CHCo4hTYPE
�,� �O�O�o# 0Bkfx�� �������C� >�P�b���������ӏ Ώ�����(�:�c��^�p�����7eWOR�D ?	�+
 �	RSc`��P�NS��C4�JO�v1��TE�P��COL�է�2��gLVP 3�����Oj�TRACECTL� 1�2��!{ �� ��Қ�q�DT Q�2�Ǡ��D �� :��f��Ԡ�Ԡ���}�ׯ���;�4��4��4� ��;�u:�q:���;�U8�	8�
8�8�U8�8�8�8�T�@:�8�8����� ���ٱ޴���ؿ�$�6��� 
�l�~�@�R�dϞϰ� ��������
��V�h� zߌߞ߰��������� 
�,�>�P�*�<�v���*� +8� (
��)��*�������� ��)�;�M�_�q��� ������������ %,�>�P�b�t����� �������С�* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6@u bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� V�߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�?��?�1�$PGTR�ACELEN  ��1  ����0��6_U�P ����2A@�1@�1_CFG �ES�3�1
@�<D�0<DZO<C�0uO�$BDEFSPD ��/L�1�0���0H_CONFI�G �E�3 U�0�0d�D��2 �1�APpDsA�A��0��0IN'@T�RL �/MOA8lpEQPE�E��G��A<D�AIL�ID(C�/M	bTG�RP 1ýI �l�1B  ������1A�3�3FC� F8п E�� @eN	��A�AsA�Y�Y�A�@� 	 vO�Fg��_ ´8cokB ;`baBo,o>oxobo�o��1>о�?B�/�o�o~�o =?%<��
C @yd��"�������  Dz@�I�@A0�q� ��� ����ˏ���ڏ��� 7�"�4�m�X���|����Ú)ґ
V7.10beta1HF @�����Aq��Q m �?� �BܠPz�p �C��&�?B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@��8�f������ҡ�R9�ܣ�Rљ���1��i�������t<B!CeQKNOW_M  lE7FbT�SV ĽJ �BoC_�b�t�������@������1�]aSM�S]ŽK ���	NB~�0���Ŀ�K���-�bb ��A�RP����0��Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1�K
 4MU�iǨj� K�]�oߠߓ� �߷�������2��#� h�G�Y��}�����@��
������,�27�9I��1�<t�H���P3^�p�����,�4 ��������,�5(:,�6Wi{��,�7����,�8��!3,�MAD��6 F,�OVL/D  KD�xO�.�PARNUM � �MC/%�SCH� E
9'!G)�3Y%UPD/��E|�/P�_CMP_���0@�0'7E�$E_R_CHK�%5H�&�/�+RS���bQG_MO�+?=5_'?~O�_RES_G6��:�I�o�?�?�?�? O�?O7O*O[ONOO�rO�O�O�{4]��< �?�Oz5���O__|3  #_B_G_|3V b_�_ �_|3� �_�_�_|3�  �_�_o|3Oo>oCo|2V 1�:�k1!��@c?�=2THR_INRc0i!}�zo5d�fMASS�o� Z�gMN�o�cM�ON_QUEUE� �:�"�j0��*O�N� U1Nv�+�DpENDFqd?`yEcXEo`u� BEnp|PAsOPTIOMw�m;DpPROGRAoM %$z%Cp�}o(/BrTASK_�I��~OCFG ��$��K�DAkTA��T���j12/ď֏���� ��+�=�O�a������𩟻�͟��INFO
�͘��3t��!�3� E�W�i�{�������ï կ�����/�A�S��e�w�����Θ� �'��FJ�a K_N�q�T��˶ENBg Hڽw1��2��GN��2�ڻ P(�O�=���]ϸ��@���v� ��u�uɡdƷ_EDIT �T�����>G�WERFL�x�c�)�RGADJ �Ҷ�A�  $�?@j00��a�Dqձӆ5�?�����<u�)%e���Ș��FӨ�2�R��	�H;pl�G�b_�>��pAod�t$��*�/� **�:�j0�$�@�5 Y�T���^��q�߈b ~�L��\�n���� �����������4� F�t�j�|��������� ����bLBT �x����:� �$,�Pb� ��/����/ ~/(/:/h/^/p/�/�/ �/�/�/�/V? ??@? 6?H?�?l?~?�?�?�? .O�?�?OO O�ODO VO�OzO�O_�O�O�O �O�Or__._\_R_d_��_�_�_�_�_�_�f	 g�io�pWo�o{d�o��~o�ozoB�P?REF �Rږp��p
�IORI�TY�w[���MP�DSP�q��pwUT�6����ODUCT�3�����OG��_TG��8�����rTOENT 1�׶� (!AF_INE�p,�7�?!tcp7�_��!udN���!icmv��ޯrkXYK�ض���q�)� ,�����p��&�	��R�9�v� ]�o�����П����� �*��N�`�*�sK���9}�ߢ���Ư �,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE� �R��:�wd��连�2s�9Ks���PORT_NUUM�s�p����_CARTREP�{p�Ω�SKSTAv�w d�LGS)��ݶ��tӁpU�nothing��������{��TEMP ޾y��'e���_a_seiban�o\��olߒ� }߶ߡ���������"� ��X�C�|�g��� ����������	�B� -�f�Q���u������� ������,<b M�q��������(L�VE�RSIyp�w} �disabl�edWSAVE �߾z	260_0H768S?��!ؿ����/ !	5(�r)og+^/yÁe{/�/�/�/�/�*��,/? �p���_��p 1�Ћ�? �����Wh?xz?�W*pURGE��aB�p}vgu,�WF�0#DO�vƲ�vW%��4�(�C�WRUP_DELAY �\���5R_HOT �%Nf�q׿GO�5R_?NORMAL&H�rx6O�OZGSEMIjO��O�O(qQSKIPF3��W3x=_9 8_J_\_]�_�_{_�_ �_�_�_�_�_	o/oAo Soowoeo�o�o�o�o �o�o�o+=a Oq������ ��'��7�]�K���x����)E�$RA{����K/�zĀÁ_�PARAM�A3���K @.�@`\�61�2C<��y�M�C�6$�BÀ�BTIF�4`�RC_VTMOUu�cŻ�ÀDCRF3��I �+Q;�/�CC�SeD��#�1=h��-0�t]�/��ޅ�����1��0��_��k_����Cd;��.<�߈<�g�<?F+<L���Ѱ��d�u�L������� ϯ����)�;�M��_���RDIO_T?YPE  M=U��k�EFPOS1 ;1�\�
 x4/�����+�$/<�� $υ�pϩ�D���h��� ���'������o�
� ��.ߤ�Rߌ������ ��5���Y���i��*� <�v���r������� ��U�@�y����8��� \�����������?��xc����2 1�KԿX�T�x��3 1�����nY�S4 1�'9K�/�|'/�S5 1����/�/�/�/:/S6 1�Q/c/u/�/�-??Q?�/S7 1��/�/
?D?�?�?�?>d?S8 1�{?�?��?�?WOBO{O�?SM?ASK 1L�8�O�D�GXNO���Fx&�^��MOTEZ�hŻ��Q_ǁ�%]�pA݂��PL_RA�NG!Q]�_QOWE/R �ŵ�P1V�SM_DRYPR/G %ź%"O�_��UTART ���^�ZUME_PR�O�_�_4o��_EX�EC_ENB  yJ�e�GSPD`pO`WhՅjbTDBro�jRM�o�hING�VERSION �Ź#o�)I_AIRPURhP� �O(�MMT_ҡ@T�P#_ÀOB�OT_ISOLC��NTV@A'qhuN�AME�l��o�JO�B_ORD_NU�M ?�X#q�H768  �j1Zc@�r
��rV�s���r�?�r?��r�pÀPC_TI�MEu�a�xÀS2�32>R1�� �LTEACH PENDANw��:GX�!O �Maintena�nce Cons�j2����"��?No UseB�׏ ������1�C�y�V��NPO�P@�YQ��cS�CH_Lf`�%^ �	ő~��!UD1:�z��R�@VAIL�q�@�Ӏ�J�QSPA�CE1 2�ż ��YRs�i�@Ct��YRԀ'{��8�?��˯���� "���7�2�c�u����� G���߯ѿ򿵿�(� �u�AC�c�u����� Ͻ�߿���ϵ��(� �=�_�qσϕ�C߹� �����߱��$��9� [�m�ߑߣ�Q����� �߭��� ���	�W�i� {���M�������5� ��.S�e�w��� ��I������� *?as��E �����/&// ;/]o����� �/2/�/?"?�/7?Y/ k/}/�/�/O?�/�/�?��?�?O0OOKA�o�*SYPpM*��8.30261 �yB5/21/2018 A �WP�fG|�H�_TX`�� !$COMM�E�$US�Ap $EN�ABLEDԀ$sINN`QpIOR�B��@RY�E_SIG�N_�`�AP�AIT\�C�BWRK�BD<��_TYP�CRIN�DXS�@W�@%VF{RI{�_GRPԀ$UFRAM�r�SRTOOL\VMY�HOL�A$LE�NGTH_VTE�BTIRST�T ? $SECLP�X�UFINV_PO�S�@$MAR�GI�A$WAI�T�`�ZX2�\�VG-2�GG1�AI�@�S��Q	g�`_WR�BNO_USE_DI�B^uQ_REQ�BC�C�]S$CUR_T�CQP�R"a^f �G�P_STATUS>�A @ �A3`X�BLk�H$zc1�h��P@���@_�F�X �@E_MLoT_CT�CH_�J6�`CO�@OL�E�C�GQQ$W�@w��b#tDEADLO�CKuDELAY_CNT�a3qGt�a�$wf 2 �R1[1$X<�2*[2�{3[3$Zwy �q%Y�y�q%V�@�c�@��b$V�`�RV�UV�3oh>b�@ � q�d�0arMSKJ��LgWaZ�C`NRK�P�S_RATE�0�$���S
`�Q�TAC���PRD���e�S�*��a4�b  �DG��A 0�P�flp3 bquS2ppI��#`
`�P 
�S�\`  �A�Ro_ENBQ ��$RUNNER�_AXI�<`ALPLx�Q�RU�THICQ?$FLIP7��D?TFEREN��R��IF_CHSU�I0W��%V)�G1�����$PřA�Q�Pݖ_�JF�PR_P�	��RV_DATA~�A  $��ETIM���$V�ALU$�	�OP_   ��A  2 ��SC*�	� ?�$ITP_!�SQ�]PNPOU}�o�TO�TL�o�DSP��J�OGLIb��PE_IPKpc�Of�i��P�X]PTAS�$KEPT_MIR��d¤"`M�b�APq�aE�@�y�q�g@١�c�q�PG�BRK�6�x���L�I�� � ?�SJ�q�P�ADyEz�ܠBSOCz��MOTNv�DUM�MY16Ӂ$S}V�`DE_OP���SFSPD_OViR
���@LD�����OR��TP8�L�E��F������OV���SF��F����bF��d�ƣ&c)�fQc�L�CHDLY��REGCOV���`��W�P1M��gŢ�RO����r��_F�?� @v�=S �NVER�@�`�OFS�PC,�CSWDٱc�ձ���B�����TRG�š�`E_�FDO��MB_CiM}���B��BLQ��¢	�Q�̄Vza�BU�P�g��G
��A�M���@`KՊ�e�_M!�d�AMf�Q��OT$CA����DF���HBKd�v���+IOU��I'R��PA����������p���і�DVC_DB �S!�x�Q�!�s�d�9�1A��9�3A��ATIO�0��͠��aUS����WaAB�� R+c�`tá`DؾA���_AUXw�SUB'CPUP���S�`�����3Եжc���3�F�LA�B�HW_C wp"�Ns&�]sAa���$UNITS�|M�F�ATTRIz��Z�CYCL�CN�ECA���FLT�R_2_FI��TARTUPJp��ь�A��LP������_�SCT*cF_F�F1_P���b�FS��+�K�CHA/Q��*�d�RSD��Q��ص�Q���_TH�PRqOr���հEMPJ�䢠G�T� ��Q�DI�@y�R�AILAC/�bM�X�LOf�xS��ځ`���拁���PR#�S`app�C� �	��FUNC���RIN`QQP�� ԱRA)]R ���AƠ��AWAR֓��BLZaWraAkg�ngDAQ�0B�rkLD�र�&q�M�K���TaI���j��$�@�RIA_SW��AF��Pñ#��%%p�p9r1��MOIQ����DF_~P(�PD�"LM-�FA�PHwRDY�DORG��H; _QP�s%MU�LSE~Pz���*��� J��Jײ��F�AN_ALMLV�G��!WRN�%HA#RDP��UcO�� �K2$SHADO�W]�kp�a02��� S�TOf�+�_^�w�A�U{`R��eP_SBR�z5���:F��| �3MPINF?��\�4��3REGLV/1DG�+cVm L�C�CFL(��?��DAiP���Z`�� q�����Z�	 �Pv(Q$�A$Z�Q� V�@�[�
� ��EG߀o���kA#AR���㌵2�axGܘ�AXE��RO]B��RED��W�Q2D�_�Mh�SYA��AtF��FS�GWRI�P~F&�STR����E��˰EH�)��D�a�\2kPB6P��=V��D.v�OTO�1)���ARYL�tR�v�3�淡FI&�ͣ$LGINKb!\��Q��_3S���E��QX�YZ2�Z5�VOFIF���R�R�XxP	B��ds�G�cFI�03g�������_J��'�ɲ �S&qR0LTV[6���a#TBja�"�bC����DU�F7�TU�R� X��e�Q�2XP�ЊgFL�E���x@�`�U9Z8���� W1	)�K��Mw���F9��劂����OCRQj��G;W3�� �#�Ґd ���uz�����1�tOVE�q_�M ��ё?C�uEC�uKB�v '0�x-�wH��t� ��& `��qڠ�B�ё �u�q�wh�ECh����SER��K	�EPH����AT�K�6e�9e�W���AX s�'��v�/�R �� ��!�� ��P��`���`�3p�Yp�1 �p�� �� �� (� � 8�� H�� X�� h��� x�� ������DEBU�$%3�I��·RAB���ٱr�sV��� 
d� J、��@񘧕���� ���Q���a���a��3q���Yq+$�`%"<�cL�AB0b�u�'�G�RO���b<��B_s��"Tҳ*`�0A��u��uq�p1}�AND Gp�������U��p1�� �ѷ0�Qθuݸ���PNT0���SE�RVE �Z@ $�`EAV�!�PO����nP!�P@��$!Y@  ]$>�TRQ�b
=�d�BG�K�%"2\���� _  l8��5�D6ERRVb(��I��V0`;���TO	Q:�7�L�@
�R��Je G�%�Q�� <�50F� ,�`�z��>�RA� 2' d!�����S�  M��pxU �����OCuG� � ��COUNT�6Q��FZN_CFGF� 4#��6��TG4�_�=�����ü��VC ���M  �"��$6��q ��CFA E� &��X�@@�������A���r�AP��P@HEL�0~�� 5b`�B_BAS��RS)R�6�CSH��R��1�Ǌ�2��3��U4��5��6��7��98��}�ROO���̚P�PNLEA�cAB�)ë ��ACKu�IeNO�T��(B$UR08� =�_PU��!0��OU+�Pd�8j���� V��TPFWD_KAR��� ��RE(ĉ P�P�>7QUE�:RO�p�`r0P1I� x�j�Pp�f��6�QSEM���0��� A��STYfL�SO j�DIX��&�����S!_TM>CMANRQ��P�ENDIt$KEYSWITCH��ذ�kHE�`BE�ATM83PE{@L�E��>]��U��F���SpDO_H�OM# O�@�EF�pPRaB�A#PY��C� O�!���OV�_M|b<0 IOCqM�dFQ��h�;HKYA D�Q�7��UF2��M���p޸cFORC�3WA�R�"�OM|@ G @S�#o0U)SUP�@1�2&3&Q4E���T�O��L�y��8UNLOv��D4K$EDU1  ��SY�HDDN�F� M�BLO�B  p�SN�PX_AS�� �0@�0��81$S{IZ�1$VA{�~��MULTIP-���# A� � $��� /4`��BS��0�C���&F'RIFBO�S����3� NF�ODB�UP߰�%@3;9(������Z@ x��S�I��TEs�r�cSKGL�1T�Rp&���3B��@�0STMTdq�3Pg@VBW�p��4SHOW�5@��SV��_G�� 3p$PCJ�PИ���kFB�PHSP 1AW�EP@VD�0WC�� ���A00��PB XG XG �XG$ XG5VI6VI7�VI8VI9VIAVIB�VI�XG�YF�0XGFPVH��XbI1oI1|IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1Y1YU2UI2bI2oI2|I2�I2�I�`�X�I2pT�X�I2�I2�I2�I2�I2Y2Y�p�h�bI3oI3|I3�I3��I3�I3�I3�I3��I3�I3�I3�I3��I3Y3Y4�i4�bI4oI4|I4�I4��I4�I4�I4�I4��I4�I4�I4�I4��I4Y4Y5�i5�bI5oI5|I5�I5��I5�I5�I5�I5��I5�I5�I5�I5��I5Y5Y6�i6�bI6oI6|I6�I6��I6�I6�I6�I6��I6�I6�I6�I6��I6Y6Y7�i7�bI7oI7|I7�I7��I7�I7�I7�I7��I7�I7�I7�I7��I7Y7T́V5P� UD�y"ՠ���
<A62��:t�R��CMD� ���M5�Rv�]��Q_h�R���e����<��YSL���  � �%\2��+4�'�W�BVALU���b��'���FH�IgD_L���HI��9I���LE_���f��$0C�SACѿ! h �V?E_BLCK���|�1%�D_CPU5� � 5ɛ �����C�� ���R " � �PWj��#0��LA�1SBћì���RUN_FLG�� �����ĳ ��������B��H���ХĽ��TBC2��# � @ B��e �S�p8=�FTDC�����V���3d�Q�T!HF�����R�L�?ESERVE9��F��3�2�E��Н��X -$��LE�N9��F��f�RA���W"G�W_5�b�14��д2�MO-�T%	S60U�Ik�0�ܱF����[�DEk�21LgACEi0�CCS#0�� _MA� j��z��TCV����z�T�������.Bi�'AH�z�'AJh�#EM5�"��J��@@i�V�z���2Q �0&@o�h�6��JK��VK9��0{���щ�J0�����JJ��JJ��AAAL���������4��5�ӕ N1����딨�.�LD�_�1�* �CF�"% `�GROU���1��AN4�C�#m RE�QUIR��EBqU�#��6�$Tk�2$���zя #��& \�APPR� C� 0�
$OP{EN�CLOS"�St��	i�
��&' �MfЩ����W"-_MG�7C�B@�A���BBR=K@NOLD@�0RTMO_5ӆp1J��P�������������60��1�@ m1�>#�(� ������'��+#PATH''@!6#@!�<#� r� '��1SCA�؆�6IN��UChJ�[1� C0@UM�(Y ��#�"�����*����*��� PAYLO�A~J2LؠR_AN^�3L��91��)1AR_F2L3SHg2B4LO4�!�F7�#T7�#ACRL�_�%�0�'�$��H���.�$HA�2FWLEX��J!�) P�2�D߽߫����0��* : ����z�FG]D����z���%�F1]A�E�G�4�F�X�j�|���BE ������������ (��X�T*�A���@�X I�[�m�\At�T$g�QX<�=��2TX���e mX��������������@����+	�J>+ �-�K]o|��٠AT�F�4�ELPFPѪs�J� *� ;JEmCTR�!�A�TN�vzHAN/D_VB.��1��n$, $8`F2Av���SW�
"-� $$M*0 .�]W�lg��PZ����A��� 1�����:AK��]AkA�z��LN�]DkD�zPZ G��C�ST�_K�lK�N}DY ��� A����0��<7 ]A<7W1�'��d�@g`�P��������"
"J"�. �M�2D%"��H����A'SYMj%0�� j&!-��-W1�/_�{8 � �$�����/�/�/�/ 3J<�:9�/�\89�D_VI�v�|���V_UNI�����cD1J����╴� W<��n5Ŵ�w=4��9 ��?�?<�uc�4�3ɴ�%�H���/0�j��0�DIzu�O�İ�k�>0) �`��I��A��# ���@ģ���@��IP�l� 1 � /�ME.Qp��9�ơT}�PT�;pG �+ Gt� ���'���T�0 $�DUMMY1��o$PS_�@RF�@�;�$b�'FL�A@ YP(c|��?$GLB_TP�ŀ����9 P�q��2c X� z!ST9��� SBRM M2�1_V�T$SV_ER*0O�p����SCL����AGPO�¶f�GL~�EW>�3s 4H �$Yr�ZrW@�x�A1+�A����";�"�U&�4 �8`NZ�"�$G�I�p}$&� p-� �Y�>�5 LH \{��}$F�E��NEAR(PN�CF<��%PTANC�B;��JOG�@� 6�9�$JOINTxwa?pd�MSET>�7  x�E��HQtp�S{r��up>�8�k �pU.Q?�� LOCK_FOV0�6���BGLV�sG�Lt�TEST_X9M� 3�EMP��q���_�$U&@�%�w`24� Y��5Љ�2�d��3��CE�- ���� $KAR��QM��TPDRA8)�����VECn@���IU��6��HE�f�TOOL�C2Vv�DRE IS3ErR6��@ACH��� 7?Ox �Q�2�9Z�H I�  �@$RAIL_B�OXEwa�RO�BO��?��HOWWAR�1�_�zROLMj��:qw��jq� �@ O_Fkp! d�l>�]9�� �R O8B�: �@�c�O%U�;�Һ�3ơ�r|�q_�$PIP��N&`H�l�@��~#@CORDEDd��p >f�fpO�� �< D ��OB ⁴sd���Kӕ����qSYS�ADqR�qf��TCHt�� = ,8`ENTo��1Ak�_{�-$xCq7�f�VWVA��?> �  &���PREV_RT~�$EDITr&_VSHWRkq��(� &R:�v�D��JA��$�a$HEA�D�6�� �z#K�E:�E�CPSPD.�&JMP�L~��0R*P��?��1%&�I��S�rC�pNEx; �q�wTICK�Cb��M�13�3HN��@ @� 1Gu�!�_GPp6��0STY'"xLO��:�2|l2?�A t 
m MG3%%$R!{�=��S�`!$��w`��Ȃճ���Pˠp6SQ�U��E��u�TER�C�0��TSUtB ����hw&`gw��Q)�pO����@I�Z��{��^�PR`�kюB1XPU��ΞE_DO��, XS:�K~�AXI�@���UR�pGS�r� �^0�&��p_) �EET�BPm��o��0�Fo��0A|����Rԍ��a<�S=R�Cl>@P� �b_�yUr��Y��yU�� yS��yS���UЇ�U�� �U���U�]��Ul[��Y�bXk�]Cm������YRSC�� 7D h�DS~0��fQ�SP���eATހ��A]0,2N�AD�DRES<B} S�HIF{s��_2C�H�p�I��=q�+TVsrI��E"����a�Ce�
��
;�V8W�A��F \��qA��0l|\A@�rC��_B"R{zp�ҩq�T�XSCREE�Gzv��1TINA����t{�XQ�A�b?�H T1�ЂB��р��I��A��BE�y RRO������ B��D�: �UE4I ��g�!p�S��RSyM]0�GUNEX(@~Ƴ�j�S_S�ӆ�� Á։񇣣�ACY��0� 2H�pUE�;�J�����@GM�T��Lֱ�A��O^	�BBL_| W8�N��K ��0s�OM��LE/r��� TyO!�s�RIGH���BRD
�%qCKG9R8л�TEX�@��>��WIDTH�� ��B�|�< �U�I_��Hi� L 8K���_�!=r���R:�_��Y�1R�O6q�Mg0璴�U��h�Rm��L�UMh��FpERV�w��P���`�Nz��&�GEUR��iFP)�)� LP��(RE%@�a)ק�a�P!��f �5�6�7�8Ǣ#B�É@����tP�fW�S@�M�USR&�O <����U�Qs��FOC)��PRI�;Qm� :���TRI}P�m�UN��
��Pv��0��f%�p�'���@�0 Q�\���AG �0T� ��a>q�OS�%�R Po���8�R/�A� H�L4N���U¡��SU�g��¢5��OSFF���T�}�=O�� 1R���:��S�GUN��}6�B_SUB?Ҝ��,�SRTN�`TU0g2��mCOR| D�'RAUrPE�TZ�#'��VCC��	3V �AC36MFB�1f$XRPPG ��W (#��ASTE�M�����0PEt��T3G�X �\ ��MOVEz�<���AN�� ���M���LIM_X��2�� 2��7�,�����ı�
��VF�`E���~�d�04Y��IB�7���5S��_Rp� 2���� WİG�p+@��}СP��3�Z�x ���3 ���A�ݠCZ�GDRID����Vy0�8�90� De�MY_UBYd���6��@���!��X��P_�S��3��L�KBMv,�$+0DEY(#�EX`�����UM_�MU� X����ȀU�S�� ���G0`PACI���а@��:���:,�:����RE/�3qL�+��:�[��TARG��P��r��R<�\ !d`��A��$�	��A�R��SW2 ��-$��@Oz�%qA7p��yREU�U�01�,V�HK�2]g0`�qP� N� �EAM0�GWOR���MwRCV3�^ ���UO�0M�C�s	�8��|�REF_�� �x(�+T� ����������3_RCH4(a�P�І�hr�j�NAۑXQ��0�_ ���2����L@��n�@@OU~7w6����Z��a2[��RE�p�@;0\�c�a'2]K�@SUL��]���C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��Q5(I�]7q�}�Tg`4D�`�0.`0�AP_�HUC�5SA��CMPz�F�6�5�5�0_�aR��a�1I\!�X�9|"GFS��a/d ��M��0p�UF_x��B� ���,RO��Q��'����UR�3GR�`.�3AIDp���)�D��;��A��~�IN��H{D���V@AJ���S͓UWmi=������TYLO*�5�����bt +��cPA� �cCACH�vR�UvQ��P�Y��p�#CF�I0s�FR�XT���Vn+$HO����P!A3� ��XBf�(1 ���$�`�VPy� ^b_SZ�313he6K3he12�J�eh chG�chWA��UMP�j��IMG�9uPAD�iiI�MRE�$�b_SI�Z�$P����0 ��A�SYNBUF��V�RTD)u5tqΓOLE_2DJ�Qu5RJ��C��U��vPQ�uECCUlVE�MV �U�r�WVIR9C�aIuVTPG����rv1s��5qMPLAHqa��v�V0�cm}� CKLAS�q	�Q�"��d  ��H�%ӑӠ@}¾�$�Q���Ue |�0!�rSr�T�#0! �r��iI��m�vK�BGf��VE�Z�PK= p�v�Q�&�_HO�0>��f � >֦3x�@Sp�SLOW>��RO��ACCE0���!� 9�VR�#���p:���AD�����PAV�j�� D�����M_B"���^�J�MPG ��g:�#E$SSC�����vP$q��hݲvQS�`qV�N��LEXc�i# T`�sӂ��Q��FLD �DEsFI�3�02���:���VP2�Vj� ��A��V�4[`MV_PIs��t����A�@��FI��|�Z ��Ȥ�����A���A���~�GAߥ1 LOO��1 JCB���Xcx��^`�#PLANE��R��1F�c�����pr�M� [`�噴��S����f����Af��R��Aw�״tU��pR�KE��d�VANCp�A���� k��q�ϲ�BR_AA� l��2� ��p�#Hć�m h���O !K�$������kЍ0SOU&A�"A�
pցpSK�TM@FVI=EM 2l ��P=���n <<��d^K�UMMYK1P�j�`D�ȡ��CU��#AU��o� $��TIT��$PR����OP����VSHIF<�r�p`J�Q�sԙ�fOxE$� _R�`U�#����s�� q������G�"G�޵r'�T�$�SCO{D7�CNTQ i�l�> a�-�a�;�a�H�a�V�P��1�+�2u1��qD����  � SMO�Uq��a�YJQ�����a_�R�[�r�n�*@LIxQ�AA/`�XVR���s�n�TL���ZABC�t�t�c��
AZIP��u,���LVbcLn"�}L�ZMPCFx�Mv:�$�� ���?DMY_LN����8���@y�w Ђ(a\�u� MCM�@Cbc�CART_�DP~N� $J71D��=NGg0S�g0�BUXW� ��U�XEUL|B yX���	������x 	���m��YH�Db  y� 80���0EIGH�3n�?(� H��9��$z ���|�,����$B� Kd'���_��L3�RVS�F8`���OVC�2@'�$|�>P&��
q�4��5D�TR�@ �9Vc��SPHX��!�{ ,� *<��$R�B2 2 ����C!�  �L� V+@b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/ ?�/�/V(7%3@/R/ d/v/�/6?�/�/�?�?@�?O4OOION;4]? o?�?�?�?SO�?�?�O�_�O0_Q_8_f_N;5 zO�O�O�O�Op_�O_ o8o�_MonoUo�oN;6�_�_�_�_�_�oo %o4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8����� Ǐ=�_�n���R���şx��ڟN;G � џ�
�� ����W�i�{����� ��ï�.�������A��dW�<�N�|� ������Ŀֿ�ޯ� ��0�B�_�R�d�� �϶������������ �*�L�^��rτ�
� �����������&�p8�J�l�~� `ҟ @�з��������-����&�,� ��9�{�����a��� ������������A 'Y����� ����a#�1�
��N;_MO�DE  ��S ��[�Y�AB���
/\/*	|/��/R4CWORK_{AD�	�
�T1/R  ���� ��/� _INTVA�L�+$��R_O�PTION6 ��q@V_DAT�A_GRP 2,7���D��P�/~? �/�?�9��?�?�?�? OO;O)OKOMO_O�O �O�O�O�O�O_�O_ 7_%_[_I__m_�_�_ �_�_�_�_�_!ooEo 3oioWoyo�o�o�o�o �o�o�o/e S�w����� ��+��O�=�s�a� ������͏���ߏ� �9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_T�IM����ΑR� ��Ƙ/��5�;#�U!P"�1!���  �?E�W�i�{�����.��ïկ�����'(~�T"2F���dR�I�Y��2�o+@a얿����)�u���� k0ϴ��_ ��  T� � ��2�D�)�T D��Q�zόϞϰ����� ����
��.�@�R�d��v߈ߚ�/V凷�����߽��R�_;�o �W��p��
�t���Diz$� �0 � �T"1!��� ������������ ��*�<�N�`�r��� ������������ &8J\n��� �����"4FX ��࿁�� �����/`4� =/O/a/s/�/�/�/�/ �/�/�!!/ �0޲k� ݵu�0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ ok$o6oHoZo lo~o�o�o�o�o1/�o �o 2DVhz �/5?������ ��&�8�J�\�n��� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-��?�Q�c�u��� �� ��`Ò�ϯ���� )�;�M�_�q������� ��˿ݿ� ����\3� ���&2,���	12345�678v�h!B_!��2�Ch���0�ϵ����� �����!�3�9ѻ�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� h�K߰���������
� �.�@�R�d�v����� ���������* <N`r���� ���&��J \n������ ��/"/4/F/X/j/ |/;�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�/�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_�? L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o=_�o�o�o�o�o �o 2DVhz@�����h��� ���u�o.�@�R���Cz  B��_   ���2&�_ � _�
����  	�_�2��Տ����_�p������ďi�{� ������ß՟���� �/�A�S�e�w����� ����N������+� =�O�a�s��������� Ϳ߿���'�9�K�"_������<v�_���$SCR_GR�P 1
� ��� t ���� ��	 �����������������_������)�a�����&�DE� D�W8���l�&�G��CR-35iA �90123456�7890��M-�20��8��CRg35 ��:�
��D�������������:֦�Ӧ�G���&������	��]�o������:���H���>��������@���&���ݯ:���j����g������B��t����������A����  @�`��s@� ( ?�=���Ht�P
��F@ F�`z�y� ����� �$ H��Gs^p��B��7�� /�0//-/f/Q/�/ u/�/�/�/8���P�� 7%?����"?W?-2<?<���]? �H�1�?t�ȭ7@�������?-4A, ��&E@�<�@G�B-1 3OZOlO-:HA��H�O�O|O P��B(�B�O�O_��E�L_DEFAUL�T  �����`SHO�TSTR#]A7RM�IPOWERFL�  i�/UYTW7FDO$V /UR�RVENT 1�����NU L�!DUM_EI�P_-8�j!AF_INE#P�_-4O!FT�_->�_r;o!��`o �*o��o!RPC_M'AIN�ojh�vo�oN�cVIS�oii��o�!TPpPU��Ydk!
P�MON_PROX	Yl�VeZ�2r���]f��!RD�M_SRV��Yg�O�!R��k��XYh>���!
�`M���\i���!RL�SYNC�-98|֏3�!ROS�_�-<�4"��!
C}E4pMTCOM����Vkn�˟!	��C'ONS̟�Wl����!��WASRCd��Vm�c�!��'USBd��XnR��� Noӯ�������!���E��i�0���WRV�ICE_KL ?�%�[ (%S?VCPRG1��-:"Ƶ2ܿ�˰3�	�"˰4,�1�˰5T�Y�"˰6|ρ�˰7�ϩϐ˰�����9���� ȴf�!�˱οI�˱�� q�˱ϙ�˱F���˱ n���˱���˱��9� ˱��a�˱߉��7� ���_������� ��)����Q����y� �'���O����w� �������� ˰��İd�c��� ���=(a s^������ /�/9/$/]/H/�/ l/�/�/�/�/�/�/�/ #??G?2?k?V?}?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O��O�O�O	_�O-_��_�DEV �Y��MC:5Xd��GTGRP 2�SVK ��bx 	�� 
 ,�PK 5_�_�T�_�_�_ o�_'o9o o]oDo�o hozo�o�o�o�o�o �o5{�_g�� �������� ?�&�c�u�\������� Ϗ���J\)���M� 4�q���j�����˟ݟ ğ��%���[�B� �f������ٯ���� ���3��W�i�P��� t���ÿ���ο�� �A�(�e�L�ί��R� ���ϸ������ �� O�6�s�Zߗߩߐ��� �������'�~ϐ�]� ��h�������� �����5��Y�@�R� ��v���������@�	 ��?&cu\� ������� ;M4qX���� ���/�%//I/ [/B//f/�/�/�/�/ �/�/�/�/3??W?� L?�?D?�?�?�?�?�? O�?/OAO(OeOLO�O �O�O�O�O�O�O�O_�iV �NLy�6� * 		S=>��+c"_VU@T�n_Y_B���B��2�J�j~Q��~_g_�_�Q%J?OGGING�_�^�7T(?VjZ�R{f��Y���/e�_%o7e�Tt�]/o�o {m�_�o�m?Qi�o�o�;)Kq%� �o�}os���� ��9�{`��)��� %���ɏ���ۏ�S� 8�w��k�Y���}��� ş���+��O�ٟC� 1�g�U���y������ �'����	�?�-�c� Q���ɯ����w���s� ���;�)�_ϡ��� ſOϹϧ�������� �7�y�^ߝ�'ߑ�� �ߣ��������Q�6� u���i�W��{��� ���=��M���A�/� e�S���w�������� ����=+aO ������u�� �9']��� M������/ 5/w\/�%/�/}/�/ �/�/�/�/=/"?4?�/ ?�/U?�?y?�?�?�? ?�?9?�?-OO=O?O QO�OuO�O�?�OO�O _�O)__9_;_M_�_ �O�_�Os_�_�_o�_ %oo5o�_�_�o�_[o �o�o�o�o�o�o!co H�o{��� ���; �_�S� A�w�e�������я� ��7���+��O�=�s� a������П���� �'��K�9�o����� ��_���[�ɯ���#� �G���n���7����� ����ſ����a�F� ���y�gϝϋϭϯ� ����9��]���Q�?� u�cߙ߇ߩ���%��� 5���)��M�;�q�_� ���߼��߅������ %��I�7�m������ ]�����������! E��l��5��� ����_D� we����� %
//���=/s/ a/�/�/�/��/!/�/ ??%?'?9?o?]?�? �/�?�/�?�?�?O�? !O#O5OkO�?�O�?[O �O�O�O�O_�O_sO �Oj_�OC_�_�_�_�_ �_�_	oK_0oo_�_co �_so�o�o�o�o�o#o Go�o;)_Mo ����o��� �7�%�[�I�k���� ������ُ���3� !�W���~���G�i�C� ���՟���/�q�V� �����w�������� ѯ�I�.�m���a�O� ��s�������߿!�� E�Ͽ9�'�]�Kρ�o� ������Ϸ���� 5�#�Y�G�}߿Ϥ��� m���i������1�� U��|��E����� ����	���-�o�T��� ���u����������� G�,k���_M� q����� ��%[Im� ��	���// !/W/E/{/��/�k/ �/�/�/�/	???S? �/z?�/C?�?�?�?�? �?�?O[?�?RO�?+O �OsO�O�O�O�O�O3O _WO�OK_�O[_�_o_ �_�_�__�_/_�_#o oGo5oWo}oko�o�_ �oo�o�o�oC 1Sy�o��oi� ����	�?��f� x�/�Q�+���Ϗ��� ��Y�>�}��q�_� ������˟���1�� U�ߟI�7�m�[�}�� ��ǯ	��-���!�� E�3�i�W�y�ϯ��ƿ ��������A�/� eϧ���˿UϿ�Q��� ������=��dߣ� -ߗ߅߻ߩ������� �W�<�{��o�]�� ��������/��S� ��G�5�k�Y���}��� ������������C 1gU������{ ����	?-c ���S���� ��/;/}b/�+/ �/�/�/�/�/�/�/C/ i/:?y/?m?[?�?? �?�?�?? O??�?3O �?COiOWO�O{O�O�? �OO�O_�O/__?_ e_S_�_�O�_�Oy_�_ �_o�_+oo;oao�_ �o�_Qo�o�o�o�o �o'ioN`9 ������A&� e�Y�G�i�k�}��� ��׏���=�Ǐ1�� U�C�e�g�y����֟ ���	���-��Q�?� a���ݟ��퟇��ϯ ��)��M���t��� =���9���ݿ˿�� %�g�Lϋ���mϣ� �ϳ�������?�$�c� ��W�E�{�iߟߍ߯� �����;���/��S� A�w�e��������� �����+��O�=�s� �����c��������� ��'K��r��; �������# eJ�}k�� ���+Q"/a� U/C/y/g/�/�/�// �/'/�/?�/+?Q??? u?c?�?�/�?�/�?�? �?OO'OMO;OqO�? �O�?aO�O�O�O�O_ _#_I_�Op_�O9_�_ �_�_�_�_�_oQ_6o Ho�_!o�_io�o�o�o �o�o)oMo�oA/ QSe�����%{,p�$SER�V_MAIL  �+u!��+q�O�UTPUT��$�@�RV 2��v  $� (�q�}��SAVE�7�(�TOP10 �2W� d O6 *_�π(_� �����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u�����`����Ͽݷ��YP���'�FZN_CFGw �u$��~����GRP �2�D� ,B�   A[�+qD;� B\��  �B4~�RB2�1��HELL�!�u��j�k�2���>��%RSR���� ���
�C�.�g�Rߋ� v߈��߬�����	����-�?�Q��  �_�%Q���_�슨�,p����)ޖ�g�2,pd��ﾆ�HK 1�� ��E�@�R�d��� �������������� *<e`r���?OMM ������FTOV_EN�B�_���HOW_?REG_UI�(��IMIOFWDL� �^�)WAIT���$V1��^�NTIM���VA�_)_UNIT�����LCTRY�B�
�MB_HDD�N 2W�  2�:%0 �pQ/�qL/ ^/�/�/�/�/�/�/�/��"!ON_ALI_AS ?e�	f�he�A?S?e?w?�: /?�?�?�?�?�?OO &O8OJO�?nO�O�O�O �OaO�O�O�O_"_�O F_X_j_|_'_�_�_�_ �_�_�_oo0oBoTo �_xo�o�o�o�oko�o �o,�oPbt �1������ �(�:�L�^�	����� ����ʏu�� ��$� Ϗ5�Z�l�~���;��� Ɵ؟����� �2�D� V�h��������¯ԯ ���
��.�ٯR�d� v�����E���п��� ϱ�*�<�N�`�r�� �ϨϺ���w����� &�8���\�n߀ߒߤ� O�����������4� F�X�j�|�'����� �������0�B��� f�x�������Y����� ����>Pbt ������ (:L�p�� ��c�� //$/ �H/Z/l/~/)/�/�/ �/�/�/�/? ?2?D?�V?]3�$SMON�_DEFPRO ����1� *S�YSTEM*0�m6RECALL �?}9 ( ��}
xyzrat�e 61 >14�7.87.149�.40:1253�2 =�=3148y �1�95172]?�O+M}�7�=2896 �?�?O�O�O�8Ctpdisc 0IO[@\OnO�O_�#_6Etpconn 0�=�O�O�O�_8�_1J�611 J_\_ n_�_o#o6OHOZO�_ �_�o�o�_�QJo\ono �o#6oHo�o�o�o ���o�oXj|� �2D������� ��T�f�x�	��.��@�ҏ������,�8�copy frs�:orderfi�l.dat vi�rt:\tmpback\I�[�y�
���/�/��mdb:*.*ԟ�����l��7�3x��:\H� ɠZ�[�s����(�;�4��aǯٯV���� ������ΟW�r���� '�:�տ^��ϓϥ� ��K�]���#�6� ����l��Ϗߡߴ��1 J�\�n߀��#�6�H�844 ������ ���J�\�n���#�26�?��602[��� �������9�9��ѿ@I�[�y�
/�0?� ��R�����8�H����V�t�) }5?������ ����Xs�/(/; �_�/�/�/�L ^��/?$?7�/�/ m�/�?�?��P/� }?O O3/E/�?i/�? �O�O�/�/V?�/yO
_ _/?A?�Oe?�O+_�_ ���Q_c_u_�_o*o=�O�192^��_o �o�o�_Jo\ono�ox#6�H�9308]���o���s�$S�NPX_ASG �2����q�� P 0� '%R[?1]@1.1��y?��s%�!��E� (�:�{�^�������Տ ��ʏ���A�$�e� H�Z���~���џ���� ؟�+��5�a�D��� h�z�����ů�ԯ� ��
�K�.�U���d��� ����ۿ������5� �*�k�N�uϡτ��� �Ϻ������1��U� 8�Jߋ�nߕ��ߤ��� �������%�Q�4�u� X�j��������� ����;��E�q�T��� x�����������% [>e�t� �����!E (:{^���� ��/�/A/$/e/ H/Z/�/~/�/�/�/�/ �/�/+??5?a?D?�? h?z?�?�?�?�?�?O �?
OKO.OUO�OdO�O �O�O�O�O�O_�O5_ _*_k_N_u_�_�_�_ �_�_�_�_o1ooUo 8oJo�ono�o�o�d�t�PARAM ��u�q �	U��jP�d9p�h�t��pOFT_�KB_CFG  ��c�u�sOPIN_SIM  �{�vn��p�pR�VQSTP_DS�BW~r"t�HtS�R Zy �� &!pINGS EL_5SEM����vTOP_O�N_ERR  �uCy8�PTN �Zuk�A:4�R�_PR�D���`VCNT_GOP 2Zuq�!px 	r��ɍ����׏��wVD��RP' 1�i p�y ��K�]�o��������� ɟ۟����#�5�G� Y���}�������ůׯ �����F�C�U�g� y���������ӿ�� 	��-�?�Q�c�uχ� �ϫ����������� )�;�M�_�qߘߕߧ� ����������%�7� ^�[�m������� ������$�!�3�E�W� i�{������������� ��/ASew ������� +=Ovs�� �����//</ 9/K/]/o/�/�/�/�/ �/�/?�/?#?5?G? Y?k?}?�?�?�?�?�?��?�?OO)�PRG�_COUNT8vq�k�GuKBENB���FEMpC:t}O_UP�D 1�{T  
4Or�O�O�O_ _!_3_\_W_i_{_�_ �_�_�_�_�_�_o4o /oAoSo|owo�o�o�o �o�o�o+T Oas����� ���,�'�9�K�t� o���������ɏۏ� ���#�L�G�Y�k��� ������ܟן���$� �1�C�l�g�y����� ����ӯ����	��D� ?�Q�c���������Կ Ͽ����)�;�d��_�q�=L_INFO� 1�E�@ �2@����������� �ٽ`y*��d�h'����¬��=`y�;MYSDEBUG�U@�@���d�If�S�P_PASSUE�B?x�LOG U ���C��*�Α�  ��A��UD1:\�ԘΥ�_MPC�ݵE&�8A��V� �A�SAV !�����l��X���SVZ��TEM_TIME� 1"���@ �0  3X���X�X����$T1?SVGUNS�@VE�'�E��ASK_OPTIONU@�E�A�A+�_DI���qOG�BC2_GRP 2#�I���~��@�  C����<Ko�CFG %�z��� �����`��	�.>d O�s����� ��*N9r] �������/ �8/#/\/n/��Z+�/ Z/�/�/H/�/?�/'? ?K?]�k?=�@0s?�? �?�?�?�?�?O�?O O)O_OMO�OqO�O�O �O�O�O_�O%__I_ 7_m_[_}__�_�_�X � �_�_oo/o�_So Aoco�owo�o�o�o�o �o�o=+MO a������� ��9�'�]�K���o� ��������ɏ���#� �_;�M�k�}������ ��ß�ן��1��� U�C�y�g��������� ������	�?�-�c� Q�s����������Ͽ ����)�_�Mσ� 9��ϭ�������m�� �#�I�7�m�ߑ�_� �ߣ����������� !�W�E�{�i����� ����������A�/� e�S�u�w��������� ����+=O��s a������� 9']Kmo �������#/ /3/Y/G/}/k/�/�/ �/�/�/�/�/??C? ��[?m?�?�?�?-?�? �?�?	O�?-O?OQOO uOcO�O�O�O�O�O�O �O__;_)___M_�_ q_�_�_�_�_�_o�_ %oo5o7oIoomo�o Y?�o�o�o�o�o3 !CiW��� ������-�/� A�w�e���������� я���=�+�a�O� ��s�������ߟ͟� �o�-�K�]�o�ퟓ������ɯ���צ���$TBCSG_G�RP 2&ץ�  ��� 
 ?�   6�H�2�l�V���z���@ƿ�������(��d�E+�?~�	 HC����>���G����C�  A�.�e�q�wC��>ǳ33��"S�/]϶�Y��=Ȑ� C\  Bȹ���B���>���X�P���B�Y�z�"�L�H�0�$���� J�\�n�����@�Ҿ ���������=�Z�%�07����?3������	V3.0�0.�	cr35��	*����
���0������ 3���4�   {�CaT�v�}��J2��)������CFG� +ץ'� �*������I����.<
 �<bM�q�� �����(L 7p[���� ��/�6/!/Z/E/ W/�/{/�/�/�/�/.� H��/??�/L?7?\? �?m?�?�?�?�?�? O O$O�?HO3OlOWO|O �O����Oӯ�O�O�O !__E_3_i_W_�_{_ �_�_�_�_�_o�_/o o?oAoSo�owo�o�o �o�o�o�o+O =s�E���Y� ����9�'�]�K� m�������u�Ǐɏۏ ���5�G�Y�k�%��� }�����ßşן��� 1��U�C�y�g����� ��ӯ������	�+� -�?�u�c��������� �Ͽ���/�A�S� ����qϓϕϧ����� ���%�7�I�[��� mߣߑ߳������߷� �3�!�W�E�{�i�� ������������ A�/�e�S�u������� ��������+ aO�s��e�� ���'K9o ]������ �#//G/5/k/}/�/ �/[/�/�/�/�/�/? ?C?1?g?U?�?y?�? �?�?�?�?	O�?-OO QO?OaO�OuO�O�O�O �O�O�O___M_� e_w_�_3_�_�_�_�_ �_oo7o%o[omoo �oOo�o�o�o�o�o !3�o�oiW�{ �������/� �S�A�w�e������� я�������=�+� M�s�a���������ߟ �_	���_ן]�K� ��o�������ۯɯ�� �#���Y�G�}�k� ����ſ׿������ ��U�C�y�gϝϋ� �ϯ��������	�?� -�c�Q�s�u߇߽߫� �������)��9�_� M����/����i�� ����%��I�7�m�[� ���������������� ��EWi{5� ������� A/eS�w�� ���/�+//O/ =/_/a/s/�/�/�/�/ �/�/?'?��??Q?c? ?�?�?�?�?�?�?�? O�?5OGOYOkO)O�O�}O�O�O�O�N  �@S V_R��$TBJOP_�GRP 2,�E��  K?�V	-R4S.;\{��@|u0�{SPU >�<�UT @�@LR	 �C� �Vf  C���U<LQLQ>�33�U�R�����U�Y?�@=��ZC��P���ͥR��P  Bq��W$o/gC��@g�dDb�^Ǚ��eeao�P&f�f�e=�7LC/�kaB o�o�P���P�efb-C�p���^g`�d�o�PL��Pt<�eVC\[  �Q@�'p�`�  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�ana�a`C�;�`L �w�aQoxp�x�p?:��XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb��� �X�	��1��)�W� ��c����������� �󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSocr35QT*��QT�A�� E��'E�i�F�V#F"wqF�>��FZ� F�v�RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG�G#
��D��E'
�EMKE����E�ɑE�ۘ�E��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF�u��<#�
<t���ٵ=�_��V �R�p�V�9� ]ESTPARbtp�HFP*SHR\�ABLE 1/;[I%�SG�� �W�G�G�G� WQ*G�	G�
G�GȖ�*QG�G�G�ܱNv�RDI~�EQ��@�Ϲ�������W�O_߀q�{ߍߟ߱���w�S]�CS !ڄ���� ��������&�8�J� \�n�������������  ]\�`��	��(� :�����
��.�@�w�~NUM  �E�EQ�P	P �۰ܰw�_CFG �0��)r-PIM?EBF_TTb��8CSo�,VERڳ-zB,R 11;[O 8��R�@2� �@&  �� �����//)/ ;/M/_/q/�/�/�/�/ �/?�/?J?%?7?M? [?m?>�@�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_H�_�_l_�Y@c�Y�MI_CHA�N8 c cDB'GLV��:cX��	`ETHERADW ?f�\`���?�_uo�oQ�	`R�OUTV!	
!��d�o�lSNMA�SKQhcba255.uߣ'9ߣ�Y�OOLOFS_�DIb��U;iOR�QCTRL 2$		�Ϸ~T�� ���#�5�G�Y�k� }�������ŏ׏������.��R�V�PE?_DETAI/h|z�PGL_CONF�IG 8�	����/cell/�$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c�u��� ��(���ϯ���� ��;�M�_�q�����$� 6�˿ݿ���%ϴ� I�[�m�ϑϣ�2��� �������!߰���W�@i�{ߍߟ߱�%}F� ������/�A�C�i�H�Eߞ������ ����?��.�@�R�d� v�������������� ��*<N`r� ������ &8J\n��! �����/�4/ F/X/j/|/�//�/�/ �/�/�/??�/B?T? f?x?�?�?+?�?�?�? �?OO�?>OPObOtO��O�O�O���U�ser View� ��}}1234?567890�O�O �O_#_5_=T�P��]_���I2�I:O�_�_��_�_�_�_X_j_�B3 �_GoYoko}o�o�o o�op^46o�o1 CU�ovp^5�o� ����	�h*�p^6�c�u����������ޏp^7R��)�;�@M�_�q�Џ��p^8� ˟ݟ���%���F��L� lCamera�J��@������ӯ���E~� �!�3��OM�_�q��������y  e��Yz� ��	��-�?�Q���u� �ϙ�俽���������>��e�5i��c�u� �ߙ߽߫�d������ P�)�;�M�_�q��*� <��i��������� )���M�_�q������ ����������<�û�� =Oas��>�� ��*'9K ]f�Q����� ��/�%/7/I/� m//�/�/�/�/n<� �^/?%?7?I?[?m? /�?�?�? ?�?�?�? O!O3O�/<׹��?O �O�O�O�O�O�?�O_ !_lOE_W_i_{_�_�_FOXG9+_�_�_oo (o:o�OKopo�o)_�o��o�o�o�o ��	g�0�oM_q�� �No����o�%� 7�I�[�m�&l�n� �Ə؏���� �� D�V�h��������� ԟ柍�g�ڻ}�2�D� V�h�z���3���¯ԯ ���
��.�@�R��� 3uF�鯞���¿Կ� �����.�@ϋ�d�v� �ϚϬϾ�e�w���U� 
��.�@�R�d�ψ� �߬����������� *���w���v��� �����w�����c� <�N�`�r�����=�w� �-�����*< ��`r�����������   ��1CUgy�������   -/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_�W_i_�  
��(�  �%( 	 y_�_�_�_�_�_ �_o	o+o-o?ouocoЙo�o�o�Z* �Q&�J\ n������o�� �9�(�:�L�^�p� ��������܏� � �$�6�}�Z�l�~�ŏ ����Ɵ؟���C�U� 2�D�V���z������� ¯ԯ���
��c�@� R�d�v�����᯾�п �)���*�<�N�`� �����ϨϺ������ ��&�8��\�n߀� �Ϥ߶���������E� "�4�F��j�|��� ����������e� B�T�f�x��������� ����+�,>P b��������� �(o�^p ������� / G$/6/H/�l/~/�/ �/�/�//�/�/?U/ 2?D?V?h?z?�?�/�`@ �2�?�?�?�3��7�P��!fr�h:\tpgl\�robots\m�20ia\cr35ia.xml�? ;OMO_OqO�O�O�O�O8�O�O�O ���O_ (_:_L_^_p_�_�_�_ �_�_�_�O�_o$o6o HoZolo~o�o�o�o�o �o�_�o 2DV hz������o �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟�ݟ��&� 8�J�\�n��������� ȯߟٯ���"�4�F� X�j�|�������Ŀ־:�8.1 �?@88�?�ֻ �ֿ�3�5�G�iϓ� }ϟ��ϳ�������� 5��A�k�U�wߡ߿���$TPGL_O�UTPUT ;|�!�! ��������,�>�P� b�t��������� ����(�:�L�^�p�Ђ����������23�45678901 ���������" ��BTfx��4������
} $L^p��,> ��� //$/�2/ Z/l/~/�/�/:/�/�/ �/�/? ?�/�/V?h? z?�?�?�?H?�?�?�? 
OO.O�?<OdOvO�O �O�ODOVO�O�O__ *_<_�OJ_r_�_�_�_ �_R_�_�_oo&o8o �_�_no�o�o�o�o�o `o�o�o"4F�o T|����\��}�����0�B�T��e�@������� ( 	 ��Џ�� ����<�*�L�N� `���������ޟ̟� ��8�&�\�J���n� ��������ȯ���"�������*�X�j�F� ����|�¿Կ��C��� ϱ�3�E�#�i�{�� �ϱ�S���������� /ߙ�S�e�߉ߛ�y� ����;�������=� O�-�s���ߩ��]� �������'����]� o������������E� ����5G%W} ������g��� 1�Ug	w� {��=O	//� ?/Q///u/�/��/�/ _/�/�/�/�/)?;?�/ _?q??�?�?�?�?�? G?�?O�?OIO[O9O O�O�?�O�OiO�O�O �O!_3_�O_i_{__��_�_�_�_�_�R�$�TPOFF_LI�M >�op:���mqbN_SV�`  l�jP_MON <6�Sdopop2l��aSTRTCHK' =6�f� b�VTCOMPAT�-h�afVWVAR� >Mm�h1d K�o �oop`b�a_DEFPR�OG %|j%�ZERO ZUZ�AUN	�j_DISPLAY`|n"r�INST_MSK�  t| ^zI�NUSER�odtL�CK�|}{QUIC�KMEJp�"rSC�RE�p6��btpscdt�q�h�b*�_.�ST�j�iRACE_CF�G ?Mi�d�`	�d
?�u�H_NL 2@|i����k r͏ߏ����'�9�K�]�w�IT�EM 2A�� ��%$12345�67890���� � =<��П�� G !���p�� =��c��^������� ���.���R��v�"� H�ί��Я������ *�ֿ���r�2ϖ��� ��4�޿�ϰ���&��� J�\�n���@ߤ�d�v� �ς������4���X� �*��@������ ��������T���x� ������l������ ��,�>�P�������F X��d������ :�p"��o �����F6H Zt~��N/t/�/ ��// /2/�/V/? (?:?�/F?�/�/�/j? �??�?�?R?�?v?�? QO�?lO�?�O�OO�O *O|O_`O _�O0_V_ h_�Ot_�O__�_8_ �_
oo�_@o�_�_�_ Lodo�_�o�o4o�oXo jo3�oN�or��o���s�S�B|���z�  h���z ��C�:y
 �P�v�]����UoD1:\�����q�R_GRP 1C���� 	 @Cp���$��H�6�l�Z��|�����f�৏˟���ڕ?�  
���<�*�`�N� ��r�������ޯ̯���&��J�8�Z���	��u�����sSCBw 2D� �� ���(�:�L�^�p�����|V_CONFIG E���@�����ϖ�OUTPU�T F�������6�H�Z�l�~� �ߢߴ���������� ��#�6�H�Z�l�~�� ������������� 2�D�V�h�z������� ��������
�.@ Rdv����� ��)<N` r������� //%8/J/\/n/�/ �/�/�/�/�/�/�/? !/4?F?X?j?|?�?�? �?�?�?�?�?OO/? BOTOfOxO�O�O�O�O �O�O�O__+O>_P_ b_t_�_�_�_�_�_�_ �_oo'_:oLo^opo �o�o�o�o�o�o�o  $����!�bt� �������� (�:�-o^�p������� ��ʏ܏� ��$�6� G�Z�l�~�������Ɵ ؟���� �2�D�U� h�z�������¯ԯ� ��
��.�@�Q�d�v� ��������п���� �*�<�M�`�rτϖ� �Ϻ���������&� 8�J�[�n߀ߒߤ߶� ���������"�4�F� W�j�|�������� ������0�B�S�f� x��������������� ,>Pa�t� �������(:L/x���k}gV�K� ��//&/8/J/\/ n/�/�/�/W�/�/�/ �/?"?4?F?X?j?|? �?�?�?�/�?�?�?O O0OBOTOfOxO�O�O �O�?�O�O�O__,_ >_P_b_t_�_�_�_�O �_�_�_oo(o:oLo ^opo�o�o�o�o�_�o �o $6HZl ~����o��� � �2�D�V�h�z��� �����ԏ���
�� .�@�R�d�v������� ��Ϗ�����*�<� N�`�r���������˟ ޯ���&�8�J�\��n���������Ż�$�TX_SCREE�N 1G�g�}ip�nl/��gen.htmſ�*�<�N��`ϽPanel setupd�}�dϥϷ����������ω�6�H�Z�l� ~ߐ�ߴ�+������� � �2�߻�h�z�� �����9�g�]�
�� .�@�R�d������� ��������}���< N`r��;1 ��&8�\ �������Q�ȾUALRM_M_SG ?��� �Ȫ-/?/p/c/ �/�/�/�/�/�/�/?�?6?)?Z?%SEV7  -�6"ECFG I嵻�  ȥ@�  A�1   ;B�Ȥ
 [?ϣ ��?OO%O7OIO[O�mOO�O�O�G�1GR�P 2J�; 0�Ȧ	 �?�O I�_BBL_NOT�E K�:T��lϢ�ѡ��0RDEFPR�O %+ (% N?u_Ѡc_�_�_�_�_ �_�_o�_o>o)obo�Mo�o\INUSE�R  R]�O�oI�_MENHIST� 1L�9  �(�0 ��)/�SOFTPART�/GENLINK�?current�=menupag�e,1133,1��oDVhz~�� }9361�� ���r�$�6�H�Z� l�~������Ə؏� ���� �2�D�V�h�z� 	�����ԟ���
� ��.�@�R�d�v���� ����Я�����9R q��B�T�f�x����� ����ҿ����ϩ� >�P�b�tφϘ�'�9� ��������(߷�L� ^�p߂ߔߦ�5����� �� ��$����Z�l� ~����C������� � �2��/�h�z��� ������������
 .@��dv��� ��_�*< N�r����� [�//&/8/J/\/ ��/�/�/�/�/�/i/ �/?"?4?F?X?C�U� �?�?�?�?�?�?�/O O0OBOTOfO�?�O�O �O�O�O�O�O�O_,_ >_P_b_t__�_�_�_ �_�_�_�_o(o:oLo ^opo�oo�o�o�o�o �o �o$6HZl ~i?{?����� �2�D�V�h�z��� �-�ԏ���
�� ��@�R�d�v�����)� ��П��������� N�`�r�������7�̯ ޯ���&���J�\��n����������$�UI_PANED�ATA 1N����ڱ  	�}�����0!�3�E�W� )Y�}� 7�뿨Ϻ�������� i�&��J�\�C߀�g� �ߋ�����������"�p4��X�7�� �q}�ϕ������� ��B����%�I�[�m� �����
��������� ��!E,i{b�������l� ܳ7�<N`r� ���-���// &/8/�\/n/U/�/y/ �/�/�/�/�/?�/4? F?-?j?Q?�?�?% �?�?�?OO0O�?TO �xO�O�O�O�O�O�O KO_�O,__P_b_I_ �_m_�_�_�_�_�_o o�_:o�?�?po�o�o �o�o�oo�o sO$ 6HZl~�o�� ����� �2�� V�=�z���s�����ԏ GoYo�.�@�R�d� v�ɏ����П��� ���<�N�5�r�Y� ������̯���ׯ� &��J�1�n����� ��ȿڿ����c�4� ��X�j�|ώϠϲ��� +��������0�B�)� f�Mߊߜ߃��ߧ��� ������P�b�t� ����������S�� �(�:�L�^����i� ���������� �� 6ZlS�w�'�9�}���"4FX)�}��l �����/j'/ /K/2/D/�/h/�/�/ �/�/�/�/�/#?5??�Y?��C�=��$UI�_POSTYPE�  C�� 	 e?�?�2�QUICKMEN  �;�?�?�0�RESTORE �1OC� � �L?��6OCC1O��maO�O�O �O�O�OuO�O__,_ >_�Ob_t_�_�_�_UO �_�_�_M_o(o:oLo ^oo�o�o�o�o�o�o o $6H�_U gy�o����� � �2�D�V�h���� ����ԏ���� w�)�R�d�v�����=� ��П������*�<� N�`�r�������� ޯ���&�ɯJ�\� n�������G�ȿڿ�x����7SCRE�0�?�=u1�sc+@u2K�3�K�4K�5K�6K�7�K�8K��2USER�-�2�D�ksMì�3���4��5��6��7��8���0NDO_?CFG P�;� ���0PDATE ����No�ne�2��_INF/O 1QC�@��10%�[���Iߊ�m� ���ߣ���������� >�P�3�t��i���<�-�OFFSET T�=�ﲳ$@�� ����1�^�U�g��� �������������$ -ZQcu���?��
����UFR�AME  �����*�RTOL_A�BRT	(�!EN�B*GRP 1�UI�1Cz  A��~��~��������0�UJ�9MSK � M@�;N�%8�%��/�2VC�CM��V�ͣ#RG�#Y�9���/�����D�BH�p,71C���3711�?�C0�$MRf2A_�*S�Ҵ�	����~XC56# *�?�6���1$k�5���A@3;C��. ��8�?��OOKOx1FODsO�5�51��_O��O�� B����A2�DWO�O7O_ �O8_#_\_G_�_k_}_ �__�_�_�_�_"o�O�FoXo�%TCC�#`�mI1�i�����n� GFS��2aZ;� �| 2345?678901�o�b �����o��!5aH�4BwB�`56 3~11:�o=L�B r5v1�1~1�2��}/� �o�a��#�GY k}�p������ �ُ�1�C�U�6�H� ��5�~���ߏ���	����4�dSELEC�)M!v1b3�VI�RTSYNC�� ����%�SIONOTMOU�������F��#bU���U�(u _FR:\H�\��A\�� �� wMC��LOG��   UD1���EX����' ?B@ ����̡�m��̡  OBC�L�1�H� ��  =	 1-� n6  -������[�,S�A�`O=��͗��ˢ}��TRAIN�P�b�a1l�
0d�$tj�T2cZ; (a E2ϖ�i��;�)�_� M�g�qσϕϧ���������	��F�STAOT dm~2@��zߌ�*j$i߾��_�GE�#eZ;�`�0�
� 02��H�OMIN� fU?��U� ~������БC�g�X���J�MPERR 2gZ;
  ��*jl� V�7������������ ��
��2�@�q�d�v�ZB�_ߠRE� hW�.�$LEX��iZ;�a�1-e��VMPH?ASE  5��c9&��!OFF/�FV�P2n�j�0�)�㜳E1@��0xϒE1!1?s33�����ak/�kxk(䜣!W�m[�䦲��[����o3;� [i{� ���/�O �?/M/_/q/��/� �//�/'/9/�/=?7? I?s?�/�?�/�/�?�? ?Om?O%O3OEO�? �?�O�?�O�O�?�O�O �O__gO\_�OE_�O �_�O�O/_�_�_�_o Q_Fou_�_|o�o�_�o o�o�o�o�o;oMo? qof-�oI��� ��7�[P� ��������ˏ�� !�3�(�:�i�[�ŏg��}������TD_F�ILTEW�n��3 �ֲ:���@�� �+�=�O�a�s����� ����֯������0�B�T�f�x���SH�IFTMENU [1o[�<��%�� ֿ����ڿ����I�  �2��V�hώ��Ϟ����������3�
�	�LIVE/SNA�P'�vsfli�v��E����I�ON * Ub�h�menu~߃������أ���p���	0����E�.�50�sU�P�@� ��Aɠ+B8z�z��}��x�~�P�� X���MEb���j<�0���MO���q���z�WAITDINEND��1����OK1�'OUT���SD��wTIM����o�G���#���C���b�������RELEAcSE������TM��������_ACT�[�����_DATOA r��%L�x���xRDISb�~E�$XVR��s���$ZABC_GRP 1t�UQ�,#�0�2�.��ZIP�u'��&����[MPC?F_G 1v�Q�!0�/� w��ɤ� 	�Z/  85�/�/H/�/l$?��+�/�/�/�?�/�/???r?�?  �D0�?�?�?@�?�?�;���x�|]hYLIND֑�y� ��� ,(  *VOgM.�`SO�OwO�O�M i? �O�O^PO1_�OU_<_ N_�_�O�_�_�__�_ �_x_-ooQo8o�_�o��oY&#2z� ���oC�e?a?�>N|�oq����qA��$DSPHERE 2{6M��_�;o ���!�io|W�i� �_��,��Ï���Ώ @��/�v���e�؏�� p����������ZZ�� �N