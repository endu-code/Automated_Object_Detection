��   u��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����UI_CON�FIG_T  �� A$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�62�ODE�
3�CFOCA �4VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�;s�� &USTOM~0 t $} RT_SPID�r,DC4D*PAG� �?^DEVIC�EPISCREuE�F��IGN�@$oFLAG�@ B��1  h 	$�PWD_ACCES� E �8���C�!�%)$LAB=E� $Tz ja�@�3�B�	B�USRVI 1  < `�B*�B���APRI�mx� t1RPTRIP�"m�$$CLA�@? ���sQ��eR��RhP\ SI��qW  ;�5�QIRTs1q_��P'2 L3hL�3!pR�	 ,���?����Q�PQ�R�T�Q����>�P� `�S�/o��
 ��)/�SOFTP.@/G�EN�1?curr�ent=menu�page,1133,18o�o�o�o��|Mo_o,1388vop/A �'�o�n9�o�����ocmc480|�%�7�I� �zQa�s��� ������͏\���� '�9�K�ڏo������� ��ɟX�����#�5� G�Y��}�������ů ׯf�����1�C�U���� TP�TX��y�򨑿o�� s �o���$�/softpar�t/genlin�k?help=/�md/tpia.d�gd����"�4��r&ɿۻpwd꿁ϓ� �Ϸ���������#� 5���Y�k�}ߏߡ߳� B�T�������1�C�V���zQf	bN� ($�ߕ�����p�����i zQ@�Q�c*oc����"�
)��Qa��
ae����  ��M	����@��n������P#`  ��V������SB 1��XR \� }%`REG VED�� �wholemo�d.htm4	si�nglEdou�b\trip�tbrows �@�!���� /AS|�/�Adev.sJlh�o�1�	t� ��w�G/Y/k/5/��/�/�/�/�/ ?� �P?*?<?N?`?r? �?�?�?�?�6�@?�? �?�? O2ODOE	�/ �/wO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_��_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -??z���� ���
��O@�R� !�3�����QOcOI� ݏ��*�%�7�I�r� m��������ǟٟ� ����_/�)�W�i�{� ������ïկ���� �/�A�S�e�w����� iֿ�����0�B� T�f�x�s��Ϯ�}Ϗ� ���ϭ�����>�9�K� ]߆߁ߓߥ������� ����#�5�^�Y�k� 9������������� ��1�C�U�g�y��� ������������ſ2 DVhz���� ����
��@R 	������� ��/*/%/7/I/r/ m//�/�/�/�/���/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSO!�O�O�O �O�O�O�O__0_+�T_f_5_G_�_�_�Z��$UI_TOPMENU 1�P��QR 
�d�QfA)*d?efaultqOZM�*level�0 *\K	 �o� So�_Qocbtpio[23]�(tpst[1�h�eo�ouo3oEo�-
h�58e01.gi�f�(	menu15&ypHq13&zGr�%zEt4M{4�a�� �������eB �C�U�g�y�����,��prim=Hqp�age,1422,1��ݏ���%� 0�I�[�m������2����class,5������)�4���130�f�x���h����5���53ʏ@���� �2�5���8ٯm��������4��ٿ����!�3�^I �P�Q�_k�m]��a[���ϝfty�m�o�aOmf[0�o��	���c[164�g.�5�9�h�a���k�Ax2 uK}��azmWw%{�� �sK�]�6�H�Z�l�~� ɿ������������  �2�D�V�h�z�	���2����������	�� ʟ?Qcu�( T�������Ѥ1$�N`r������ainedi�c����//��config=s�ingle&��wintpĀ /`/r/��/�/E�W��/{���gl[47��ow�?���!8��� 6�i.?h?>82ڀ??�?�?zl\rLz\r4s&x �? OVx`�6O��O�O �O�O�O�O��O_#_ 5_G_Y_k_�O�_�_�_��_�_�_,$;4$dokub?%o��13ؠ�&duali38�#�,4�_Pobo�_9 o,n'o9ato�o�o�o }_,>Pbt ���������� �o4�F�X�j�|����@��ď֏���=J�/ ,�wω¯���YOw���As�͔����ϡ�u�� l�V�ȟ.��?RO<���4�ߚ�6��u7���  �����/�A���e� w���������N����@��+�=�O�."$13�ϛϭϿ���ܿ ����+�=�O���s� �ߗߩ߻�����"�߀�'�9�K�]�����6 d��������,$۬74��/�A�S�e��C����?�	TP?TX[209�,����2�(��������1@I8��
����0P�2���1_�1�Y�tAv������0�
��1�
ïqC:4$treeviewA#�.f3�m381,26=o���l�� ��//+/�O/a/�s/�/�/�/�_B�5 $oq�?)?;?F/_? q?�?�?�?�?H?�?�?�OO%O7O�/�/�1��/r2V��O�O�O �6XO�edit 2azO�O_._@_�? ���OSL_�_�_�_~� �_�_G�o}o�Co Uogoyo�o�o�o�o/o �o�o	-?Qd uӥ������ ��?2�D�V�h�z��� ���ԏ���
��� �@�R�d�v�����)� ��П�������<� N�`�r�����%���̯ ޯ���&���J�\� n�������3�ȿڿ� ���"��_�_X�o|� �o��ϱ��������� �ߋ�)�S�e�x߉� �߭߿��ߓ��,� >�P�b�t￿���� ��������(�:�L� ^�p������������ �� ��$6HZl ~������ � 2DVhz� �����
/� ./@/R/d/v/�/7�I� �/m��/I���??)? ;?M?`?q?�?�/�?�? �?�?�?OO%O7O�� nO�O�O�O�O�O�O%/ �O_"_4_F_X_�O|_ �_�_�_�_�_e_�_o o0oBoTofo�_�o�o �o�o�o�oso, >Pb�o���� �����(�:�L� ^�p��������ʏ܏ /�/$��/H��?MO k�}�������ş؟� W����1�C�U�h�y� ����_Oԯ���
�� .�y�@�d�v������� ��M������*�<� ˿`�rτϖϨϺ�I� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F���X�|� ��������e������0�B�T���*defaulta��2�*level�8���������{� �tpst[1�]��ytpio[23���u������	m�enu7.gif��
�13�	�5��
��
�4�u6 �
ʯ?Qcu�� �����//� ;/M/_/q/�/�/�/6"�prim=�p�age,74,1��/�/�/??+?6"��&class,130?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO~O�O�O�O�/�"18�/�O_ _'_9_DON26@_u_��_�_�_�_��$U�I_USERVI�EW 1���R 
����_>��_
o�m (oQocouo�o�o<o�o �o�o�o�o);M _qo~��� ���%��I�[�m� �����F�Ǐُ��� ���.�@���{��� ����ßf������ /�ҟS�e�w�����F��*zoom��ZOOM��W�I�� $�6�H�Z���~����� ��ƿi����� �2��DϦ�maxres�H�MAXRES ߯E�㿬Ͼ������� ���*�<�N�`�߄� �ߨߺ���w������� o�%�J�\�n���5� �����������"�4� F�X�j��w������ ��������BT fx��?��� ���'=�t ����_��/ /(/�L/^/p/�/�/ ?�/�/�/7/�/?$? 6?H?Z?�/~?�?�?�? �?i?�?�?O O2O�/ ?OUOcO�?�O�O�O�O �O�O
__._@_R_d_ _�_�_�_�_�_sQ