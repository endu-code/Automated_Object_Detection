��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�� RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DIS�� S�MB�	"�BC�J@"CI2AI<P6EXPS�!�gPAR��TCL�/
 <(C�0��SPTM�E� PW�R��X�X�QoC l5��!�"%�7�ICC�%� kf�R�0leP� _DLIV��YNo3 �<oNbX_�P~#Z�_INDE
C�`O�FF� ~UR�iD���c�   �t �!�`MON��%sD�&rHOU�#EWA,vSq;vSqJv�LOCA� Y$�N�0H_HE����@I"/ 3 �$ARPz&�1FF�W_\ �I!F�`�;FA�Dk01#�H{O_� INFO�s;EL	% P K � !k0WO` $ACCE� �LVZk�2H#IcCE�L�V �$�s�# ���k���
���
`�K`SQi��  �5|�I�0ALh�z�'�0 ��
���F��p�����܅�$� 2ċ$b�w�������� č��!`r�Z���4���Ċ�!147.87.224.20h�S���96����܁�܁3�_{p_  �ċ� bfh.ch̟�1�C�U� g�y���������ӯ^��� _FLTR  l��π � �������n�nxč2�n��rSH�PD 1�ĉ  P!�
robstat�ion֯՚!k�.�Q�ſ������ ��޿?��c�&χ� JϫϽπ��Ϥ���� )���M��"߃�Fߧ� j��ߎ��߲���%��� I��m�0��T��x� ��������3���W� �{���P���t����� ��������Sw :�^����� �= a$Zׯm$ _L�A1��x!1.�ğP��1�Q2551.%�S���2��E �//*/<&3F/�� l/~/�/�/<&4�/�50�/�/??<&56?��0\?n?�?�?<&6�?�%@��?�?�?
O1�?P���MY� MY���c���� Q� �VN< �O�O_�O+_=_O_"_s_�_NPd_�_�_�_ �_�_o!o3o�_Woio{oVNLoM��o�l��oAo
.@U}�iRConnect: irc\t�//alerts E����Pu�@���1�C�Uу9P_R8�d��H�~� ������Ə؏����  �2�D�V�S$���8�(p����o͟ߟ�$�QA8��d�A��B4��j�h9�Q�+��@DM_�A�+��SMB 	 X�8%ğVO��߯����_CLNT 2
.X� 4C�ɯ0� �l�c�B�T���x��� Ͽ������)�;���_�q�Pϕ��MTP�_CTRL ��%���ϙdc���߀���?�*�c߳l��N���@{�Vߵ�Ƥ=�������ѓC���USTOM �{���}�@ |}�DTCPIPu��{��h�E�TE�L�{��A���H�!Ta�t�ç�roblolr� � ���!KC�L���F��!CRT��������!CONS&�$���n+���