��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����DRYRUN�_T   � �$'ENB �4 NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��SAW_� G �%$INIT�	RESUME_/TYPEN &J�_  4 �$($FST_IcDX�P_ICI�0 �MIX_BG�-A
_NAM�c MODc_U�Sd�IFY_TqI�.yMKR-�  $LI�Nc   �_SIZ�w� k. �, $USE_FL4 ��8&i*SIMA��Q#QB6'SCAmN�AXS+INS*}I��_COUNr�RO��_!_TM�R_VA�g�h>�i) �'` ���R��!�+WA-R�$}H�!{#�NPCH��$�$CLASS  ����01��5z��5%0VERS��.7  =�@2IRTU� .?�@0'/ l55�������Y0�6!m071�5��%71�?����?
O��}5I2�;�GOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_��%FW�?N8�0 ����_�_�_��@��o { 2�; �4%L_AND�_Bt_���QI���%L Jo��~:dLmu�%[oČo7g�1zo�o 
�X�o�o�o�o���p
Oa@� dvu�S���=�9Y0 ma`�s�1�t�a�r Y0�>�&�8�J�\�n� ��������ȏڏ��� �6�1��1 �2�D�V� h�z�������ԟ����
�44�6�S!2>�9 �[� m��������ǯٯ� ���!�3� �M�f�x� ��������ҿ���� �,�>�I�b�tφϘ� �ϼ���������(� :�L�W�p߂ߔߦ߸� ������ ��$�6�H� S�e�~�������� ����� �2�D�V�a� z��������������� 
.@Rdo�� ������ *<N`k}�� ����//&/8/ J/\/n/F