��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTTpe&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STPS_L�OG_P N��$��T�N�  �6 COUNT_D�OWN�$EN�B_PCMPWD� � DV�I�N!$C� C{RE�PARM:z� T:DIAG:�)�LVCHK|!FULLM0�YXT�CNTyD�MENU��AUTO,�FG�_DSP�RLS��U� &ENC�/  C�RYPTE  }���$$CL(   ���;!��� D 0 V� IO�� :&+ �}5L!IRTUA� �:/�$DCS_C�OD@���?%��  W�'_S � v*�!x �&��A91�"w!� 
 $B!���- �/? ?6?D?Z?h?~? �?�?�?�?�?�?�?OpO2O,#'SUP� ��+4OFO�#F�fOxO�O��  !�L�A���O � ��� V�[t&W��j���D�O N_��W
_��+!�U�U��YWALUGH 1}w) + �)�_�_�_oo)o ;oMo_oqo�o�o�o�' �_�o�o�o/A Sew����o� ����+�=�O�a� s���������ߏ� ��'�9�K�]�o��� ������Ə۟���� #�5�G�Y�k�}����� ��¯�����1� C�U�g�y��������� Я���	��-�?�Q� c�uχϙϫϽ�̿�� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� �%