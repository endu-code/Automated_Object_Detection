��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk"J 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A g /�C2�T�SST̀ 7���CH�r�F_�RVd�Ln�N�E2_�F�_�AC��_��C]q�2}��ck�_M&��DC�$_�V�3k�	V����W������d�q��d���RTN���i�T�A����AL�GO_S~�$P��a��x�REV_3IT!��MU�t�`CCCOF�Q>���X���GAM�PAS����_O�NTR���Fѐ��TR�V�CNPL��E���*�rtCNC`+1"�ZѐO�CHW�L��_�F-�r�;�d�OV�M/�QR�!֢�IO©�D���hע�JTHl#d�PA������PDA  i��DS�PVsCNMONL�S��*�w$8�RC��V<�P�KPGRI�j�RGfu�˔x��u�)O��g�T��O�Ae�Rvb����V�13���PD���AGWA֗�THӃ%��q3�aM��E����VRYac� �g�M��g���OVK���� /յ�;֧��VL^�!���cTCO���_�TR�/1u�MG�sI�o���.y@%a8INDE�sqϐTM9�זZC�C��ZRGCUSPF>����qp�ՇTWD�Ʊɖ�S�R��7t���O�L&�?��q<NS�K܀P`��sAXC�P_P�r+R�(SR��-DI7�-E�p�$J,E�RTY�LUFFIXE�sREG�1�����!F��Ѐ1sM����CNFC��EN��0�V��E�R�TV*TMU�R�G �4 Z��4 DU�?-'TS Y(**�@S�s�z%PQz$|z%IP/�4 AP���(�!IV]C2"N,�0P�M���!�н�#RC��(!8'�@QPY0H�5&B4��_sC3���r"[R_p�d`U��@VA}DCMVROU
b��1PERIO�sF31P���2D-��32%T��1_D��2H�ĺ3��T����K�95K��K�7CL����0�ADJ����_Uvdr�I�AUX�@��	 4�@C�P?a$� A�&�n@� qUX_AXS���P[PMC�� 
 h�D�rӠ �Cd��C�t�C�F�@�H��G1P�FOXp4XAX{ISU� Tj� �D͡Na�E��AP@M@� 	BQ܀HR
C$IDX\PRV�QSa��GRT�L ;$F�E_Uנ��=�TTOOL�R�p`;�Aѡp�y1DOf`� \��0R_P�KG�RQ BQ �NR�PBQS�P[Q H��R�P32�S�P2�Q�Q�ba	�1�ad�$VFLfw0IM�,�LT�r �:a��Tc�6Tb�����$DYG��C$d0JgGUg	�d�4�d��cMPSWP  ��$ @��  �����a�@&�@ &��`VERSION��h  ��5�aIRTUAaL�o�avS?�h&�  �a L|J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f��x��a+u|P11 29{\�@p��� ֓Ә�� � ?�a �@�@����A�   �����#����3��-�?�Q�?�g�U�����  D  Bp  =��Ϳ�??333?�a�̠d�̤@��ߥA ���/  & G�P� ?fffˡ>��ߥ�������0� ܙD���̤ˡ��k� C�Z�[��`�0�����Xӿٲ��B�ђǟ�I�ÿ��;���F�@ K���������Dz��l�W�I��ٺ��"ܑ�P`��w���ēV��'�9�K�]�o� 5ߓ���_�q�ۿ�� �����#�9�G�y�7� I�j�߳��������� ��a��!���y�3����ϋ�9�K�]�o� �ϓϙ���x���D�� ���������,> �b������� ����ɤ����ȗ�Đؓ� ��2/d���L����^/\�Ϣ�]�ĐW��"�@�"��'B������p���/"  $đƚ�$1>B,4_��(����1?��?�?�8>����ā�// @/�?T/f/?O�/�/�/ �/�/�/�O??,?>? P?b?;_�?__�?�?�? �?�?OO(O�_o^O pO�O�O�O�O�O�O�O  __$_�oH_Z_3~_��W��fx���2@�����	���o2�2-�V�h�z����� ��ԏ�������� Dqdd�����l��ߩߩ �b�����o����ğ���cd�p(�����(�qT�@� a>Ho��
}��[��c|�>L�Š���_v���<#�	
�Qsbp|��X��o�C��� a?e?a��3�T`��@ �G _�
�T���_����x�2bo%{Bta��������1��U�g�k�`>�X�ؤ����ϑ�Itk$ ��$$�>�٢	
���A��߭�'�x����4�+���s��.���Ճa$�{����(4$ܛռS�e�;��.��>���H�Ճa5�=���8M�Y��;��=���3��a�B�	 9�R�=�v�a�ߡ�� ��������m����  �b\'� �����`k�S�K�X�,� w�������/�����C���Q�??33�3;�s�<��saD/�  C``G�P /?fff/a>$��� ?_	W�_��0��_ g�;�5c?�4�'e��u�j� F@ ��[�� DzI ���w58���y ܃� ����/���/�/ 7I�_I/[/m//�/ �/�/�?�?�?�/?!? 3?E?W?i?{?�?kO}O�?�?�L�Oq�O� ������O���O �O�_
__._@_R_d_ o�_�_,o�_o�_�_ oobo%`&/ $.(��?��>� "��o����}��o��E +̰�B��+��ȴC� �8�����{j4�~gĠ {t��"�������$��3t7�q�����>���3t�cu� ��������� )�W���_�q������� ����ݏ�ȯ�%�7� I�k�%����j���ǟ ٟ���Ϳ3�E�W� i�{�a�������կ�L@�o0��������2Q /�A�S�e�v�Uώ�2�߲���������� �0�B�T�[Ru�� �������7M;	;	/� DO*GT�V� �M�D�i���Op�����������A>�a��f�p�B�BH���>L! �H���g�<#�
�ϲp��w�E�v������A��7������@\A�b� f��D?B,��7J���_���Bб���Z{@�p��N���>��4_�U�/��It$� //$��>�5
/a'A��a/	/�/-/�?&��+����%.�����%��$�=��%(4$��%�/��+;��.#5>���H/5��5���?58M�YK5��=@ g5��8�x?�+	�/ �?�?�?�7?�?O$O�6OHOZO�o�GnlG  ;¸`�X ���E�E��A��O��O�O	_�2 _^����`=�e?333����B�����D/ � C��G�P ?fff��>���e �Y�Q�iȌOVb�m�� ���W�i�]ooo�o���k��_wo�o�`F�@ uawU�`Dz�P$to�o�j"���� ��_�_o o'o�KoU�)��o �oﯥ����� 1���"�Y�k�}��� ����ŏ׏�ǟٟX�1��̸k��oC��o '9KQ���0�B� ��f�x���������z� ������l�>�P�b� t���lu�ς\�nπ��x�O������� 4�����C�<���R (����c�$�C � ���׺��ڷ  �� ��~Jk���_V�؏���/�?�Q�]�>�����]�������� ��+��O�a�s߅� ��U����������� ��9�K�$o���� ��������#�5� G�u�k�)�������� ������1ǼZ� ��/0/B/X%2�l�/��/�/�/�-��"2 �/? ?2?D?V?h?z? �?�?�?�d�n�>� GYGZ<���Y�Y��� ����ijO|O�O�O�FK �GLO^Ib!W
�#�> �'_��8��4U>L}PdQx�.B�<#�
K+p4_�B�t�FB�����SU�RkU@��lT��o� δ���ζ��0o��eB,TUPo�o�o�o �o��P>a�T�O�OrICIt$ Z�$�&>��R
k�wAHD�e���v��@+���+�.����7��A$敕G�(4$�S����;��.�>��yH���A5����O8M�Y���==dP Å�B�ԏ�{	�
� ��.��g�Y�n����������%o�=��ȗ  B��R�T_b �P#��J��X/�A�@S�e��|�j�B�	�y�S��?333�E�+��D7IcaD/  �CG�P ?fff�A>�Q8D��� �O=X蟲��M�O ���o��˿���?�Y�ӿ-�Kl�F@� _�k�ӥbl�Dz ���k�]�/��~!^/P) �;�M�_�q� ��Iߧ���s߅��� K��%�7�M�[ߍ� K�]�~���������� �!�3�u�#�5����Sl���)ϟ�M�_�q� �ϕϧϭ�GR����X ��������
�@ R�v����� ��/�ϸ����ȫ�� viڗ� N.k_=C��/o�㢄` s���U�"�d�Q�f�P cEci3�/6|P3$��ښ�$E>�Us��(���)o�<�?�8>�����:/-/?/Q/c/ u/�/`O�/�/�/�/? �O?)?;?M?_?q?J_ �?�?�_�?�?�?O#O �_7OIO"omOO�O�O �O�O�o�O�O_!_3_ oW_i_B�_{���z���u2	���H��.�F�2A� j�|�������ď֏� ����
�-�Xqxd�� ���l�����b���� �Ɵ؟���!�wd�p<������qh�T�_a>\��}z�o� s��>L٠�� o<��y<#�
�Q�b�p��/�l��o.�c���_aSeWa��G�h`ǥ@�Ȥ[s��T ���_�V�ꌿFbo9{B�a�����3�E�(�i�{�.k�>l���x��ϥ�It$ ��-$8�>��
���A�����;�����H��+��̇�.��y���G�$敕�Տ(4$ܯ�g�y�;���.��>��H���G�5����8'M�Y�O�=���G��a0�V�	M�f�Q� ��u��ߵ������� �����'��$�  �bp;����� �g�_�l�@����������C�����c��e<��S?333O����P���ñD/  C�t`G�P ?fffO�>8���Ss	k �_!xD�s{�O�I wS�'H;e#���/��j� F@ `��/o�� Dz]  ����I�q��y ܗ���� �//�/�/K]�_ ]/o/�/�/�/�/�/�? �?�??#?5?G?Y?k? }?�?�?O�OO�?g|�#O��O���� �/	_���O�O�__ 0_B_T_f_x_2o�_�_ @o�_$o�_oo,ovo�$%t:/&8B(�OPp\cҹ6��o�~ ǯ���o��E?��B Pp?��ܴW���L��� ���jH��gؠ�tPq6�@#������8�GtK������	��>��� Gt�w����� �����+�=�k�� s���������͏��� �ܯ'�9�K�]��9� ����~�ɟ۟���-� #��G�Y�k�}���u� ��ů���lD�������2eC�U�g�$yߊ�iϢ�2���� ������� �2�D�V� h�of���Դ���� ��KMO	O	C�XO>Ghπj"�4�a�X�}�Ӵ�И��������p�>�a��z��B�B\���>L5 \���{�<#�
��p������E,ϊ�����p������İ#@pA$�b�z�B�SB�@�KJ���s���B �n�������t >�Hs�i��*/�It$ C/$���>�I
#/u'A� �u//�/A/S&��+�����%.�����%��$敕�%(�4$�5�/�+;�{�.75>��HC5ޣ�5��S58M�Y_5��= {5��L��?�+	�/�?�?�? �7?O&O8OJO\OnO�}K�$CCSCH�_GRP12 2�����A&� \��|Xo��  O� �`�lt �E�E�� �A�__,_>_�2U_�C^����`Q�e?333��R����#�D/  CаGÿP ?fff��> ���e�Y�Q�}��O jb�m����W�i��o �o�o���2o�o�E`F@ 8uDa�U�E`Dz�PYtDo6��j6��� � o&o8oJo\o"��o� L�^��o�o���� �&�4�f�$�6�W��� ����ď֏����N� �����f���� x�&8J\n��� ��e�w�1�������ѯ ������+���O��� s��������u�Ϸ0�ϣϵϿxȄ��� ٳ.��i�'�#��x� q�H��R<L������ 8�W� ���� �4 ����J���sLV�����/�t����>����Ē��� ��*�<�N�`�9��� �ߨߺ��ߊ����� &�8�J�#n��Y�� ���������"�� F�X�j�|�����^�� �������0B/ f�����S/e/w/�%�2�l�/�/�/�/=�22?C?U?g?y? �?�?�?�?�?�?�d�n N1!Q|Y|Zqȝ�Y �Y�՟����i�O�O�O�O�FP� W�OP�I�!AW-3�>5��\_�S�H��iU>�L�P�Q�cB�<#�
�`pi_RE�8�V<B���, 0�U bA�U@푡T 4�Lo��В�fȚeo��Ba�U�o �oBT�P�>Ea�T�O�O�~CI�t$ �$6>��R
��wA}D������v!P+��̞`�.���l� Q$�敕|�(4$�x��@�R�;��.���>��H�� Q5{��Ѕ8M�Y܅(M=�P�� R�	�/�	&�?�*�c�N����� ����ǟٟ�Zo Mؾ>��  �I� b�T�b�PX�@�8JE� hd�v�����������<B�>��S,�?3�33(U`�)TlI�aD�/  CMG�P_ ?fff(Q>a mD,�L�D����� L�TM(_"�P�,� � !��?���bπ��F@ �Š��Hb��Dz6��Ġ���d�p"ʳ!�/�) �p� ��������~�ܿ�Ϩ� ��$�6π6�H�Z�l� �ߐ��߀������� � �2�D�V�h��X�j���������^��� �ϔϦϸ�������|R �������	-? Qu���� ��O��M/���/����) 5 �i���.�_nC��/ ����`��) e�"�d 0a�f%`�E�ih!?k �Ph$)!��$z>�U��8 $$�^o�<�?�8>��� $�:P/b/ t/�/�/�/�/�O�/�/ ??D?�OL?^?p?�? �?�?_�?�?�_ OO $O6OXOolO~OWo�O �O�O�O_�O�o _2_ D_V_h_No�_�_w�_�l�/����u2@>��.�@�R�c�B{�2v�����ÏՏ� ����/�A�H�?�b� �q�dةت�l$�(�(� r1��AC����:�1�V��d�pq�ݟ�(�q����Ia>����S}���5sť>L����5o��Ty<#�	
�Q�bpůd���c�����Ia�e�a�|��`��@I���� ��Sd,�o۶$���{bLon{B�a��Gπh�z�]Ϟϰ�ckM�>���!�L�B��ړItk$ �$m�>�"�	
��N�AٔN���p�x�,�}�+��̼��.�����|�$�{����(4$��ռ�߮�;��.�>���H�|�5�=�,�8M�Y8儝�=��T�|�%qe��	 �ߛ���������� �#�5�G���\�4Y�  (r�p� E��M���������u� ��������x��������*��?33�3����ș��D/�  C�`G�P /?fff��>m�ɔ ��	��_Vxy�C� ����~���J\}�peX��d��j� F@ ��d��� Dz� $���~8���y ��� ��/8B/?? ���_�/�/�/�/�/ �/?�?�?OF?X?j? |?�?�?�?�?O�O�OEOO�L�XO�0_� �//&/8/>_آ_ /_�_S_e_w_�_�_�_ go�_�_uooYo+o=o Ooao�oY%�o/I[mw(�<O�p�c� k�!�~��Γ0)� U t�R�pt�P�Č� 0Ɓ������j}��g� �t�qk�X�֎L�m��|t�ߺ�,�>�J�>���|tJ���� �����<�N�`� r���B�����̏ޏ�� �ۯ&�8��\�n��� ����n�ȟڟ����� "�4�b�X��|����� ��į��������p�@Gy��/�E�2� xߊߜ߮߿�����2������1�C�U� g�y�������� 	�4	4
)̀M�	�	x� �OsG�ϟW�i��������8���9�K�O����� Q>�a��pR R��!>Lj �Q����<#�
8��p!���EaϿ����� Q��@���X@�AY�b ��w��Bu�7�Jײ����B�A=��@���/��� >��}����_/6�It$� x/$��>�~
X/�'A5��/R/�/v/��&��+���5.����$5��$�=�45(4$�@5�/�
;;��.l5>���Hx5��5����58M�Y�5��=@Q �5����?�+	�/ �?�?OGT?FO[OmO�O�O�O��n�G  ��p�� L� U�E���A�_�._@_R_�2i_W^�����`��e?333���R��$�XD/ � C�G�P ?fff��>�-��e i�Q<����O�b}� ���Wy��o�o�o̵���Fo�o8�Y`F�@ LuXa�U Y`Dz�PmtXoJ�jk�K�=� �(o:oLo ^opo6��o�`�r��o �o8�� ��$�:�H� z�8�J�k�����Ə؏ ���� �b��"���z�4������:L ^p����4y��� E�����ӯ���	�ÿ -�?�ѿc��������� ��ϵu���Ϸ����xȘ����c�G }�;�X&�υ�\��R q`������m�� � P�P ���#�i  � ���J��2�`V������/����>����Ħ���,�>� P�b�t�M��ߪ߼��� �ߞ���(�:�L�^� 7���m�������� ��$�6�Z�l�~� ������r������  DV//z��� ��g/y/�/�%2�l�/��/�/
?=�322 .?W?i?{?�?�?�?�? �?�?�? t�nNE!e �Y�Z�ܝ�Y�Y�� ϗ��i�O�O�O�OVd� )W�O�I�!UW
A3L>I�p_-g�8\��}U>L�P�Qx�wB)<#�
�tp}_RY��VPB��L@D�U4bU�U@��TH�`o/ ����fܚyo3&+Bu�U�o�o 2 Vh`>Ya�T�_�O��CIt$ Z�$%6>��R
��A�D��(���v�5P+���t�.������4Q$敕��(4$ܜ�T�f��;��.ȅ>��yHԅ4Q5���O8M�Y��<M=�P �4R��C�	:�S� >�w�b�������ɟ۟����noM��  �]�(b�T�b `l�T�LJY�-hx���@����0�ů��PB�R�y�S@�?333<U�t�=T�I�aD/  �CaG�P ?fff<Q>%a�D@�`� X��(1���`�hM<_ 6�d�@��5�(Oࢿ�vϔ��F@� �Ŵ��\b��Dz J��Ĵ���x�6��!�/�) ܄������� ̿����ϼ���8�J� �J�\�n߀ߖߤ��� ��������"�4�F� X�j�|��l�~���������r����ϨϺ� ���������R����� /ASe� �-��� c�a/'�//%//����= I�i#�� �.�_~C��/��,��` ��= ,e2�dDa�f9` �E�i|5?�P|$=!�#�4�>e��%84$�8�ro�<�?H>���4$Jd/v/�/�/�/ �/�/�O�/??*?X? �O`?r?�?�?�?�?�_ �?�?�_O&O8OJOlO &o�O�Oko�O�O�O�O __�o4_F_X_j_|_ bo�_�_��_(l�1/����u2R�0�B�HT�f�w�V��2�� ��ŏ׏�����1� C�U�\�S�v��q�d� ��l8�<�<�0rE�+� UW��!�N�E�j��d�p���������]a>�̯g}���Is٥>L"�	�Io<Ӓhy<#�
�Q�b�pٯx���w�����]a�e�a�����`�@]�����g/d @�-o�8�տ�b`o�{B�a����[�|ώ�q�����wka�>��5�`�xV���It$ 0�-$��>�6�
�b�A�b�
߄�.�@֑��+�����.��y��Ր�$敕�Տ(4$��հ���;���.$�>��H�0吡5��@�8'M�YL嘝=	�h���9qy��	�߯�� �������%�7�I��[�j��$CCSC�H_GRP13 �2������&� \��~E�y   <r���Y��a����� ������+��(B0����>��?333����ܙ��D/  C�`G�P ?fff��>��ᔜ�	��_jx ��W�ĝ������ ���el���<�j2F@ %%1���2Dz� F$1�#/��#���y �%7I?m w/9?K?���_�/�/ �/�/?!?S?O#ODO {?�?�?�?�?�?�?�?@;O�O�OzOSO\��O �e_/%/7/I/[/m/ s_�R_d_o�_�_�_ �_�_�_�ooo�o<o �o`oro�o�o�o�%�`�/~���(�qO �p�cɠ�V��ޓ e^�5U�)�9R�p�� ��%Ġ�Dƕ����j ���g!��t�q�����`�9���t��οa�<s��>����t� ����)�;�M�&� q�������Տw�ݏ� ��%�7��[�m�F� ������ǟ韣���� �3�E�W�i�����K� ��ïկ���߿�/� �S���|�@�R�d�z�2��߿�������	���2�0�B�T� f�x��������� ����>�i	i
^̵M �	�	���O�G����� ��������=�m��n�����.�ڱ>�"qI��@R5R��V�>L� �ƿP���<'#�
m�M�pV��p2U����)���ڱ@��u.��@�A �!r9�Ϭ��B��l �JR�ݿ��BN�v r��/�//A/��� >2������/k�It$ �/$��>%��
�/�'Aj��/��/?�/�& +��=�M5.���Y5�$敕i5(4$��u5-??;;��.��5>��H�55����58M�Y�5�=� �5���?;	?,OOPO;G�? {O�O�O�O�O�OG��|�n�G  �� 6p��� EU-U%� 2QQ_c_u_�_	B�_��^)��+p�u?333MRY���D/  C:�GÿP ?fff> �Z�u9i1aq���
_ �b9}A�g=y/�o �o���{o�oOm��`F@ �u�a�U5�`Dz#`�t�o�Qz�р�r� � ]ooo�o�o�ok��o� ����#m�#�5�G� Y�o�}���m����׏ �����1�C�U��� E�W�֟��i���K ��o�����ϯ i����z������ ,�>���b�t�Ϙ�� ��ο��<��u:� �0��������͟� "Ø�G��pލW��� �ߑ�b������ �����U�� XǞ U���J��g���V���?K������>������=� O�a�s߅ߗߩ߂��� �����1���9�K�]� o���l������ ���#�E��Y�k�D ������������� 1CU;y�d/ ���
ߜ/�/�/�%�2+|	??-???P=//h22c?�?�?�?�? �?�?�?
OO.O5t,~ ONz!��Y�Z��i i	"��./0y�O�O'__CV�� ^W�OP�I�!�Wv3��>~���_@-����"#�U>�L�P�Q"�BA)<#�
��p�_QR��8�PV�B����u y�Uib��U@6��T }o@/��f��oh9[+B��U�o 4UgJ��P:`�>�ad9_/_��CI�t$ 	�$Z6>�b
�;�A�D;���]���jP+��̞��.�����iQ$�敕Ņ(4$�xх����;��.���>��H	�iQ5{���8M�Y%�qM=�PA�iR!R�x�	o���s������ן ����"�4��oIM!�>F�  "�� ]b2d�b:`�����J�� bh����ѯ�e����ʅB���cu�?3�33qU��rT�I�aD�/  C�G�P_ ?fffqQ>Za �Duŕ����C(f�0� �͝Mq_k���u7�I� j�]EO׿Qϫ���F@ ���Q��b�Dz�����ϭ�pk��!�/�) ܹ� ˿ݿ����%�/��� �m���ߑߣߵ� �����������3�E� W�i�{���������2�����E��� ��������%�+�R 
�@Rdv� �T��b�F *<N�FՖ/\�6/H/Z/d��)�r ~ �iX�/�.�_�C/? ��a�p��r ae=2�d yavn`�E�i�j?� �P�$r!X�E4�>9e�Z8i$m��oL+O7H>���i$7J�/�/ �/�/�/�/?�O)?;? M?_?�?/_�?�?�?�? �?�?�_O%O�_IO[O mOO�O[o�O�O�o�O �O_!_O_E_i_{_ �_�_�_�o�_�_�o�]l4/f/�
��2�2@��e�w��������Ă2�������0� B�T�f�x����ĈΫ� �q�d!�!�|m�q�q� erz�`����D�V���z����d%���&�8�(<��҃��>����}����~s�>L�W�>�~o��y<#�	
%arp�����N��������e�a-�Ų�`E�@��F�� �ddu�bo$�m�
��b�o�{Bq.�*ϐπ���Ϧ����Ϭk��>��j�����L�#�Itk$ e�$��>�k�	
Eߗ�A"���?߹�xc�u�Ơ+�����.����š$�{��!�(4$�-�����;��.Y�>���He�š5�=�u�8M�Y��͝�=>���Ţnq����	 ���������A�3�H� Z�l�~�������}��  qr��� ��9�����ݚ�� 	-?��VD����s��?33�3ͥΤ�E�D/�  C�`G�P /?fff͡>��� ��	�)o�x���� ��ͯ���ϓ����e��3�/%zFF@ 9%E��FDz� Z$E7/	/�8X�8�*� �' 9K]#?��/M?_? ��%o�/�/�/?'? 5?g?%O7OXO�?�?�? �?�?�?�?OOO�O_�OgO!\��O/y_'/ 9/K/]/o/�/�_!�f_ x_2o�_�_�_�_�_�_ �oo,o�oPo�oto�o �o�o�o�%��/����(ȅO�p�cP� ��j(�E��yr�IU �^�MR�p����Z�ձ y�ʰ=�=�zƏwV� ��q�������M����t���u�����>����t����� +�=�O�a�:������� ��鏋����'�9� K�$�o���Z�����ɟ ۟�����#���G�Y� k�}�����_�ůׯ� ����1�C��g���@��T�f�xߎ�2� ����������� �2�D�V�h�z��� �����������2� R�}	}
r��M�	�	�� �O�G�������������Q���������B.�9�>6q]��pTRIR��j>L� �ڿd���<#�
��a�pj	FU��=���9�-�1��!B��@�A�5rM �����B����Jf ���Bb����/@//C/U/�� >F�������/�It$� �/$�>��
�/�'A~��/�/?�/��&" +���a5.����m5!$�=�}5(4$܉5A?�S;;��.�5>���H�5!5����58M�Y�5)�=@� �5!��
O0;	'? @O+OdOOG�?�O�O�O��O�O�O[��n�G  ��Jp� �� YUAU9�FQe_�w_�_�_B�_�^=���?p�-u?333�)aR*m��D/ � CN�G�P ?fff)>n�-u MiEa����_�bM}U� )#gQy-/�o"����o	c�ʢ`F�@ �u�a	eI�`Dz7`�t�o�e#z���߆� �qo�o�o �o�o��o�����% 7��7�I�[�m����� Ï����������!� 3�E�W�i���Y�k��ß}����_կ�� �����}¯ԯ ����
��.�@�R�� v���Ϭ���п��� �P��uN���� �����*�6ìW �τޡk����ߥ�b ���*��Ҷ1� &���i�"�lǲ i� *�Z��{���V�!��%?_������>���!���Q�c�u߇� �߽߫ߖ������� E���M�_�q���� �������%�7� Y�m��X������ �����!3EW iO��x/��� ߰/�/�/�%2?|?�/?A?S?d=C/|22 w?�?�?�?�?�?�?O O0OBOIt@~cN�!� �Y�Z�%�)i)i"2� �B/Dy�O_;_2_WV�� rW�O�I�!�W
�3J>���_T-��8��6#�U>L`�Qx6�BU)<#�
��p�_eR��/dV�B��J���U}b��U@J��T�©oT/ -��f%��o|Mo+B��U�oHi{ ^��dN`>�a"d�M_C_��CIt$ Z�$n6>�#b
�O�A�DO��q��-��~P+��̽�.����Ʌ}Q$敕م(4$�兝����;��.�>��yH�}Q5��-�O8M�Y9��M=�P U�}R&!f���	���� ��������� ��$��6�H�W��$CCS�CH_GRP14 2���y��&� �\m.2�p)  )"��qbFd�bN`֥ ���Jávh�����Py�/���B���+c��?333�Uޢ�T|�I�aD/  C��G�P ?fff�Q>na�D��ʹ±� W(��D©ͱM�_���� �l�~ϟ�qYOφ�x����F@ �0����b�Dz��3Ԁ���Ϡ�1�/�) �� ��$�6��� Z�d�&�8�ϴ���� ������ ��@���� 1�h�z����������(�����g�@���� z���R ��$�6�H� Z�`�R?Qu� ������� ){M_q��{���/��k/}/�/��� ^�� �y��C/>�_ �CR/K?"��p&�  uer2t�a1v�`�E�i ��?�`�$�!��z4 �>Me&��8�$���oxNL`OlH>����$ lJ�/�/�/??(?:? _^?p?�?�?�?d_�? �?�? OO$O�_HOZO 3o~O�O�O�O�O�o�O �O�o _2_D_V_�_z_ 8�_�_�_�_�_�o
o o�@o�li/�/-�?�Q�g�2�̚�����Џ����2��/� A�S�e�w��������� �Ľ����+tV�V�K| �������r�������@y�������Ԧ*tZ�@�[�m�q����a>!6��}-"�sC�>L��s��o=��yO<#�
Za:rpC����������au
qb���pz�@ ��{�"&���d��o@YƢ�?��b�o�{B;q c�_����������.��k˰>���ʯ����^X�It$ ��$�K>���
z���AW����t��ߘߪ���+�{��:�.���F����$敕V�(4�$�b��,�;��=.��>��H�����5����8M�	Y���=s������q��	�	 ���=�(� v�h�}���������4��ڝ���   �r# �ôn�˰2 ��>Pbt��(�y�� ��%?333�:�F��z�D/  C'pG�P ?fff�>�G�%&^o�x ���&-.���*)� ����e֟h�</<Zz{F@ n%z�"�{Dz�$z�l/>/���m�_� �J\n��X?� �/�?�?�/Zo?"? 4?F?\?j?�?ZOlO�O �?�?�?�?OO0OBO@�O2_D_�O�OV\��O 8/�_\/n/�/�/�/�/ �_V��_�_go�_�_�_ oo+o�oOoao�o�o �o�o�o�o�o)�%'�`�/����(ȺO �s�����]�z�H� ���~U����R�� ΂��
�����r�r�Bz ��Ew��B����քT�ʵ���t��8Ϫ�<��Ș>����tȚ *�<�N�`�r�����o� ��̏ޏ�����&�8� J�\�n���Y������� ڟ����2��F�X� 1�|��������֯�� ����0�B�(�f�x� Qߜ�����ߛ߭���2,����,�=�	�U�2P�y��� ����������	��"$ .<�gчĲ	�
���M ��_�G�)�� ��0����K�������wc�#�>�kq�-݉R~Rӟ�>L� �ϙ�.�<'#�
����p�>p{U��=r���#�@b�f��Vw��@#Q �jr�-���R� �J�U�&�H�B��� �!/B/T/7/x/�/=�'>{�&�/��It$ �/$G�>%��
�/(7A��(?��/J?�/6W +��=̖5.����5V�$敕�5(4$�ܾ5v?�;;��.��5>��H�5V5���E8M�YE^�=� .EV��?Oe;	\?uO`O�O�G�? �O�O�O�O_!_�6�|~3W  � pJ�'�UvUn� {QO�_�_�_�_RB�_��^r��tpbu?333^�R_����D/  C��GÿP ?fff^> G��bu�iza��0�S_ r�}��^Xg�yb/$ 6WJ�2��o>����`F@ �u�a>e~�`Dzl`�t�o���Xz���߻� � �o�o�o�o�o��� ޏ��Zl��l�~��� ����Ə����ȟ� � 2�D�V�h�z������� ����������2�� 
����� ��� ���	�ÿ-�?�Q�c� u���Aϫ���O��3� ��)�;υ�3���I�0#�5�G�Q���_� k��EW�Ϲ����
� �ڥNb�ޢ_�N*� �f
&[�����W� ��� ��_�EZ2��&�VG�V�Z?���$�>���V�$��� �ߪ߼���������� (�:�L�z����� ������ ���6� H�Z�l���H����� ������<2�V hz������/ �J!�S��/�/	?5�2t|R?d?v?�?�=x/�22�?�?�?�?O O/OAOSOeOwO~tu~ �N�!�ij,Z�^i ^iR"g�M�w/yy1_C_p_g_�V�0�W_P%Y)1�W�3>����_�-�ڢk#�U>�LD`+ak�B�)<#�
�p�_�Rץ8;/�V�B��� �e�b�2e@�3d ���o�/Qb�OvZ��o���+B�e }�������`�>�aWd�_x_9�SI�t$ R�$�6>�Xb
2���AT��,��P�b��P+��̞�.������Q$�敕�(4$�x�ҏ�;��.F��>��HR��Q5{��b�8M�Yn��M=+`���R[!����	��џ������.� � 5�G�Y�k�}��o�Mj�>��  ^"�� �b{d&r�`�ҥ�Jס �h����,���C�1���B���`c��?3�33�U�T�I2qD�/  C�G�P_ ?fff�Q>�a �D��޹ֱ�(��y� ���M�_���ɾ�ϒ� �Ϧ�O Ϛ���*3�F@ &�2����b3�DzȰG�2�$���p��E1%?9 �� �&�8�J��n�x�:� L������������ �"�T��$�E�|�� �����������<�����{�T������f �&�8�J�\�n�tb Se����� ���=�a s������/��/�/�/���r�� � =y��W/>2o�Cf/_? 6��Kp:� �e�2Gt �afv�`*U*y��?� C`�$�!���4N�e:��8�$���obLtO�H>����$�J�/�/ ??*?<?N?'_r?�? �?�?�?x_�?�?OO &O8Oo\OnOGo�O�O �O�O�O�o�O_�o4_ F_X_j_�_�_L�_�_ �_�_�_�oo0o	�To��l}/�/A�S�e�{�2@�̮���ҏ�����2�1�C�U�g�y� ��������ӟ������ �?tj�j�_|������ �r������ɍ���̯ï�>tn��o���(��/���a>#!J���}A6�sW�>L࠰���oQ��y<#�	
naNrpW���3���*����auqv��/p��@��"" :���d��omƶ�S�r�o �BOqw�s��π�����0�B��k߰>�3���ޯԯ��l�Itk$ ��$��>���	
����Ak��߈��x�߾��+���N��.���Z��$�{��j�(4$�v�.�@�;��.��>���H���5�=���8M�Y����=������q���	 �-��Q�<���|��� ��������H�����  �r7 � ״��߰F.&�3� Rdv�
��*���, ��%?33�3�N�Z���D/�  C;pG�P /?fff�>��[� %:2ro�x�:- B��>)���/�u�|�P/nz�F@ �%��6Dz$�$��/R/*8����s� �^p ���l?��/�?�? /$/no$?6?H?Z?p? ~?�?nO�O�O�?�?�? O O2ODOVO�OF_X_�O�Oj\��OL/�_p/ �/�/�/�/�/�_j��_ �_{o�_�_	oo-o?o �ocouo�o�o�o�o �o�o=�%;�?���	8��O�#s�� ���q���`�����U ���R��₣�� �������Vz�Yw�� V�����h�޵������LϾ�Пܘ>����ܚ>�P�b� t���������Ώ��� �2�ԯ:�L�^�p��� ��m���ʟ��� �� $�F� �Z�l�Eϐ��� ��Ư��ꯨ�� �2� D�V�<�z���e߰��@���߯�����2,, 
��.�@�Q�0�i�2d���������� ����/�6$-.P�{� ���	�
��]
� _W/�1)����(D����_�������w�7�>q�A�p�R�R#ӳ>L� ��#ϭ�B�<#�
ʱ��p�R�U��Q����7�v�z��j���@7Q�~r� A�	�R��Z�i�:�\�B����5/V/@h/K/�/�/Q�;>��:0�/��It$� 
?$[�>�
�/<7A��<?�/^??�6k +��̪5.�����5j$�=��5(4$��5�?ޜ;;��.�5>���H
Ej5���E8M�Y&Er�=@� BEj�SOy;	p? �OtO�O�G�?�O�O�O�_#_5_D[�$CC�SCH_GRP1�5 2����fQ&� �\Z�]�  ғp^3�; �U�U���Qc�_�_�_�ofBo
n����p<vu?333r�R�s���D/  C���G�P ?fffr>[��vu�i�a οD؈_1r�}��r�g �yv/Yk�^�F��o�s���pF@ `�uqse�pDz�`  ����z������ ��o�o�o# �GQ��%���ʿ ����ŏ׏���-�� ���U�g�y������� ��ӟ�ïկT�-���g��?����#� 5�G�M��,�>���b� t���������v��� ���h�:�L�^�pϺπh���~�X�j�|߆��K��Р��zW0��� ���?�8���b � ��b_��z&o�� ��ʌ���� �Ԕ�zZ@g���:f|��n?�;�M�Y�>��� ��Y����������� '� K�]�o���Q ������������5� G� k�}�������} �����1Cq g%/������ �	�/-V߈�?,?>?T52�|�?�?�?$�?�=�/�22�?
O O.O@OROdOvO�O�O �O�t�~�N�!$CiCj 8,���i�i�"�����/��yf_x_�_�_�V$�G0�WH_ZY^1g�3�>��#o�-���#0e>Ly``a�*R��)<#�
G'"p�0o�R�p/�VR�����Oe�b ge@��hd���/�����Fv��,���+B (!PeL����	����`>q�d�_�_�n�ESIt$ ��$��6>��b
g���A�DT��a�ۏ�����P+����'�.����3��Q$敕C�(�4$�O���;�{�.{�>��H����Q5����8M�Y���M=``���R�!П��	���*� �c�U�j�|��������!�M��ħ  �"��b�d[r�`� ��J��h+�=�O�a�P�x�f�R���c��?333�U'��T|3YgqD/  C �G�P ?fff�Q>�a4T����K �(䯮��]�_�� ���������OU���x)�G*h�F@ [�0g�ϵrh�Dz��|Ԁg�Y�+���z1Z?L9 �7�I�[�m��E� �ϭ�o������G�� �!�3�I�W��G�Y� z��������������/�q�1����C� ��%ߛI�[�m�ߑ� �ߩCb��T�� ���<N� r�����/���?�ߴ/�/�/��� ��� �ry֧�/J>go 1S�/�?k߲�po�  �e�2|t�a�v�`_U_y /*�?2'x`/4�!֪�4 AN�eo��8�$�%x�L�O�H>����$ �J?)?;?M?_?q?�? \_�?�?�?�?O�_O %O7OIO[OmOFo�O�O |o�O�O�O�O_�o3_ E_i_{_�_�_�_�_ ��_�_oo/oSo eo>��o�l�/�/v�������2������*�	�B�2=�f�x� ��������ҟ���� ��)�T�tt�����| �����r�����
�@¯ԯ����st��@8�������d�P�q>X!��vk�s��>Lհ���o���O<#�
�a�rp���+�h�*�_����qOuSq��C�dpõ@ ĴW"o���d���o@������Br5�B�q �����/�A�$�e�w�*{�>h���	���^��It$ ��$4�K>��
���A�����7�����D�+�{�̃�.������C�$敕��(4�$ܫ�c�u�;��=.��>��H��C��5����8M�	Y��K�=���C��q,�R�	I�b�M���q� �����������}��#��    �rl 7�ķ��{c [�h<ȇ���?�(��_��a �O%?333K��L������D/  CppG�P ?fffK�>4���O%og�o� @
"o-w�K�Es)O� /#/D/7u��+/�/<�z�F@ �%�+k��DzY�$���/�/E*ց���� ܓ�����?� 	?�?�?G/Y/�oY?k? }?�?�?�?�?�O�O�O OO1OCOUOgOyO�O@�O{_�__�O�\�_ �/�_�/�/�/�/�/�/ o���_�_�oo,o>o Poboto.�o�o<�o  �o(r 5p�`6?�"�4�>8�_ L�Xs��2���ÿ�� ����U;���RL�;� ���S���H����ɋz D��w԰��L�2
�����4�C�G���<��>���C�� s���������͏ߏ�� ��'�9�g�	�o��� ������ɟ�����ؿ #�5�G�Y�{�5Ϗ��� z�ůׯ���)���� C�U�g�y���qϯ��� ���7��@��������2a,?�Q�c�u��	eߞ�2�������� ��
��.�@�R�d�k$ b.�������	�
��G] KK?�T_:Wd�f) 0]Ty���Д� 	����l�>��q�v��R�RX���>L1X���w�<'#�
����p��p�U(߆����l�@�ů����@lQ  �r�v�>�OR<�� GZ���oϑ�B�� /j/�/�/�/�/�/��p>�Doe&?��It$ ??$��>%�E
?q7A��q?�?�?=?O6� +��=��5.����5��$敕�5(4$��E�?�;;��.�3E>��H?E�5���OE8M�Y[E��=wE�HшO�;	�?�O�O�O�GO _"_4_F_X_j_��|W~|W  K� �p�h"p�U�U�� �Q��_�_oo�B0o�n����pM�u?333��R���!�D/  C��GÿP ?fff�> ����u�i�a�y؜_ fr�}����g�y�/m ���{����� pF@ �q�e� pDz�`4�����z2��� � �o%7��[e� '�9�������Ǐُ ���A����2�i� {�������ß՟�)� ׯ�h�A����{�� S���%�7�I�[�a� �@�R��v������� ��п����Ϙ�*�|� N�`�rτ���|��ߒ�0l�~ߐߚ��_��� ��*)�WD����S� L�#��b8 '��Зs� 4$�S&�)�ʠ� ��0�ԨюZ{���o'f����?�O�a�m�>�����m��� ������)�;�_� q�����e������ ��%��I�[�4� �������������� !3EW�{9/� ������/ A�jߜ�.?@?R?h5�2�|�?�?�?�?�=�/�22�?O0OBOTO fOxO�O�O�O�O�t�~ �N1,$WiWjL,���i �i�"�����/�yz_�_�_�_�V+$[0�W\_PnYr1gC�>��7o�-.�#��#De>�L�`ta�>R�)<#�
[;"pDo�R �8�/�VR���% !ce�b {e@ȡ|d �'�/����Zv��@���+B<!de` �����/���`�> q�d�_�_��YSI�t$ ��$�6>��b
{�͇AXT͏u������P+��̞;�.���G��Q$�敕W�(4$�xc��-�;��.���>��H���Q5{����8M�Y��]=t`ӕ�R�!�
�	���>�)�w�i� ~�������Ư5�M��>ا  �"$� �b�dor�`3��Z � �h?�Q�c�u�����z��R���c�?3�33e;�dGY{qD�/  C( G�P_ ?fffa>�a HT�'��_�(���� '�/]o��+������ ����Oi���=�[*|�F@ o�{��#r|�Dz���{�m�?�p�ʎ1n?`9 �K� ]�oρϓ�Y���߃� �����[�#�5�G� ]�k��[�m������� ������1�C���3E����W���9߯ ]�o߁ߓߥ߷߽Wb ��h��� ,�Pb���� ���*/��(?���/�/�/��Ȼ�0# �yꧠ/^>{oES�/�? �p�0�e�2�t q�v psUsyC*�?F' �`C41��4UN�e���8�$��9�L�O�H>����$�J+?=? O?a?s?�?�?p_�?�? �?�?O�_'O9OKO]O oO�OZo�O�O�o�O�O �O_3_�oG_Y_2}_ �_�_�_�_�_��_o o1oCo)goyoR��o��l�/�/������ą2@���	��-�>��V�2Q�z������� ԟ���
��#��=� h��t�����|���� �r����֯���1��t��L���ʩ(΁x�d�$q>l!���.�����>L��б��/�<#�	
�a�rp��?�|�>�s���$qcugq��W�xp׵@$شk" ��.��d�o������Vr'I�B�q����"߀C�U�8�yߋ�>{(�>�|���'���ߵ�Itk$ ��$H�>���	
��)�A��)���K�x���X�+��̗��.�����W�$�{����(4$ܿ�w��;��.��>���H��W�5�=��8M�Y�_��=а/�W� �@�f�	 ]�v�a����������������"1�$C�CSCH_GRP�16 2����S&� �\G�/J�  �� K� ��� (���o��Pȼ�@��S�	�s��u y�c%?333_��`�����D/  �C�pG�P ?fff_�>H���c%� ��o1�u"�-��_� z�)c�F/X/y/Ku3���`/�/�z�F@� �%�`��Dz �4��/�/z*�ʏ�� ����� /�?4/>? OO|/�/ �o�?�?�?�?�?�?O �O�O_BOTOfOxO�O �O�O�O_�_�_A__�\�T_�/,o�/�/�/ ?"?4?:o��o+o�o Ooaoso�o�o�oc�o �oqU'9K] �U5��k?E�W�i�s8�8_���s��g� ێ׿��,�%��Up��  b��O�L���g��\� ϥ���zy��w������g
T�Ҟ'� i�x��[��(�:�F�>���x�F�����̏ޏ�� ���8�J�\�n��� >�����ȟڟ���׿ "�4��X�j�|����� j�į֯������0� ^�T��x��������� ��������l�C�u���+�A�2�,t��H��������2�� ��	��-�?�Q�c�u� �����$�.�����0 0%�|]��t҉_oW �ߛ)Se����4��5G	K������>�q��b�R��>LfM��<��<#�
4�ҁp��U]߻����������<���T@�QU�r /��s� �Rq�3&|Z/�¤���B�=9/�/�/�/�/�/?�˥>�y�x�[?2It$ t?-$��>�z
T?�7A1�?N?�?r?�6� �+���E.��y� E�$敕0E�(4$�<E�?K;���.hE>��H�tE�5���E8'M�Y�E��=M�E�}ѽO�;	�?�O�O _WPOB_W_i_{_�_��_/���~�W  ���p��H"� e�U���Q�o*o<o�No�BeoSn����p<��u?333�b�� 	T!D/  C��G�P ?fff�>�!�u y�a 8Ϯ��_�r ���g ��/����Ű�B��4�UpF@ `H�Tq�e�UpDz�` i�TF���zg�G�9� �$6HZl 2����\�n���4� ���� �6�D�v�4� F�g�����ԟ��� 
��^�����v�0�������6�H�Z�l� ~�����0u���Aϫ� ��Ͽ��Ͽ�)�;� ��_ϱσϕϧϹ�߀���Ǐ�߳���ψȔ�����_)�Wy�7� T�߁�X��bm \� �����i$��&�L L)����e����Z@��.��\f�����?�/������>��� �Ԣ���(�:�L�^� p�I��������  ��$�6�H�Z�3~� ��i���������  2/Vhz�� �n/���
/ @R+?v�����c?u?�?�52�|�?�?�?$OM�//B2*OSO eOwO�O�O�O�O�O�O �O�t�~^A1a$�i�j �,ح�i�i�"�˧�/��y�_�_�_�_
f`$��0%g�_�Y�1Qg=C�>E�lo=c�X��#ye>L�`�a�sR�9<#�
�p"p�yobU��/fLR���<%@!�e0rQ �e@���dD�\?�ࢀ��vتu/" /";B q!�e���.��R�d�+p>Uq�d o�_����SIt$ Џ$�!F>��b
���A��T���$�Ώ��1`+����p�.����|�0a$敕��(�4$ܘ�P�b�;�{�.ĕ>��HЕ�0a5����8M�Y�8]=�`�0b�!�?�	6�O�:�s� ^�������ůׯ����j]���  �"Y�$r�d�rph� P�HZU�)xt�������P,�����LR�N��c<�?3338ep�9d||Y�qD/  C] �G�P ?fff8a>!q}T<�\�T�� 
8-���\�d]8o2�`� <����1�$%_���xrߐ*��F@ ��0���Xr��DzF��Ԁ�Ϣ�t�2��1�?�9 ܀ϒϤ϶��ώ� ���߸���4�FߐF� X�j�|�������� ������0�B�T�f��x���hz������ n���ߤ߶����� ����b��� +=Oa/��)/ �/��//_/��]?#��/?!?+�� ��90E#�y��/�>�o zS�/�?�(��p�90 (uB�t@q�v5p�U�y x*1O{'�`x491�D �N u��!H044�nx�L�O�H>���04 �J`?r?�?�?�?�?�? �_�?OO&OTO�_\O nO�O�O�O�O�o�O�O �o_"_4_F_h_"|_ �_g�_�_�_�_oo �0oBoTofoxo^�o �o���o$|�/-?��я���2N�,�>�P�b�s�R���2������ ӟ���	��-�?�Q� X�O�r����t���| 48�8�,�A'Q�S�@��J�A�f��t�@����������Yq>�!ȿc���E�յ>L��EϢd�O<#�
�a�rpտ�t���s������Yq�u�q���­p�@ YĠ"��c�+t<)@��4
�ϋr\~�B�q ����W�xߊ�m߮���s{]�>��1�\�R��^�It$ ,�$}�K>�2�
�^�A��^���*�<捰+�{����.�����ތ�$敕��(4�$�����;��=. �>��H,����5��<�8M�	YH���=�d���5�u���	��������� ���!3EW���l�D.i   8�� ��U� �]��� ����������(���� :Ø%?333�����ة��D/  C�pG�P ?fff��>}�٤�%���of� �S"�-������)�� Z/l/�/�uh��t/�/<�z F@  5!t�� Dz�!4/��/�/�*���� ��� //$/�?H/ R?O&O�/�/�o�?�? �?�?�?�?.O�O�O_ VOhOzO�O�O�O�O�O@_�_�_U_._�\�h_ �/@o�/ ??$?6?H? No�-o?o�ocouo�o �o�o�ow�o�o� i;M_q�i5��`?Y�k�}��8�L_ ���s�{1���֣ @�9�e�%�b���� `�!Ԝ�@֑����z ���w�Ԅ��{
h��\�}�������<�<N�Z�>�����Z� ��Ώ�����(�� L�^�p�����R���ʟ ܟ� ���6�H�!� l�~�����į~�د� ��� �2�D�r�h�&� ������¿Կ����
� ��.π�W����-�?�U�2�,�������	����2����/� A�S�e�w��������$ �.�����DD9ܐ] ���ҝ_�W�߯)g y����H���I[	_�	����>��q$��bb��1�>Lza��+��<'#�
H�(�p1�peq������@����P�	�h@�Q i�r/�߇ĘR��G& �Z-/�¸���B)�Q M/�/�/�/�/
??���>!���o?F�It$ �?$��>%��
h?�7AE�?�b?�?�?�6� +��=�(E.���4E��$敕DE(4$��PEOK;��.�|E>��H�E�5����E8M�Y�E��=a�E����O�;	�?_�O+_WdO V_k_}_�_�_�_"/��|�~�W  �� ���\"� ee 
 a�,o>oPobo�Byo�gn����u?333�(b�4	h!�D/  C�GÿP ?fff�> �5�uyqL����_ �r���g��/� ������V�*�H�ipF@ \�hq�e"ipDz�`}�hZ��,��z{�[�M� � 8J\n�F���� p�����H����"� 4�J�X���H�Z�{��� ğ֟�����0�r�  �2�����D��į&� ��J�\�n��������� D����UϿ�ѿ��� ����=�O���s��� �ϩϻ����Ņ�ۏ0�������Ȩ��� ��s)�W��K�h2�� ��l��b� p������ }$��&�``)0��� 3�y0����Z��B��pf�����?&/������>����Զ�� *�<�N�`�r��]�� ���������&�8� J�\�n�G����}�� ������ �4F/ j|�����/� �0/Tf?? ������w?�?�?�5�2��?�?OO+M
?CB2>OgOyO�O�O �O�O�O�O�O	_�� *^U1u$�i�j�,��i �i�"��ߧ	?��_�_o�_ft$�09g�_P�Y�1egQC!>Y���o=w�l��#�e>�L�`�a��R9<#�
��"p�o,bi�8�/+f`R��!P% T!�eDre �e@��d X�p?�����v��C"/6;B�!�e� �0�B�%�f�x�++p�>iq�do
oˏ�SI�t$ �$5F>��b
ď�A�T����8���E`+��̞��.�����Da$�敕��(4$�x��d�v�;��.ؕ�>��H�Da5{����8M�Y �L]=�`�Db�!-�S�	J�c�N���r������ǯٯ������$�CCSCH_GR�P17 2����@�&�� \4>��79  �"m�8rt �rp����\Z��=x�����Ϳ߿@����`R��b��cP�?333�Le��Md�Y�qD/ � Cq G�P ?fffLa>5q�TP� �ɉ��8b��p�x] Log�t�P�3�E�f�8%� _��Mߧߤ*��F�@ ����M�lr��Dz{������ߩ�g��1�?�9 ܵ����� ������!�+�����i� {ߤ{�������� �������/�A�S�e� w�����������.��A������ �����!�'�b �<N`r��P/ ��^/�B//&/8/ J/�/B�q?X�2?D?V?`��%n0z#�yT� 
?�>�o�S?O�]� �p�n0<u9B�tTq�v Ip�U�y�*fO�'�`�4 n1T�AD�Nu�VHe4�H��\'_3X>���e43Z�?�?�?�? �?�?O�_%O7OIO[O �O+o�O�O�O�O�O�O �o_!_�oE_W_i_{_ �_W�_�_��_�_o oKoAo�eowo�o�o �o��o�o��Y|0? b?���.�2��a��s�����������2 �������,�>�P� b�t����Ԅާ�ҁ�t ���im�m�a�v \����@�R��v����t!���"�4�8��
Γ�q>�!�����8�z�
�>LS�:�xz���<#�
!q�p
ϩ��J���ݢ���q�u�q)����pA�@�B��"�Ϙ� `tq^ �i
��r���B�*�&ߌ߭߿� �����ߨ{��>��f�𑿇�H��It$ Za�$��>�g�
A���A���;��_�q��°+����.�������$敕�(4$�)������;��.U�>��yHa���5��q�O8M�Y}�ɭ=:� ����j�����	���� ����=�/DVh�z���$CCS�CH_GRP18 2�����&� �\��v/��  m�� ��5Ғ� ٪��&8J\P��saݢ�� o��%?333ɵ"ʴ|�A�D/  C�p�G�P ?fffɱ>����%)!% ����"�-��ɿ��) �߰/�/�/�u��P/�/x$?!�c F@ V50b!���c Dz�w4�b/T?&?�*T�4�&� �2/D/V/h/z/@O �/�?jO|O�/�/!�? 
OO.ODORO�OB_T_ u_�O�O�O�O�O__�*_l_o,o�_�_>l� �_ ?�oD?V?h?z?�? �?�oo�oO�o�o �o�o�7I� m�������5���?����ӏ�8� �_��sL����E�A� �����fe�Z�jb� �Ŷ�V���u���9�9� *��-�R�*���
�� <���jӘ�����x������>���� ���$�6�H�Z�l�~� W�����Ɵ؟����  �2�D�V�h�Aό��� w�¯ԯ������.� @��d�v�����ȿ�� |������*��N� `�9���̭�ߏq�����2 <������%��=�28�a�s� �������������� 
4>$O�oԚ��� �]�����_�W�9@����n���@3��	��_K��>S�z�qbfb�Ӈ>L���ρ�O<#�
��~�p��&ce��%Z����J�NѦ>"_о@ a�R�j/����R��@�&�Z�/=��0�B� ��/	?*?<??`?r?%� >c!��?^�It$ �?$/�K>��
�?GA��O�?2O�?�6?+�{��~E.����E�>$敕�E(4�$ܦE^OpK;��=.�E>��H�E>�5���E8M�	Y�EF=�U>��'_MK	DO]_H_�_lW �O�_�_�_�_�_	ok��$CCSCH_�GRP19 2����:a?&� \.��>1�  ��g� 2"$�" �eeV
�a 7(�o�o�o�o:R�o�n�Z�\��J�?3�33F�bG�	�!D�/  Ck�G�P_ ?fffF>/! �J��y�q���\o� j�rFawn�J?-�?� `�2��G������pF@ Ӆ�qGuf"�pDzup��я��pa����� ܯ �������%�� ��c�u���u������� ��ϟ���ѯ�)�;� M�_�q�������鯗���(�����;���� ��ӏ���	��!Ϛ  ����6�H�Z�l�~� ��Jߴ���X���<��  �2�Dߎ�<�k�R�,�>�P�Z���h�t� �)Ng������ �Wr� �h�6%3��$ N!�&C ��)��`��� ���h�Nj;���%�fP�_�BO|/!->���_�-
��� ������������1� C�U���%�������� �����	�?Q cu�Q/���/� �E;�/_q ����/���?/�S,*�\��? OO(E2@}�[OmOO�O�M�?�B2�O�O�O__&_ 8_J_\_n_�_��~��^ �1�$yz<c�gygy [2p�V��?��:oLoyopo�f�$@�go.i(2A�g�C�!>���o��=��t3u>L�Mp4qt/�R�9<#�	
!�"p�b�D?�f�R���!�%�!#u�r� ;u@��<t�� ��?Z$k�X/�c� ��"�/�;B�!$u ����������ݏ+�p>��q`t�o�oB�cItk$ [�$�F>�ar	
;���Ad��5���xY�k��`+������.�����a$�{���(4$�#��۟�;��.O�>���H[��a5�=�k�8M�Yw��]�=4p���bd1��ʛ	 ��گů���7�)�>��P�b�t������$C�CSCH_GRP�1A 2������&� �\�>p߮9  g2�Яr�t/� �p����Z��x �2�@D�VϷ�m�[��R���yis��?333�e���di;�D/  �C� G�P ?fff�a>�qd���  �/�8ٿ�����]�o ����Ǐ�߼��߯%�_�J����:]�F@� P�\����r]�Dz ��q�\�N� ���NA.O I �,�>�P�b� t�:��ߢ�d�v����� /����(�>�L�~� <No����������  $f&�~8���>�P�b� t���r}�I/ �����/�/1/ C/�/g/�/�/�/�/�/ ?���?��?�?�?��Ȝ�0�#F�˷�? ?N;c�?�O`��T� d�0�u�BP��qo��p 3e3�$:�O'7Lp$D�1�˺�D6^�ud��H�4࿟��\�_�X>����4�ZOO0OBOTO fOxOQo�O�O�O�O _ �o__,_>_P_b_; �_�_q�_�_�_�_o �(o:o�^opo�o�o �o�ov��o�o $ 
�HZ3�~�|�?�?k�}�����2��؟�H������7�22� [�m��������ǯٯ �������I�i��� �ʉ������؂�� ���ٷ�ɿ����h���-Ǚ�����Y�E��>M1t��k`��>L�����<{��<#�
�qx��p�� �]���T����D�H���8�Y���@��L2d���t �����
}�7��*�By��ŝ��$�6��Z�l��	�>]����x���It$ ��-$)�>���
��
�A��
���,�����9��+���x�.��y���8�$敕���(4$ܠ�X�j�;���.��>��H���8�5����8'M�Y��@�=��8��!G�	>�WB {f���������$CCSC�H_GRP1B �2���4�&� \�(��/+�   �a0,�Ԭ�	Бy P�~1؝���4(��T��V0��D5?333@řAĄ����D/  Ce�G�P ?fff@�>)х�D5�)}!�� V�"d=l�@�['h9D� '?9?Z?,���/A?�?<��� F@ �5�!A%`�� Dzo �4�/��?�?[:ˑ���� ܩ/�/�/�/�/�O? O�O�O]?o?�oO�O �O�O�O�O�O�_�_�_ #_5_G_Y_k_}_�_�_@�_�o�o"o�_�l�5o �?�?�?�?�?OO ���o�0BT fx�D���R�� 6���,�>���6Ee�`LO&�8�J�TH�o b�n���H�����ς� ���eQ"���bb�0� -���H���=а��١� Z�������b�H5�����J�Y�<�v�	�<�'�>���Y�'� ��������џ���ο �+�=�O�}�υ��� ����ͯ߯������ 9�K�]�o���Kߥ��� ��ۿ����?�5��� Y�k�}Ϗϡχ����� ����M�$�V������"�2w<U�g�y�����	{��2��������  2DVhz�4 x>�����)*�]m a)a)U�joPgz�|94 Fsj�����(,������>�ʁ����b�bn���>LG .!n����<'#�
���p��p�e>������@����%�"��5%@�a 6$ɂ�/��T�ebR�6 ]j�/�҅ߧ�B��% ?�?�?�?�?�?�?��� >�!Z$�{<O�It$ UO$��>%�["
5O�GA�O�/O�OSOeF�+��=��E.���U��$敕U(4$��U�O�K;��.�IU>��HUU�5���eU8M�YqU�=. �U�^�_�K	�O�_�_�_�W1_�#o8oJo\ono�o�k��$CCSCH_G�RP1C 2�����a&� \��j���  a�ހ�" ~$)2� u�e�
�a�( ,>P�RgU~���Ӏc#��?33�3�r�51D/�  C��G�P /?fff�>�! ����qߏ��o|�� ���w��?����׏��ՑD�����W�F@ J�V��u�"W�Dz�pk�V�H��؊8H�(�� �&�8� J�\�n�4�����^�p� ڏ������"�8� F�x�6�H�i�����į ֯�����`�� ���x�2̸�����8� J�\�n�������"w� ��C߭Ͽ�������� ��+�=���a߳߅ߗ� �߻�ﳕ��ɟ�����јȖ�����@9 �g{�9�5/����Z� �rN0^���%��J4�! i6� --9���!�F  ����j��0�%^v������O�/���>�����
��*� <�N�`�r�K������ �����&8J \5/��k/��� ��/"4?Xj |���p?��� //?B/T/-Ox/�,@����eOwO�O�E2� �O�O�O_]�?1R2,_U_g_y_�_�_�_ �_�_�_�_����nCA c4�y�z�<ڽ�y�y�2 �ͷ�?���o�o�o�ovb4�@'w�o�i�ASw?S�!>G�n	Mpe�Z��3{u>L�p�q�/ub
I<#�
�!r2p{rWŻ?vNb���!>5B1�u2�S0�u@���tF�^� 	O�$��/��ںw�12?$KBs1�u�����@0��T�f�;�>W���t�o���cIt$� ҟ$#V>��r
���A�d���&�П��3p+���r�.����~�2q$�=���(4$ܚ�R��d�;��.ƥ>���Hҥ2q5����8M�Y�:m=@�p
�2r�1�A�	8� Q�<�u�`�������ǿ�ٿ�����$CC�SCH_GRP1�D 2����.�&� �\"N��%I  �2[�&��t��� ��s�Jjx�+��ϩϻϠ��.�����Nb�P�<�s>�?333:u���;t~i��D/  C�_0G�P ?fff:q>#�d>��w� �/HP���^�fm:U� b�>�!�3�T�&5o���;��:��F@ `����;�Z���Dzi� �������U��A�O�I ܣߵ������� ��������W�i�/ i�{������������ ��/ASew ��������/��/�������� ���/�r�/�/*/ </N/`/r/�/>?�/�/ L?�/0???&?8?�?�0�_OF� O2ODON��\@h3��B��?�N �|cO _�K�ˀ� \@*�'RǄB��7��e ���:T_�7�p�D\AB�@/T�^���DXSD6��p�lo!h>��� SD!j�O�O�O�O�O�O �O�o_%_7_I_w_ _�_�_�_�_�_��_ o�3oEoWoio�oE� �o�o���o�o�o9 /�Sew���� �����G�OPO�����2q�O�a�s�$����u���2��ү �����,�>�P�b� t�{�r������  �W[�[�O�dJt��v�.�@�m�dω�߄�����"�&��Ǽ�|�>�1�φ���h���>LA�(�h�򲞇�<#�
��p��ϗ��8���˲��|�����կ�Ѐ/�@|0��2�߆�N�_�L��W�߮����B ����z���������>��T��uϼ6��It$ O�$���>�U�
/���A�ā�)���M�_���+������.��������$敕(�4$�����;�{�.C>��HOޯ�5��_8M�Yk��=(Ї��X����	����� �+2DVhz���$CCSCH�_GRP1E 2�����&� \��|d?��  [� �0��x�#��%�Ǻ ���/&/8/J/�a/�O.˲��0]ӻ5?333��"����/��D/  C܀GÿP ?fff��> �����5�)�!���� v2�=㽷��'�9��? �?�?����>?�?O�Q0F@ DEP1�%��Q0Dz� eDP?BO�O�:B�"�� �  ?2?D?V?h?._�?�O X_j_�?�?��O�O
_ _2_@_r_0oBoco�_ �_�_�_�_�_ooZo �oro,|��oO �2ODOVOhOzO�O� �q�=����� ����%�7�ɏ[��� ����������Eܟ�O0�������HȐoِ �:�u�3�/����� }�Tu�"H�Xrِ�դ� D��c��'�'��ѯ �@��ّ���*��X&��Д���߀�����>���Д�� � �$�6�H�Z�l�Eϐ� ����Ư������� � 2�D�V�/�z���e߰� ¿Կ�����.�� R�d�vψ϶Ϭ�j��� ��������<�N�'� r��ܛ�͟_�q������2�<��������+2&Oas� �������4�> =�]�)�*}��m�) �)���o�g���9����&\���!'�P���M'9��>A��h/�_rTr��u%>�L� �!��o�<#�
��l�pu/"Qu8��&H����8� <�%,2M�%@�a�$ @�X?����b�ߋ6�jq?+����Bm�%�? �?O*OONO`O�� �>Q1�$���O�I�t$ �O$>��"
�O�GA��O�O� _�O�F- +��̞lU.���xU,!$�敕�U(4$�x�UL_^[;��.�U�>��H�U,!5{���U8M�Y�U4=� e,"��o;[	2_Ko6oooZg�_�o��o�o�o�o�o{�$�CCSCH_GR�P1F 2����(q&�� \���  ��U� 2�$ �2� �umuDrq%8�����(b��~H��J��#8�?333�4%�r5$x�1D/ � CY�G�P ?fff4!>1y8� y�q����J�X�` 4/O�\�8O�-�N� ����5�����΀F�@ ��́5�T2΀Dzc��͏����O������� ܝ����� ӏ叫�	��կ�Q� c���c�u��������� ﯭ�����)�;�M� _�q�����׿�ϗ��￩̸)ϋ�߯��� ӟ���	�߈"�� � ��$�6�H�Z�l�~�8� �ߴ�F���*���� � 2�|�*�Y�@��,�>�H���V�b�9<w ����/v�����E� �0��V�$5!�4<1�6 10��9��N�� �� V�<z)��%�v>M��0_j?�>���M�}������� �������1C q/y����� �/�	�/-?Qc �??���?��� /3/)/�?M/_/q/�/ �/{?�/�/�O�/A<� J��O�O _U2k�I_�[_m__�]oO�R2 �_�_�_�_oo&o8o Jo\onou�l��n�A�4 ���<Q�U�U�IB^� D�nOp�(:g^�v�4	P�w
y Q�w
�Sv1>����M��8��bC�u>L;�"�xb?�b�I<#�
	1�2p��r��2O�v�b��v1�5�1����0)�@v�*���Տ�O H4Y�F?�Q�2y?�KB�1��t����� ��˟ݟ�;z�>΁N��yo0�sIt$ ZI�$�V>�O�
)�{�At{�#���G�Y�ުp+����.�������q$敕�(4$��ɯ۫�;��.=�>��yHI��q5��Y�O8M�Ye��m="� ���rRA����	��ȿ ���׷%��,�>�P��b�tσ��$CCS�CH_GRP1G 2������&� �\�N^�I  UB����r��z�� ���j����� �2�D�P��[�I��b���W���?333�u
Ҳt|�i)�D/  C�0�G�P ?fff�q>���d������? �H��p����m����� �������5�o8��x�	JK�F@ >�0J��тK�Dz��_�J�<����<Q_Y ��,�>�P�b�( ���Rd����	?�� ��,:l*< ]������ �T//�l&,� ��~/,�>�P�b�t� ���/�k/}/7?�/�/ �/�/�/�/�??1?�? U?�?y?�?�?�?�?����O���O�O�O��� ��@�34���oO-^)� �c~Ow_N%��B�R"�@ ���R>���]���!u!� J�_G:�T�A�ʦT $ny�RֻX�D���xzl�o�h>����D �j�O__0_B_T_f_ ?�_�_�_�_�_��_ oo,o>oPo)�to�o _��o�o�o�o�� (�L^p��� d���� ����6� H�!�l����O�OY�k�}���2��Ưد�����%�2 �I�[� m��������ǿٿ� �����7�W��ق�w� �����ƒ�����@�Ϸ����� �V���@ׇϙɝ�G�3��>;Ab���Y"N"ߓo�>L�П�ߏi���O<#�
��f�po���K%���B�����2�6���&�G���@ ���:BR���ń�Ï@���k�%����Bg� �Ջ����$��H�Z����>K������ϭ�^��It$ ��$�K>���
����A�����������'�+�{��f.���r�&�$敕�(4�$܎FX;��=.�>��H�&��5���8M�	Y�.�=���&�ϑ5	,E0iT ������� +��$CCSCH_�GRP1H 2����"!?&� \��?>�  ҒO@ ��Ԛ���%g%>�l! �/�/�/�/"�/�.�B��D@��2E?3�33.Շ"/�rɦ�D�/  CS�G�P_ ?fff.�>� s�2Es9k1�� �D/�2 RMZ�.�I7VI2�O'O HO�ϵ?/O�O���0F@ �E�1/5N��0Dz]0�D�?�O�OpIJ������ ܗ? �?�?�?�?�_O_�_ �_KO]O��]_o_�_�_ �_�_�_�o�o�oo#o 5oGoYoko}o�o�o��o�|�#�O� �O�O�O�O�O_	��� �����0�B�T�f� x�2�����@�ҏ$��� ��,�v�$US�:_�&�8�BX�P�\� ��6'쟪���p����� �u?2���rP����� 6���+��Ş鏚H��� �Џ�P�6*#������&8�G�*d���	��>���G��w��� ������ѯ㯼��� +�=�k��s������� ��Ϳ������'�9� K�]��9�ϥ�~��� ������-�#���G�Y� k�}ߏ�u���ߞ��߀;��D�������2@eLCUgy�i��2�����  2DVhoDfN� �����)�*��K}O9O9 C�X>wh�jI"/4/a/X/}&�� �'/)(�'�p�>���/�z��r�r\��%>L�501\��{�<#�	
���p�/�"�u,��&���p���5�2��#5@pq$4�� �?z�B�Sr@�FKz�?��s��B��5OnO��O�O�O�O�O��t0>��1H4s/i/*_#Itk$ C_$�>�I2	
#_uWA $u__�_xA_SV� +����U�.����U�!$�{���U(4$�e��_�[;��.7e>���HCe�!5�=�Se8M�Y_e��=0{e�"L�o�[	 �_�o�o�o�go&�8J\n}{�$C�CSCH_GRP�1I 2�����q&� �\��X���  O�̐�2l4B t0�u�u��q�8��@,�>��bU�C�����yQ3��?333�%���$�#AD/  �C��G�P ?fff�!>�1����� ��}��j�ϝ��/ Ƈә�O����ş���2�����E�F@� 8�D����2E�Dz ڀY�D�6��ƚ6	 ��&�8�J� \�"�����L�^�ȟڟ �گ����&�4�f� $�6�Wώ�����Ŀֿ ����N���ߍ�f� ܸ���x�&�8�J� \�n������"e�w�1� �߭߿������߯�� +��O��s���� �������������Ȅ�����.I�wi� '#?�x�qHռ�<@ L���5�8D�1WF�0 %I���40��z�s5L�����_�?t��>��������*< N`9/����� �/�&8J#? n�Y?����� �?/"/�?F/X/j/|/ �/�/^O�/�/�/�/? �?0?B?_f?�<����S_e_w_�U2��_�_H�_�_m�Ob2o CoUogoyo�o�o�o�o �o�o��~1QQD|� |�qL��̉̉�B�ϻ� �O癟����vPD�P���y�QA�-c�1>5�\��MS�H��Ci�>L�����?<cr�I<#�
�1`B�pi��EթO�<r���1,E0A�� �A@��@����4�L��O�4 �½?���e�B�?[BaA��������B�T�K�>E�ń�x���~sIt$ ��-$f>�Ƃ
���A}t򯚯���Ц!��+���`�.��y�l� �$敕|��(4$܈�@�R�;���.��>��H��� �5��е8'M�Yܵ(}=���� ��A	�/�	&�?�*� c�Nǜ��ϣϵ�����������$CCSC�H_GRP1J �2�����&� \�^��Y   �BI��鄔��y�a� 8zf���ߗߩ߻��(����<r�>�΃,�?333(���)�ly���D/  CM@G�P ?fff(�>�mt,�m�e�?�H >���L�T}(�C�P�,� �!�B�E�o��)���<�J��F@ ����)�H���DzW����������C��Q�_�Y ܑ��������� ��E�W��?Wi {������� /ASew�@�y/�/
/��,�/ ��/������������ ?|��/�/�??*?<? N?`?r?,O�?�?:O�? O�?OO&OpOM_`4_ _2_<�/ JPVC��0��O�^��js �O�_�%9⹐�"JP� b��0�Ԗ%��u���J Bo�G���TJQ0�d�n����2hAT$�^��l<x>���ATz q_�_�_�_�_�_�_� oo%o7oeo�moo �o�o�o�o���o�o֏ !3EWy3��� x�����'��۟ A�S�e�w���o����� ���5�_>_Я���
�2_�=�O�a�s���	c���2����ҿ� ����,�>�P�b�i� `��ή�Δ�����E- I�I�=�R/8'b�d�� .�[�R�w�͔���נ�����ת�j�>��A��t��"�"V����>L/��V���u�<'#�
��ݒp�߅�p�%&��ֹ���j�@�����⾐�@j! �B��t�<�M":��� E*�m���Bޑ� �h�����~�������n�>��B�m�c�$�ïIt$ =$��>%�C�
oA��o��;M��+��=��.�������$敕�(4$����;��.�1>��H=��5���M8M�YY��=�u��F���	������/ /2/D/V/h/w+��$CCSCH_G�RP1K 2�����!&� \��RO��  I��@�� f��n��%�%���!�� ??&?8?�O?=>�����@K�E?33�3���"�����D/�  CʐG�P /?fff��>���� �E�9�1�w��/dB�M �ͥ��7�I���O�O�O���y�,O�O _��?@F@ 2U>A�5��?@Dz�0ST>O0__�J80��� �O O 2ODOVOozO�_FoXo �O�O���_�_�_
o o .o`o0Q�o�o�o �o�o�o�oH���`����Or� _ 2_D_V_h_z_����_� q�+�������ˏݏ� ���%���I���m�� ����ퟛUʯ�_�������X�~Ǡӓ(� �'c�!����r�k�B� �26�F�Ǡ�咲2��� Q��������	�.� �ǡ�*���m�F6��������ǹό�>�������� �� $�6�H�Z�3�~����� ��⿄����� �2� D��h�z�S�ϰ��� ���ϰ�
����@�R� d�vߤߚ�X������� �����*�<�`��@����M_q�2�L ������2=Oas�� �����D�N .+ K�v9v:k��}�9�9�� ��w���I�/�/�/�/�&J�z 7{/�)�;7'��>/�V?��pM�B���c5>L�0�1��]"��<#�
z�Z�pc?2?���66"����&�*�5B;�5@�q�4.�FO �����r��yF�z_O���B[�5O�O_@_�O<_N_��0>?A�4�/�/�_x#It$� �_$>��2
�_�WAw$�_�_o�_��V0+���Ze.����fe1$�=�ve(4$܂e:o�Lk;��.�e>���H�e15����e8M�Y�e"-=@�0�e2��)k	 o 9$]Hw�o��� ���$[