��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA!R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B!SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sA�TB�d�5�MO<� �cE D [�M�c��^qREV��BILrw!XI�� QrR  �� OD�P�q$NO^PM�Wp�t�r/"�w� �u��q�r�0D`S �p E RD_E��pCq$FSSB�n&$CHKBD_[SE^eAG G�"$SLOT_�H�2=�� V�d�%�x�3 a_EDIm   � �"���PS�`(4%$�EP�1�1$OP��0�2�a�p_OKv�UST1P_C� ुd��U �PLACI4!�Q�4�( ra�COMM� ,0$D����0�`��EOWB�n�IGALLOW�� (K�"(2�0VARa��@�2a�o�L�0OUy� !,Kvay��PS�`�0�M_O]����CCFS_UT~p0 "�1�3�#�ؗ�`X"�}R0  4�F IMCM�`O#S@�`��upi �_�pB�B}�a���M/� h�pIMPEE_F�N��N��0�@O��r�D_�~��n�Dy�F� dCCq_�r0  T� '��'�DI�n0"���p�P�$�I������F�t X� GRP0��=M=qNFLI�7��0UIRE��$g"~� SWITCH5��AX_N�PSs"C�F_LIM�� � �0EED���!��qP�t�`PJz_dVЦMODEh��.Z`�PӺ�ELBOF� ������p@� ���3���� FB�/��0�>�G�� �� WARNM��`/��qP��n�N�ST� COR-�0bFLTRh�TR�AT�PT1�� $ACC1a��N ��r$ORI�o"V��RT�P_S� C�HG�0I��rT(2��1�I��T�I1���� x pi#�Q��HDRBQJ; CQ�2L�3L�U4L�5L�6L�7L֤ N�9F3��O`S <F +�=�O��#�92��LLECy�>"MULTI�b�"�N��1�!���0T�� ;�STY�"�R`�=l�)2`����*�`T  |� �&$��۱m��P�̱�U�TO���E��EX�T����ÁB���"�2� (䈴![0�������<�b+�� "D"���ŽQ��<�$��kcl�9�#��與1��ÂM�ԽP��"� '�3�$ L@� E���P<��`A�$JOBn�T���l��TRIG3�% d K�������<���\��4+�Y���_M��o& t�pFLܐ�BNG AgTBA � ���M��
�!��p � �q��0�P[`�,�O�'[���0t�na*���"J��_R���CDJ��IdJk�D�%C�`�Z���0��P_�P��@ 7( @F RO.��&��t�IT�c�NOAM�
����Sp�P`T)w@���Z�1P�d���RA�0��p2b"����
$T��.��MD3�T��`QU31���p(5!HGb��T1�*E�7��c�KAb�WAb�cA4#Y�NT���PDBG�D�� *(��PU�t@X��W���AX���a��eTAI^cB�UF��0!+ g� 7n�PIW��*5 P�7M�8M�9
0�6F�7SIMsQS@>KEE�3PATn�^�a" 2`#��"�L64FIX!, ���!d��D�12Bus=CCI�:FgPCH�P:BAD렀aHCEhAOGhA]HW�_�0>�0_h@�f�Ak� ��F�q\'M`#�"�:DE3�- l�p3G@��@FSOES]FgH�BSU�IBS9WC��.� ` ��MARqG쀳��FACLp�SLEWxQ�e�ӿ��MC��/�\pSM_JB M����QYC	g�e���Д0 ā�C�HN-�MP�$G� Jg�_� #���1_FP$�!TC uf!õ#�����d�#a���V&��r�a;�fJ�R���rSEGFR�PIO� STReT��N��cPV5���!41�r��
r>�İ�b�B�O�2` +�[���,qE` &�,q`y�Ԣ}t��yaSIZ%���t�v�T�s� �z�y,qRSINF}Oбc���k ��`��`�`L�ĸ �T`7�CRCf�ԣCC/�9��`a�uah�ub'�MIN��uaDs�T#�G�D�YC��C������e�q0��� �E�V�q�F�_�eF��N3�s�ah��Xa+ep,5!�#1�!OVSCA?� A��rs1�"!3 ��` F/k��_�U��g��]��PC�� a�s���R�4� ����N�����5a�R�HANC��$LG��P�f1�$+@NDP�t�AR5@N^��a�q���c��ME�18���}0��3RAө�AZ �t���%O��FCTKѐ�s`"�S�PFADIJ�OJ�ʠ�ʠ����<���Ր��G8I�p�BMP�d�p8�Dba��AES�@	�vK�W_��BAS��| �G�5  M�=I�T�CSX[@@��!62�	$X�R��T9�{sC��N�`��a~P_HEIGH�s1;�WID�0�aV�T ACϰ�1Ap�Pl�<���EXPg�܈�|��CU�0MM�ENU��7�TI-T,AE�%)�ap2��a��8 P� �a�ED�E�Н�P;DT��REM.���AUTH_KEY#  ������ �b��O	���}1ERR9LH� �9 \� �q�-�OR�DB�_IDx�@l �PUN_O��>Y�$SYS0��4�g�-�I�E�EVx�#��(�PXWO��z �: $SK7!�f2�(�Td�TRLn��; �'AC�`ܱ�ĠIND9DJ$.D��_��f1��f����PL�A�RWA�j���SD�A��!�+r|��UMMY9d�F�10d�&���J��<��}1PR� �
3�POS��J�=� �$V)$�q�PL~�>���S�ܠK�?����CJ�@\����ENE�@T���A���S_�REC�OR��BH z5 O�@=$LA�>$~�r2�R��`�q��b`�_Du��0RO�@�aT[�Q��b�������! }У�PAU�S���dETURN,��MRU�  ;CRp�EWM�b�A�GNAL:s2$L�A�!?$P�X�@$P�y A �Ax�C0 #ܠDO�`X�k�W�v�q�GO_AWAY��MO�ae���]�C�SS_CCSCB� C �'N��CERI��гJ`u�QA�0�}��@�GAG� R�0�`��0{`��{`OF�q��5��#MA��X���.a�LL�D� �$���sU��D)E%!`���OVgR10W�,�OR|�~'�$ESC_$`>�eDSBIOQ���l ��B�VIB&� �c,�����f��=pSSW���f!V�L��PL���AR'MLO
��`�����d7%SC �bALspH�MPCh �C�h �#h �#h 5�UU ���C�'�C�'�#�$'�d�#C\4�$�pH���Ou��!Y��!�SB���`k$4�C��P3Wұ46$VOLT37$$`�*��^1��$`O1*�Y$o��0RQY��2�b4�0DH_THE�����0SЯ4�7AL�PH�4�`���7�@ ��0�qb7�rR�5 �88� ×���"���Fn�MӁVHBPFUAFLQ"D�s:�`�THR��i2�dB�����G(��PV@P�����������1�J�2�B�E�C�E�CPS u�Y@��Fb3���H� (V�H:U�G�
X0��FkQw�[�Na�'B���C� INHBcFILT���$��W�2 �T1�[ ��$����H YАAF�sDO��Y�Rp� fg�Q �+�c5h�Q�iSh��QPL���Wqi�QTMOU�#c�i�Q\Ѐ�X�gmb��vi�h�bA4i�fI�aHIG��c�a	xO��ܰ��W��"vAN-u!��	#A�V�H!Pa8$PP�ד#p�R_:�A�a��B�N0�X�MCN���f1[1�q�VE�p��Z2;&f�I@�QO�u�rx�wGld�DN{G|d��aF�>!�9��aM:�U�FWA�:�Ml���X� Lu��$!����!l�ZAO����0%O�lF�sL�13�DI�W�@���Q���_��!C�URVA԰0rCR41ͰZ�C<�r�H�v����<�`��<�(�f�CH�QR3�S���t���Xp�VS_�`�ד��F��ژ�����NSTCY?_ E L����A1�t�1��U��24�2B�NI O7�����އDEVI|� �F��$5�RBT.xSPIB�P���#BYX����T���HNDG��G HC tn���L�@�Q�C���5��Lo0� H��閻�FBP�{tFE{�5�t�h�T��I�DO���uPMCS�v>�f�>�t�"HOTSWt�`s�?ELE��J T���e�2��2d5�� O� ��HA7�E��344�0?��A�wK �� MDL�/ 2J~PE��	A���s��tːÈ�s�J ÆG!��rD"�ó���L��\�TO��W�	���/��SLAV�wL  \0INPڐp���`%ن_CFd�M� $��ENU��OG��b�ϑ]զP�0`ҕ�]�IDMA�Sa��\��WR�#��"]�VE\�$a�SKI�STs�H�sk$��2u���J�À�����	��Q���_�SVh�EXCLU8MqJ2M!ONL��D�Y��|�PE ղI�_V�APPLYZP��HID-@Y�r��_M�2��VRF�Y�0��r�1�cIO#C_f�� 1����2��O��u�LS���R�$DUMMY3ҏ!���S� L_TP/Bv�"���AӞ�>ّ N ����RT_u�� ��G&r[�O D���P_BA�`��3x�!F ��_5���H��>��� ��� P $�KwA�RGI��� q�2wO ��SGNZ��Q �~P/�/PIG!Ns�l�$�^ sQ�ANNUN��@�T<�U/�ߴ�L�Azp]	Z�d~��EFwPI�@ �R @�F?IT~�	$TOTA%Š�d���!�M6�NIY�S+����E�A[�
DAYS\�ADx�@���	� �EFF_A�XI?�TI��0zC�OJA �ADJ__RTRQ��Up�!�<P�1D �r5̀Ll�T�p? ]P��"p��mtpd��V 0w�G������-��SK�SU� ���CTRL_CA��� W�TRA�NS�6PIDLE_PW���!��A��V��V_�l�V ?�DIAGS���X� /$2�_;SE�#TAC����t!�!0z*@��RRD��vPA���p ; SW�!�!�  ��o2l�U��oOH��3PP� ��IR�r���BRK'#��"A_A k���x 2x�9ϐZs2��%l�W�pt*��x%RQDW�%MS�x�t5AX�'�"��L?IFECAL���10��N�1{"�5Z��3{"dp5�ZU`}�M�OTN°Y$@FsLA�cZOVC@p��5HE	��SUPCPOQ�ݑAq� Lj �(C�1_X6�IEY
RJZRJWRJ�0TH�!�UC��6�XZ_ARl�p��Y2�HCOQ��Sf6AN��w$���ICTE�Y `>��CACHE�Cp9�M�PLAN��oUFFIQ@�� �0<�1	��6��wMSW�EZ 8䐟KEYIM�p��TM~�SwQq�wQ#�|��TROCVIE� ��[ A�BGLx��/�}�?� 	��?��D\p�ذST��!�R� �T� �T�� �T	��PEMAI�f�ҁ��_FAKUL�]�Rц�1��U�КR�DTR�E�^< �$Rc�uS�% IT��BUFW}�W��9N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTT(����sP��M��Ot�T�LwAX � ��XX~`9#�c_G�3
ЧYN_1�_�D���1 �2M�*��T�F��H@ ~g�`� 0p���Gb-sC_R�AIAK���r�t�RoQ8�u7h�qDSPq��rP��A�IM�c6�\����s2�U�@�A�s�M*`IP���s�!DҐ6�TH�@n�)�OyT�!6�HSDI3��ABSC���@ V`y��� �_D�/CONVI�G��H�@3�~`F�!�pd��psqSCZ"���sgMERk��qFB��Lk��pET���aeR�FU:@DUr`����x�CD,���@p;cJHR�A!��bp�ՔՔ+PSԕCJ���C��p��ғSp�cH *�LX�:cd�Rqa�|  ����W��U��U���U�	�U�OQU�7R�8BR�9R��0T�^�1k�U1x�1��1��1��U1��1��1ƪ2Ԫ�2^�k�2x�2��2���2��2��2��2*ƪ3Ԫ3^�3k�x��3���o���3��3ʹ�3ƪ4Ԣ�AEX9Tk!0�d <� 7h �p�6�pO��p����Na�FDRZ$eT^`V�Gr����䂴2�REM� Fj��BO�VM��A�TR�OV�DT�`-�MX<�IN��0,�W!'INDKЗ
w�׀�p$DG~q36���P�5�!D�6�RI�V���2�BGEAR��IO�%K�¾DN �p��J�82�PB@�CZ_MCM�@�1��r@U��1�f ,��a? ���P��.�"?I�E��Q�!���`m���g� _05Pfqg RI9ej��k!UP2_ h � �cTD�p����! a�����BAC�ri T�P�b�`Z�) OG��%�8��p��IFI�!�p0m�>��	�PT�"]��FMR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4�@��Uk��� �T�FS#p�Tl �P���e�qP�p$GEX_���1M�2��2� 3�5��9G ���m ��Ѝ��SW�eOe6DEBcUG���%GR���pU�#BKU_�O�1'� �@PO��I5�5MSf��OOfswSM���E�b�@�0�0_E� n �0 Y4 �TERM��o�5 �ORI�+�p�FF �GSM_���b�q�.���TA�r�Cp��UP�Rs� 9-�1�2n$�' �o$SEG,*> E�LTO��$US]E�pNFIAU"�4�e1���#$p$UFR���0ؐO!�0��f��OT�'�TAƀ�U�#NST�PA�T��P�"PTHJ�����E�P rF�V"ART�``%B`�abU!�REL:�aSHF�T��V!�!�(_SH"+@M$���� ��@rN8r����OVRq�N�rSHI%0��UN�= �aAYLO�����qIl����!�@��@ERV]��1�?:�� �'�2��%��5�%��RCq��EASYM�q�EV!WJi'��}�AE���!I�2��U@D@��q�%Ba��
5Po�X�0�p6OR�MY�& `GR��t2b5�n� � ��UPa�Uu� Ԭ")���TO�CO!S�1POP@ ��`�pC�������YOѥ`REPR3�b�aO�P�b�"eP�R�%WU.X1��e$7PWR��IMIU�2sR_	S�$VIS���#(AUD���Dv" ;v��$H���P__ADDR��H�AG�"�Q�Q�QБR~p\Dp1�w H� SZ� a��e�ex�e��cSE��r��HS���MNvx ����%Ŕ��OL����p<P��-��AC�ROlP_!QND_�C��ג�1�T �RO�UPT��B_�VpQ�A1Q�v��c_��i ���i��hx��i���il��v�ACk�IOU���D�gfsu^d�gy $|�P_D��xVB`bPRM_�b{U�ATTP_א�Haz (��OBcJEr��P��$���LE�#�s`{ � ��u�AB_�x�T~�S�@�D�BGLV��KRL~�YHITCOU�[BGY LO a�TEM��e�>�+P'��,PSS|�P�JQUERY_FLA�bG�HW��\!a|`�u@�PU�b�PIO��"�]�ӂ/dԁ=d�ԁ�� �IOLN���}����CXa�$SLZ�$INoPUT_g�$IPb#�P��'���SLvpa~��!�\�W�C-��B$�IO�pF_AuSv��$L ��w �F1G�U�B0m!a���0HY���ڑ�����UOPs� `������[� ʔ[�і"�[PP�SIP��<�іI�2�x��P�_MEMB��i`� X��IP�P�b{�C_N�`����R0�����bSP��p�$FOCUSBG�a~�UJ�Ƃ �q  � o7JOG�'n�DIS[�J7�cVx�J8�7� Im!|�)�7_LAB�!��@�A��APHI�b�Q�]�D� J�7J\���� _KE}Yt� �KՀ�LMONa����$XR��ɀ��WATCH_��3���EL��}Sy~���s� �Ю!V�g� �CTR3򲓥��LG�D� �R��I�~
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�Gȴ I�F�%SO���q �Ɩ�@��v��ƴ��K�S�����w�k�N����E��\���'�"*�U�s5��@L>�4�7DAUZ�EA�pՀX�Dp�f�GH�B��OGBOO��g� C���PIT����� ��REC��S'CRN����D_p�aMARGf�`��@:���T�L���S�s¡�W�Ԣ�Iԭ�JG=MO�MNCH�c���FN��R�Kx�PR�Gv�UF��p0��F�WD��HL��STP��V��+���Є�RS��H�@�몖C�r4��?B��� +�O�U �q��*�a28����Gh�0PO������b��M8�Ģ��EX���TUIv�I��(� 4�@�t�x�J0@J�~�P��J0��N�a��#ANA��O"�0V�AIA��dCLEA�R�6DCS_HIP"�/c�O�O��SI��S��I�GN_�vpq�uᛀTܓd� DEV-�LL�A �°BUW`�j�x0T<$U�#EM��Ł����0�A�R��x0�σ\�a�@OS1�2��3�a�`� �ࠜh�AN%-���-��IDX�DP�2MRO���Գ!�ST��R�q�Y{b! �$E&C+��p.&�A&���`� L ��ȟ%Pݘ��T\Q�U�E�`�Ua��_ � �@(��`������# �MB_PN�@ R`r��R�w�TR�IN��P��BAS8S�a	6IRQ6��{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?��?RIAt,1ID`�D�� d1��RQQp�rpDSTB
`� 1�F�HAXD2��|�G�LEXCES?R��q�BMhPa�͠D�BD4 �E�q`�`�F_A�J�C[�Ot�H� K��� \��d�bTf$� ��LI�q��SREQUIRE��#MO�\�a�XDESBU��,1L� M�� �p���P�c��AA,1N��
Q�q�0/�&���-cDC��B�sIN�a?�RSM��Gh� N#B��N�iP�ST9� � 4n��LOC�RI��v�EX�fANG���A,1ODAQ䵗ƞ@$��9�ZMF �����f��"��%u�#ЖVSUP�%`F�X�@IGGo�� �rq�"��1��#B��$���p%#by��rx����vbPDATA�K�pE;����R��M܋�*� t�`MD
�qI��)�v� �t�A��wH�`��tDIA<E��sANSW��t(h���uD��)�bԣ�(@$`� PCU�_�V6�ʠ�d�PLODr�$`�R���B����B�p�����,1R�R2�E�  ���V�A/A d$OCALI�@��G~��2��!V��<$R�SW0^D"���ABC�hD_J2�SE�Q�@�q_J3:M�
G�1SP�,��@PG�n�3m�u�3p
�@��JkC���2'A�O)IMk@{BCS�KP^:ܔ9�wܔJy�{BQܜ������`_AZ.B��?�E�L��YAOCMP0�c|A)��RT�j�ƚ�1�ﰈ��@1�茨����Z��SMG0��pԕ� ER!��m��INҠACk��p����b�n _�������D�/R͠�DIU��CDH��@
�#a�q$V��Fc�$x�$@���`@���b��̂��E�H �$B�ELP����!ACC�EL���kA°IORC_R�p�@�yT!�$PS�@
B2L$P���W3��ط9� ٶPATH��.�γ.�3���p�A�_��_�e�-B�`C����_MG�$�DD��ٰ��$FW�@�p����γ�����DE��PPABN��ROTSPEE�u��O0��DE�F>Q��$P$USSE_��JPQPC��JY����-A 6qYN�@A�L�̐�L�7MOU�NG��|�sOL�y�INCU���a�¢ĻB��ӑ�AENCS���q�B����,�D�IN�I�����pzC�VE����ҏ23_U ��b�LOWL���:�O0��0�Di�B�PҠ� ���PRC����MOS�� gTMOpp�@-GP�ERCH  M�OVӤ �����!3� yD!e�]�6�<�� ʓ	A����LIʓdWɗ���:p3�.�I�TRKӥ�AY����?Q^� ��m�b��`p�CQ�� MOM�B?R�0u��D���y�0Â���DUҐZ�S_BC?KLSH_C���� o�n��TӀ���
<c��CLALJ��pA��/PKCHKO0:�Su�RTY� �q!��M�1�q_
#c�'_UMCP�	C����SCL���LMTj�_L�0X����E�� �� ����m�h���6��PC�����H� �P�ŞC�N@�"XT����CN�_��N^C�kCSF����V6����ϡj����nCAT�SHs�����ָ1����`����������PA�&��_P���_P0� �e���O1u�$xJG0� P{#�OG���TORQU(�p�a�~����Ry������"_W��^�����4t�
5Tz�
5I;I ;Iz��F�`�!��_8�1��VEC��0�D�B�21�>p	P�?�B�5JRK�<��2�6i�DBL_S�M�Q&BMD`_DLt�&BGRV4
Dt�
Dz��1H_���31��8JCOSEKr�EHLN�0hK�5oDt�jI��@jI<1�J�LZ1�5Zc@�y��1MYqA�HQBT�HWMYTHET09�NK23z�/Rn��r@CB4VCBn�CqPASfaYR<4gQt��gQ4VSBt��R?UGTS���Cq��a���P#���Z�C$DU u ��R䂥э2�Vӑr��Q�r�f$NE�B+pIs@�|� �$R�#QA'UPeYg7EBHBA�LPHEE.b�.bS �E�c�E�c�E.b�F�c(�j�FR�VrhVghd���lV�jV�kV�kV��kV�kV�kV�iH�rh�f�r�m!�x�kH��kH�kH�kH�kH*�iOclOrhO��nUO�jO�kO�kO�kUO�kO�kO�FF.b�TQ���E��egSPB?ALANCE��R�LE�PH_'USP�衅F��F��FPFULC�3��3��E���1�l�UTO_<p �%T1T2t���2NW�����ǡ��5�`�擳�T�O�U���� INSEG��R�REV��R���gDIFH��1���6F�1�;�OB��;�C��2� �b�4L�CHWAR��i�A�BW!��$MEC�H]Q�@k�q��AX�k�P��IgU�i��� 
���!����RO�B��CR��ͥ�� �C��_s"T� � x $�WEIGHh�9��$cc�� Ih�.�I9F ќ�LAGK�8qSK��K�BIL?�cOD��U��STŰ�P�; �����
�����
�Ы�L���  2�`�"�DEKBU.�L&�n��POMMY9��NA#�δ9�$D&����$��� Q  _ �DO_�A��� <	���~��LђBX�P�N��+�_�7�L�t�OH  �/� %��T�����T�����TICYK/�C�T1��%�Ä����N��c�Ã�R� L�S���S�����P�ROMPh�E� $IR� X�~ 8���!�MAI�0��4j���_9����tt�l�R�0COD��sFU`�+�ID_" �=�����G_SU;FF<0 3�O����DO��ِ�� R��Ǔن�S����!{�������	�H)�_F�I��9��ORDfX� ����36h��X�����GR9�\S��ZDTD���|v�ŧ4 *�L_NA4���K��DEF_I[�K��� g��_���i��Ɠ������IS`i �萈�����e����4�0i�Dg�����D� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{ԓ� {ԡ�{����}��v� �Ա��g������^� ��K�Փ����!w�N�P'���^���,`b�W\�[R�	7�sTEFĨ �OULOMB_u��0�VISPI�TY�A�!OY�A�_FRId��(�SI���R�����R�3���W�W���0��0_,�EAS%��!�& "����4p�G;� h� ��7ƵCOEFF_Om���m��/�G!%�S.�߲CaA5����u�GR`� � � $hR� �X]�TME��$R�s�Z�/,)�ER��T;�:䗰�  �]�LL��S�_3SV�($~��q��@���� "�SETU��MEA���Z�x0�u������� � � �� ȰID�"���!*��&"P���*�F�'��A��)3��#����"�5;`*��RE�C���!7�SK_���� P	�1_USER��,��4p���D�0��VEL,2 �0���2�5S�I�|�w�MTN�CFG}1��  ���Oy�NORE��3��26�0SI���� ���\�UX-�ܑPD�E�A $KE�Y_����$J3OG<EנSVIA�0WC�� 1DSWy���
��CMULT�G�I�@@C��2� �4 �#t�+�z�X�YZ��|�����z� ޜ@_ERR��� ��S L�-���@��|s0BB$BUF-@qX17ࡐMOR�7� H	�CU�A3��z�1Q�
��3���'$��FV��2�,SbG�� � $SI�@ G�0�VO B`נOBJyE&�!FADJU�#EELAY' ���SD�WOU�мE1PY�.��=0QT i8�0�W�DIR$bap�pےʠDYN$բHeT�@��R�^��X����OPWOR�K}1�,�SY�SBU@p 1SOP��aR�!�jU�k�PR��2�ePA�0�!�c�u� 1OP��UJ��a'�D�QIMA�G�A	��`i�IM�ACrIN,�bsRGOVRD=a�b�0�aP�`sʠ� �^uz�LP�B�@��!PMC_E,�Q��EN@�M�rǱ��1ŲL7�=qSL&�~0���?$OVSL\G*E���*E2y�Ȑ�_ =p�w��>p�s���s	�����y��t�#}1�� @�@;���OE�R	I#A��
N��X�s��f�{��PL}1��,RTv�m�ATUS>RBTRC_T(qR��B �����$ �Ʊ8��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���UP(4����PX��؆�q�3�w� �PG��5� $S�UB������t�J?MPWAITO��s��LOyCFt�!D=��CVF	ь�y���R�`�0��CC_CT�R�Q�	�IGNR�_PLt�DBTB2m�P��z�BW)���2�0U@���IG�a��=Iy�TNLN��Z�R]aK� N��`B�0��PE�s���r��f�S�PD}1� L	�A`�`gఠ�S��UN��{���]�R!�`BDL�Y�2���6�PH_�PK�E��2RETRIEt��2�b���;FI�B� �����8� 2��0DB�GLV�LOGS�IZ$C�KTؑUdy#u�D7�_�_T1@�EM�@C\1aA��ℽR��D�FCHE3CKK�R�P�0��e��@&�(bLEc�" PA9�T���P�C�߰PN�����A�Rh�0���Ӯ�PO��BORMATT naF�f1h���2�S���UXy`	���PL|B��4�  rE�ITCH3�8PL�)�AL_ � �$��XPB�q� C�,2D�!��+2�J3�D��� T�pPD�CKyp��oC� _AgLPH���BEWQo���� ��I�wp� � �b@PA�YLOA��m�_1�t�2t���J3AR���؀դ֏�laTI�A4��5��6,2MOMCP�����������0BϐAD�����\���PUBk`R�Ԁ;���;������z4�` I$PI\D s�oӓ1yՕ�w�2�w�UZ��I��I��I�〛�p����n���y��e`�9S)bT�SPEED� G��(�Е�� /���Е�`/�e�>���M��ЕSAMP��6V��/���ЕMO�@ 2@�A��QP�� �C��n����������� LRf`kb�ІE9h�EIN09��7S.�В9
yPy�GA�MM%S���D$GGET)bP�cD]Ԛ�2
�IB�q�IN�G$HI(0;A��$LREXPA8)LWVM8z�)��g���C5�C�HKKp]�0�I_��h`eT��n�q���eT,���� ��$�� 1��iPI� RCH_D`�313\��30LE�1��1\�o(Y�7 �t�M�SWFL �M��SCRc�7�@�&��%�n�f�SV���P�B``�'�!�B�sS_�SAV&0ct5B3NO]�C\�C2^�0� mߗ�uٍa��u���u:@e;��1���8��D�P ���������)� �b9��e�GE�3���V�ve�Ml�� � �YL��QNQSRlbfqXG�P �RR#dCQp� �S:AW70�B�B[�CdgR:AMxP�KCL�H����W�r�(1n�g�M�!o�� �F�P@}t$WP�u�P r�� P5�R<�RC�R�� %�6�`��� ��qsr %X��OD�qZ�Ug��ڐ>D� ��OM#w�J?\?n?�?�?P��9�b"�L]�_��� |��X0��bf ��qf��q`�ڏgzf��9Eڐ� Ag�"��ܰ��FdPB���PM�QU�� �� 8L�QCOU�!5�QTHI�HO�QBpHYSY�ES���qUE�`�"�O.���  �P�@�\�UN���Cf�O�� P��Vu�x�!����OGRAƁ�cB2�O�tVuITxe �q:pINFO������{�qcB�e�O�I�r� (�@SLEQS��q��p�vgqyS���� 4L��ENABDRZ�PTIONt�����Q����)�GCF��G�c$J�q^r�� �R���U�g��rS�_ED����� ��F��PK��E�'NU߇وAUT<$1܅COPY���(��n�00MN��^�PRUT8R ��Nx�OU��$G�[rf���RGADJ����*�X_:@բ�$�����P��W��P���} ��)�}�EX��YCDR|�NSr.��F@r�LGO��#�NYQ_FREQR�W� �#�h�TsLAe#����ӄ ��CRE� s�IFl��sNA��%a��_Ge#STATUxI`e#MAIL�� ���q t��������ELEM�� �|/0<�FEASI?� B��n�ڢ�vA�]� � I�p��Y!q�]�t#A�ABM���E�p<�VΡY�BASR�Z��S�UZ��0�$q���RMS_TR;�qb ���S�Y�	�ǡ��$���>C��Q`	� 2� _�TM������ ̲�@ �A��)ǅ�i$'DOU�s]$Nj����PR+@3���rGR�ID�qM�BARS� �TY@��OTO��p��� Hp_}�!Ⱦ���d�O�P/�� � �p�`PORp�s��}���SRV��Y)����DI&0T��@��� #�	�#�4!�U5!�6!�7!�8��e�F�2��Ep$VALUt��%��ֱ|��/��� ;��1�q�����(_�AN�#�ғ�Rɀ(���TOTAL��S���PW�Il��REGGEN�1�cX��`ks(��a���`TR��R��_S� ��1ଃAV�����⹂Z�E���p�q��Vr���V_�H��DA�S����S�_Y,1�R4�S� A�R�P2� ^�IG_SE	s����å�_Zp��C_�Ƃ�E�NHANC�a�/ T ;�������INT�.��@F�Psİ_OVRsP��`p�`��Lv��o���7�}��Z�@�SLG�AA�~�25�	���D��S�BĤDEb�U�����TE�P>���� !Y���
�J��$2�IL_�MC�x r#_��`TQ@�`��q���'�BV��C�P_� 0�M��	V1�
V1�2��2�3�3�4�4�
�!���� � �m�A�2IN~VIABP���1�2�U2�3�3�4��4�A@-�C2���{p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KE�EP_HNADD"!!`$^�j)C�Q��A�$��"	��#O�a�_$A�!�0�#i��#REM�"�$��½%��!�(U}�e�$HP�WD  `#S�BMSK|)G�q�U2:�P	�COLLAB� �!K5�B��h ��g��pITI1p{9p#>D� ,�@�FLAP��$SY�N �<M�`C6��~�UP_DLYAA=�ErDELA�0�Z��Y�`AD�Q@a�QSKIP=E� i���XpOfPNTv�A�0P_Xp�rG�p �RU@,G��:I+�:IB1 :IG�9JT�9Ja�9Jn��9J{�9J9<��RA=s� X���4��%1�QB� NFLIC�s�@J�U�H�LwNO_H�0�"?��R�ITg��@_PAz�pG�Q� ��
^�U��W��LV�d�NGRLT�0_q���O�  " ��OS��T_�JvA V	�APPR�_WEIGH�sJg4CH?pvTOR��vT��LOO��]�+�"tVJ�е�ғA�Q�U��S�XOB'�'�@aJ�2P���7�X�T �<a43DP=`Ԡ\"<a8�q\!��RDC��LW� �рR��R�`� �RV��jr�b��RGE��*��cN�F�LG�a�Z���SP9C�s�UM_<`^2TH2NH��P.a� 1� m`E�F11��� l�Q �!#� <�p3AT � g�S�&�Vr�p�tMq��Lr���HOMQEwr�t2'r�-@?Qcu��w3'r�������w4'r�'�9�K�]�o����w5'r뤏��ȏPڏ����w6'r�!�@3�E�W�i�{��w7'r힟��ԟ����w8'r��-�?�Q�c��u��uS$0�q�p �� sF��`)a�"`P�����`/���-��IO[M�I֠���*�POWE��# ��0Za*���� �5��$DS=B GNAL���0�Cp��)�S232N3�� �~`��� �/ ICEQP��PE�p��5PIT����O�PBx0��FLOW�@TRvP��!U����CU�M��UXT��A��w�ERFACt�� U��ɲ;CH��� tQ  1_��>�Q$����SOM��A�`T�P.#UPD7 A�ct�T��UEX@�ȟÎU EFA: X"�1RsSPT�����T 
��PPA�0o񩩕`EXP�IOS���)ԭ�_���%��C�#WR�A��ѩD�ag���`ԦFRIEND�saC2UF7P����TwOOL��MYH �C2LENGTH_VTE��I��Ӆ�$SE����UFOINV_����RGI�{QITI�5B��Xv��-�G2-�G17�w�SG�X�"��_��UQQD=#�� �AS��d~C�`��|q�� �$$C/�=S�`�����S0�Ȱ����VERSIܕ ��Ȱ��5��I��������AoAVM_Y�2 �� ?0  �5��C�rO�@�r� r�A	 ����S0����������������`
?QY�BS����1��� <-���� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�Oi{CC�@XLMT��v�C�  ��D�IN�O�A�Dq�EX�E�HPV_��A�TQz
��LAR�MRECOV ��RgLMDG� *�5�OLM_IF *��`d�O�_�_�_�_j��_'o9oKo]onm, 
��odb��o�o`�o�o^��$� z, A   2D{��PPINFO u[ �Vw��������`���� ���*��&�`�J� ��n�����DQ�� ��
��.�@�R�d�v����������a
PPLoICAT��?��P��`H�andlingT�ool 
� 
�V8.30P/4�0Cpɔ_LI
�883��ɕ$M�E
F0G�4�-
398��ɘ�%�z�
�7DC3�ɜ
�NWoneɘVr��оɞ@6d� �Vq_ACTIV�U��C죴�MO�DP���C�I��HGAPON��񿰷OUP�1*��� i�m����Қ_l����1*�  �@����f�����Q����Կ�@�
���{�� ����5�Hʵl�K�HTTHKY_��/� M�SϹ��������� %�7ߑ�[�m�ߝߣ� �����������!�3� ��W�i�{������ ��������/���S� e�w������������� ��+�Oas ������� '�K]o�� ������/#/ }/G/Y/k/�/�/�/�/ �/�/�/�/??y?C? U?g?�?�?�?�?�?�? �?�?	OOuO?OQOcO �O�O�O�O�O�O�O�O __q_;_M___}_�_��_�_�_�_�_kŭ�T�Op��
�DO_C�LEAN9��pcN/M  !{衮o��o�o�o�o��DS�PDRYRwo��H	I��m@�or�� �������&�88�J���MAXݐWdak�H�h�XWd�d�|��PLUGGW��Xgd��PRC)pB��`�kaS�Oxǂ2DtSEGF0�K� �+��o�or�����������%�LAP Ob�x�� �2�D�V� h�z�������¯ԯ�>+�TOTAL�����+�USENUO��\� e�A�k­�RGDISPMMC.�e��C6�z�@@Dr�\�OMpo�:�X�_�STRING 1�	(�
�M�!�S�
��_I�TEM1Ƕ  n ������+�=�O� a�sυϗϩϻ����������'�9�I�/O SIGNA�L��Tryout Modeȵ�Inpy�Sim�ulateḏ�Out��OV�ERRLp = 1�00˲In c�ycl�̱Prog Abor���̱u�Statu�sʳ	Heart�beatƷMH� Faul	��Aler�L�:�L�^�p��������� ScûSaտ��-� ?�Q�c�u��������� ������);M8_q��WOR.�û ������ +=Oas��������//'.PO����M �6/p/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�?p�?�?�?H"DEVP. �0d/�?O*O<ONO`O rO�O�O�O�O�O�O�O�__&_8_J_\_n_PALT	��Q�o_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�op�o�o�_GRIm� û9q�_as�� �������'� 9�K�]�o�������'�R	�݁Q���� )�;�M�_�q������� ��˟ݟ���%�7�<I�ˏPREG�^�� ��[�����ͯ߯�� �'�9�K�]�o����������ɿۿ�O��$�ARG_� D ?�	���0���  	�$O�	[D�]�D��O�e�#�SBN�_CONFIG S
0˃���}��CII_SAVE  O�����#��TCELLSET�UP 0�%  OME_IOO��O�%MOV_H8������REP��J���UTOBACK�����F�RA:\o� XQ�o���'`��o���� �� f�o�����*�!�3�`�Ԉ��f��� ��������o�{��&� 8�J�\�n�������� ����������"4F Xj|����p��끁  ���_i�_\ATBC�KCTL.TMP� 6.VD GIF ��BN`r��o�N�R��f�IKNI�P�Օ�c�?MESSAG������8��ODE_D����z��O�0�c�oPAUSM!!�0�? (73�U/g+(Od/�/x/�/ �/�/�/�/�/???�P?>?t?1�0$: TSK  @-��T�f��UPDT��d��0
&XWZD_E�NB����6STAp�0��5"�XIS��?UNT 20Ž�� � 	 �� $� 1����q�T?ŵӀ��G��2�H����zF�OTo�}Cw�g�^�	���.�O�O�O�O�/_2FMET߀2�CMPTAA Q@�ԑ�A��@����@��@����rK5��5��(d5��P5��r�5F*5��338]SCRD�CFG 1�6��Ь�Ź� _�_oo(o:oLo��o�Q���_�o�o�o�o �o�o]o�o>Pb�t���o9�i�G�R<@M/�s/NA��/�	i��v_�ED�1�Y� �
 �%-5E�DT-�'�GE�TDATAU�o�9A�u?�j�H�o�f��\��A��  ���2�&�!�E���:IB���~�ŏ׏m����3��&۔�� D��ߟJ�����9�ǟ�4���ϯ�(���@�]�o�����5N� �����(�w��)�;�ѿ_��6ϊ�gϮ� (�CϮ���ϝ�+��7��V�3�z�(��z� ����i����8��&���~�]���F�ߟ�5����9~������]����Y�k�����CR�!ߖ���W� q���#�5���Y��p$�?NO_DEL��r�GE_UNUSE���tIGALLO�W 1��(�*SYSTE�M*S	$SERV_GR�V� n: REG�$�\� NUM�
���PMUB U�LAYNP\�PMPAL�COYC10#6 <$\ULSU��8:!�Lr�B�OXORI�CU�R_��PMC�NV�10|L�T4DLI�0��	����BN/`/ r/�/�/�/�/�/���p�LAL_OUT ��;���qWD_ABOR=f�q;0ITR_RTN�7y�o	;0NONS�0��6 
HCCFS�_UTIL �#<�5CC_@6A ;2#; h ?�?��?O#O6]CE_O�PTIOc8|qF@RIA_Ic Rf5Y@�2�0F�Q��=2q&}�A_�LIM�2.�k ��P�]B��K*X�P
�P�2O�QK��B�r�qF�P�Q5T1)TR�H��_:JF_PARA�MGP 1�<g^&S�_�_�_�_�V�C�  C�d��`�o!o`�`�*`�`�Cd��Ti�i:a:e>eBa�GgC��`� D� D�	�`�w?��2H=E ONFI� E?n�aG_P�1#; ���o�1CUgy�aKP7AUS�1�yC ,������ ���	�C�-�g�Q� w���������я���r�O�A�O�H�L_LECT_�B�IPV6�EN. QF�3��NDE>� �G��71234567890��sB�pTR����%
 H�/%)�������W� ��0�B���f�x���� ����ү+�����s� >�P�b���������� ο��K��(�:ϓ��^�|��B!F� |�I|�IO #��<U%e6�'�9�K߶��TR�P2$��(`9X�t�Y޼`%��x�ڥH��_MOR��3&�=��@XB��a��A�$��H�6�l�~���~S��'�=�r_A?�a�a`�᢭@K��R�dP��)<F�ha�-�_�'�9�%
�k��G� ��%Z�%��u`�@c.�PDB���+���cpmi�dbg��	�`:�  2+' �qTR���p��N  ���@e�@f/����]܌0`a�w<�^��@r�@swg�$�+�`@�wfl��q��ud1:��:J��DEF �*ۈ��)�c��buf.txt�����_L64?FIX ,���� ��l/[Y/�/}/�/�/ �/�/
?�/.?@??d? v?U?�?�?�?�?�?�?|,/>#_E -���<2ODOVOhOzO�OV6&IM��.o�YU�>���d�
�IMMC��2/����dU,�C��20�M�QT:U>w�Cz  B�i��A���A����Au�gB3�*�CG�B<�=�w�i�B.��B����B��5B��$�D�%B����ezVC�q�C��v�D���D�-lE\D�n �hw��29"��22o�D|������ ���C�ZC����
�xObfi�D4cdv`D��`�/�`v`s]E�D �D�` E4��F*� Ec���FC��u[F����E��fE��f�Fކ3FY��F�P3�Z��@��33 ;��>LS���Aw�n,a@��@e�5Y���a����`A��w�=�`<#����
��?�ozJR�SMOFST �(�,bIT1��D2 @3��
д����a���;��bw?���<�M�N/TEST�1O�CER@�4��>VC5`#A�w�Ia+a�aOR�I`CTPB�U�C��`4���r��:d�����qI?�5���qT_�PROG ��
�%$/ˏ�t���NUSER  �U������KEY_TBL  �����#a��	
��� !"#$%&�'()*+,-.�/��:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s������LCK�x
����STAT/���s_AUTO_D�O �	�c�IN?DT_ENBP���1Rpqn�`�T2�����STOr`���XCΔ� 26���8�
SONY XC�-56�"b�����@��F( А{�HR50w����>�P�7b�t�ACff����ֿ� Ŀ ����C�U�0�yϋ� fϯ��Ϝ���������-ߜ�TRL��LE�TEͦ ��T_�SCREEN }��kcs�����U�MMENU� 17�� < ܹ���w������ ���K�"�4��X�j� ������������5� ��k�B�T�z����� ����������. g>P�t��� ���Q(: �^p����/ ��;//$/J/�/Z/ l/�/�/�/�/�/�/�/ 7?? ?m?D?V?�?z? �?�?�?�?�?!O�?
O WO.O@OfO�OvO�O�O�(y��REG 8�y����`�M�ߎ�_MANUAL��k�DBCO��RI�GY�9�DBG_E7RRL��9�ۉqa��_�_�_ ^Q�NUMLI�pϡ�pd
�
^QPXW�ORK 1:����_5oGoYoko}oӍD�BTB_N� ;T�����ADB_AWAYfS��qGCP 
�=�p�f_AL�pR��bBbRY�[�
�WX_�PW 1<{y�n�,��%oc�P��h_M&��ISO��k@L��s�ONTIMX��&
���vy
��2sMOTNEND��1tRECORD ;1B�� ���sG�O�]�K��{�b ��������V�Ǐ�]� ���6�H�Z����� ����#�؟������ 2���V�şz������� �ԯC���g��.�@� R���v�寚�	���п ���c�χ�#ϫ�`� rτϖ�Ϻ�)ϳ�M� ��&�8ߧ�\�G�U����8��������K� �����6��%RC7�n���ߤ������A�4���$����H�3�A�~��; �������9���]������|�B#Zl����zTOLERE�N\�rB�'r�`L���^PCSS_CCSCB 3C>y�`IP��}�~� <�_`r�K�@����/�{�� 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�OX_�~�LL� D���fFY C[C��PZP^r_W A� p� �s�p��Q �\	 CA�p�Q�_�[? ��_�[oU�p��P�pSB�V�c��(a�PWoio{h+�o³X�o�oY���[	r�hLP����ޮ?�����:�3߮|�wc��aD@V�B��|�G����+��Kۃ �otGhXGr��So����eB �  =��Ͷa>L�tYB�� �pC�p�q�aA"�H�S�Q-� �q���ud�v������AfP ` 0��c�D^P��p@�a�
�QX��\ DaW>� �a9P��b �e:�L�^�h�Hc�́PQ�R�Q�PU�z� ֟�o\^��-�?��`c�u����zCz�	ů�b2�Щ�_�� ��S̡0��]�0�.�����.a��F�X� ѿUҁп�VSȺ�NSTCY 1E��]�@rIϫ�K� ]�oρϓϥϷ����� �����#�5�G�Y�k��}ߏߒ��DEVI�CE 1F5� E_����	� ��?�6�c��V|㰟����_HNDGD �G5�VP���R�LS 2H�ݠ��/�A��S�e�w����� ZPA?RAM I�Fg�He�RBT 2-K��8р<��WPVpC�{��,`¢PQ�Z�z��%{�C*  �2�jMT`v�,`"nPB,  s��M� }�gT�g���
B��!�bc y�[2Dchz ����/��/�gT#I%D��C��` b!�R��A���A,��Bd�ךA�;���_C4kP�!2�C��$Ɓ�]ߚffA�À�W�B�� �| ���/�/�T (��54a 5�}%/7/d?/M? _?q?�?�?�?�?�?O �?OO%O7OIO�OmO O�O�O�O�O�O�O�O J_!_3_�_�_3�_�_ �_�_�_o�_(ooLo ^oЁ=?k_IoS_�o�o �o�o�o�o�o# 5G�k}��� ����H��1�~� U�g�y�ƏAo�Տ� ��2�D�/�h�S���go ����ԟ����ϟ�� �R�)�;���_�q��� �������ݯ�<�� %�7�I�[�m������� ��}�&��J�5�n� YϒϤϏ��ϣ�ѿ� �����F��/�Aߎ� e�w��ߛ߭������� ��B��+�x�O�a�� ����������,��� %�b�M���q������� ��������L# 5�Yk}���  ��61C Ug������ ��	//h/���/w/ �/�/�/�/�/
?�/.? @?I/[/1/_?q?�? �?�?�?�?�?�?OO %OrOIO[O�OO�O�O �O�O�O&_�O_\_3_ E_W_�_?�_�_�_�_ �_"ooFo1ojoE?s_ �_�om_�o�o�o�o�o 0f=Oa� �������� �b�9�K���o���Ώ ��[o��(��L�7��I���m������$D�CSS_SLAV�E L����ё��__4D  љ�◿CFG Mѕ��������_FRA:\ĐL-��%04d.CSVn��  }�� ���[A i�CHq�z�������|�����"������Ρޯ̩�Ґ�-��*����_C�RC_OUT �N������_F�SI ?њ ����k�}��� ����ſ׿ ����� H�C�U�gϐϋϝϯ� �������� ��-�?� h�c�u߇߽߰߫��� ������@�;�M�_� ������������� ��%�7�`�[�m�� �������������� 83EW�{�� ����/ XSew���� ���/0/+/=/O/ x/s/�/�/�/�/�/�/ ???'?P?K?]?o? �?�?�?�?�?�?�?�? (O#O5OGOpOkO}O�O �O�O�O�O _�O__ H_C_U_g_�_�_�_�_ �_�_�_�_ oo-o?o hocouo�o�o�o�o�o �o�o@;M_ �������� ��%�7�`�[�m�� ������Ǐ������ 8�3�E�W���{����� ȟß՟����/� X�S�e�w��������� �����0�+�=�O� x�s���������Ϳ߿ ���'�P�K�]�o� �ϓϥϷ��������� (�#�5�G�p�k�}ߏ� �߳����� ����� H�C�U�g����� �������� ��-�?� h�c�u����������� ����@;M_ �������� %7`[m �������/ 8/3/E/W/�/{/�/�/ �/�/�/�/???/? X?S?e?w?�?�?�?�? �?�?�?O0O+O=OOO�xOsO�O�O�O�O�C��$DCS_C_F�SO ?�����A P �O�O_?_:_ L_^_�_�_�_�_�_�_ �_�_oo$o6o_oZo lo~o�o�o�o�o�o�o �o72DVz �������
� �.�W�R�d�v����� ��������/�*� <�N�w�r��������� ̟ޟ���&�O�J� \�n���������߯گ ���'�"�4�F�o�j� |�������Ŀֿ�������G�B�T��OC_RPI�N_jϳ� ���ς��O����1�Z�,U��NSL��@&�h� ����������"��/� A�j�e�w����� ��������B�=�O� a��������������� ��'9b]o �������� :5GY�}� �����/// 1/Z/U/g/y/�/�/�/ �/�/�/�/	?2?-??? Q?z?u?��ߤ߆?�? �?�?OO@O;OMO_O �O�O�O�O�O�O�O�O __%_7_`_[_m__ �_�_�_�_�_�_�_o 8o3oEoWo�o{o�o�o �o�o�o�o/ XSew���� ����0�+�=�O� x�s���������͏ߏ ���'�P�K�]�o������ �PRE_C�HK P۪�A� ��,8�2��� 	 8�9�K���+�q��� a�������ݯ�ͯ� %��I�[�9����o� ��ǿ��׿���)�3� E��i�{�YϟϱϏ� ����������-�S� 1�c߉�g�y߿��߯� ���!�+�=���a�s� Q���������� ����K�]�;����� q�������������# 5�Ak{� �����C U3y�i��� ���/-/G/c/ u/S/�/�/�/�/�/�/ ??�/;?M?+?q?�? a?�?�?�?�?�?�?�? %O?/Q/[OmOO�O�O �O�O�O�O�O_�O3_ E_#_U_{_Y_�_�_�_ �_�_�_�_o/ooSo eoGO�o�o=o�o�o�o �o�o=-s �c������ �'��K�]�woi��� 5���ɏ�������� 5�G�%�k�}�[����� ��ן�ǟ����C� U�o�A�����{���ӯ ����	��-�?��c� u�S�������Ͽ῿� ����'�M�+�=σ� ��w�����m������ %�7��[�m�K�}ߣ� �߳��߷����!��� E�W�5�{��ϱ��� e�������	�/��?� e�C�U����������� ����=O-s ����]��� �'9]oM� ������/� 5/G/%/k/}/[/�/�/ ��/�/�/�/?1?? U?g?E?�?�?{?�?�? �?�?	O�?O?OOOO uOSOeO�O�O�/�O�O �O_)__M___=_�_ �_s_�_�_�_�_o�_ �_7oIo'omoo]o�o �o�O�o�o�o!�o 1W5g�k}� �����/�A�� e�w�U�������я� �o����	�O�a�?� ����u���͟���� �'�9��]�o�M��� ������ۯ��ǯ�#� ůG�Y�7�}���m��� ſ�����ٿ�1�� A�g�E�wϝ�{ύ��� ����	�߽�?�Q�/� u߇�e߽߫ߛ����� ���)���_�q�O� ����������� ��7�I���Y��]��� ������������!3 WiG��}� ���%�A� 1w�g���� ��/+/	/O/a/?/ �/�/u/�/�/�/�/? �/9?K?�/o?�?_? �?�?�?�?�?�?O#O OGOYO7OiO�OmO�O �O�O�O�O_�O1_C_ %?g_y__�_�_�_�_ �_�_�_o�_+oQo/o Ao�o�owo�o�o�o�o �o);U__q �������� %��I�[�9����o� ��Ǐ�����ۏ!�3� M?�i��Y������� ՟�ş����A�S� 1�w���g�����������ӯ�+�=��$D�CS_SGN �QK�c��7m�� 16-MA�Y-19 10:�20   O�l�4�-JANt�08:�38}����� N.DѤ�����������M4�o���Im��P�Zۘq��  O�VE�RSION �[�V3.5.�13�EFLOG�IC 1RK���  	����P�?�P�N�!�P�ROG_ENB � ��6Ù�o�U?LSE  TŇ��!�_ACCLI�M����Ö���WRSTJNT��c��K�EMO�x̘��� ���INIT S.�G�Z����OPT_SL ?�	,��
 	�R575��Y�74j^�6_�7_�50��1��2_�@ȭ��<�TO  Hݷ���V�DEX��d�c����PATHw A[�A\��g�y��HCP_CLNTID ?��6� @ȸ�����IAG_GRP� 2XK� ,`����� �9�$�]�H������1234567�890����S�� |�������!�� ��H���;�dC�S���6�� ���.�R v�f��H�� //�</N/�"/p/ �/t/�/�/V/h/�/? &??J?\?�/l?B?�? �?�?�?�?v?O�?4O FO$OjO|OOE��O y��O�O_�O2_��_�T_y_d_�_,
�B^ 4�_�_~_`Oo�O &oLo^oI��Tjo�o.o �o�o�o�o �O'�_ K6H�l��� ����#��G�2��k�V���B]�?g��?����>ط���*��{��V>h)>���ž4	��d��D��?��ihD=P���Ƈ�����(��L�B\ډC�*����U{���>���:������ߟʟܟ���CT_�CONFIG �Y��Ӛ��egU���STBF/_TTS��
��b�����Û�u�O�MA�U��|��MSW_�CF6�Z��  ~�OCVIEW��3[ɭ������ -�?�Q�c�u�G�	��� ��¿Կ������.� @�R�d�v�ϚϬϾ� ������ߕ�*�<�N� `�r߄�ߨߺ����� ����&�8�J�\�n� ���!���������� ���4�F�X�j�|�����RC£\�e��! *�B^������C�2g{�SBL_FAULT ]��|ި�GPMSKk���*�TDIAG �^:�աI���UD1: 67�89012345�G�BSP�-? Qcu����� ��//)/;/M/t
J��
@q��/$��TRECP��

 ��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOi/{/�xO�/UMP_OP�TIONk���AT�R¢l��	�EPM�Ej��OY_TEM��È�3B��J�P�AP�DUN�I��m�Q��YN_?BRK _ɩ��EMGDI_ST�A"U�aQK�XPNCv_S1`ɫ �FO(�_�_�^
�^dpOo o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{�E�� ���y�Q��� � 2�D�V�h�z������� ԏ���
��.�@� R�d��z�������˟ ����%�7�I�[� m��������ǯٯ� ���!�3�E�W�i��� ������ÿݟ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�{�iߗߩ߻� տ������'�9�K� ]�o��������� �����#�5�G�Y�s� �ߏ�����i������� 1CUgy� ������	 -?Qk�}���� �����//)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? u?�?�?�?��?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_m?w_�_�_ �_�?�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K e_W����_�_� ���#�5�G�Y�k� }�������ŏ׏��� ��1�C�]oy��� �����ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� ��g�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�_�i�{� �ߟ߹���������� �/�A�S�e�w��� �����������+� =�W�E�s������ߧ� ������'9K ]o������ ��#5O�a�k }�E������ //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -?GYc?u?�?�?� �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_Q?[_ m__�_�?�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /I_Sew��_ �������+� =�O�a�s��������� ͏ߏ���'�A3� ]�o�������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��9�K�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ���������ߑ�C� M�_�q߃ߝ��߹��� ������%�7�I�[� m����������� ���!�;�E�W�i�{� �ߟ����������� /ASew�� �����3� !Oas����� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?+=G?Y?k? !?��?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	_#? 5??_Q_c_u_�?�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o-_7I[ m�_������ ��!�3�E�W�i�{� ������ÏՏ���� %/�A�S�e�q��� ����џ�����+� =�O�a�s��������� ͯ߯����9�K� ]�w���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� �'�1�C�U�g߁��� �߯���������	�� -�?�Q�c�u���� ��������m��)�;� M�_�y߃��������� ����%7I[ m������ ��!3EWq�{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/�/+? =?O?i_?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O��O? �$ENE�TMODE 1a�j5� + 0054_�F[PRROR_P�ROG %#Z%�6�_�YdUTABL/E  #[t?�_��_�_gdRSEV_�NUM 2R  ��-Q)`dQ_�AUTO_ENB�  PU+SaT_N�O>a b#[EQ�(b  *��`�J�`��`��`4`+�`p�o�o�oZdHIS%c�1+PSk_ALM �1c#[ �4�l0+�o;M_�q���o_b``  #[aFR�zP�TCP_VER �!#Z!�_�$E�XTLOG_RE�Q�f�Qi,�SI�Z5�'�STKR��oe�)�TOL � 1Dz�b�{A '�_BWD�pp��Hf��D�_DI��7 dj5SdDTx1KRņSTEPя��P��OP_DO�t�QFACTOR_Y_TUN�gd<��DR_GRP 19e#YNad 	����FP��x��� ��� ��$�f??�� ���ǖ�� ٟ�ԟ���1��U� @�y�d�v�����ӯ�����LW
 J��^�,��tۯ�j��U���y�B�  B�୰���$  Ay@��s�@UUUӾ��������E�� �E�`F@ F��5U/�,��L����M��Jk��Lzp�JP�ߣFg�f�?��  s��9�Y�9}�9���8j
�6���6�;��������� �!�� ��~�ߢ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����⣆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7���; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  C��0����(7�?�<B�?B����2�ٸ*9�N SMTT#t�[)��X�4�$HO�STCd1ux����?�� MC�x��;zOx��  27.0�@1�O  e�O�O	_ _-_;Z�O^_p_�_�_��LN_HS	anonymous�_�_�_�oo1o yO��Fh Fk�O�_�o�O�o�o�o �oJ_'9K]�o �_�����4o �XojoG�~�o^��� ����ŏ����� 1�T���y������� ����,�>�@�-�t� Q�c�u���������ϯ ���(�^��M�_� q�����ܟ� �ݿ� �H�%�7�I�[Ϣ�� �ϣϵ����l�2�� !�3�E�Wߞ���¿Կ ����
�������/� v�S�e�w������ �������+�r߄� ��s�����߻����� �����'9K]�� �������4� F�X�j�l>��}� �����// 1/T��y/�/�/�/��/.D\AENT 1=v
; P!J/?  ��/3?"? W??{?>?�?b?�?�? �?�?�?O�?AOOeO (O�OLO^O�O�O�O�O _�O+_�O _a_$_�_ H_�_l_�_�_�_o�_ 'o�_Koooo2o{oVo �o�o�o�o�o�o5 �oY.�R�v���zQUICCA0���3��t14��"����t2��`�r��ӏ!ROUTE�Rԏ��#�!P�CJOG$���!�192.168�.0.10��sC�AMPRTt�P�!�d�1m�����RT�폟�����$NAM�E !�*!R�OBO���S_C�FG 1u�) ��Aut�o-starte�dFTP& ��=?/֯s���� 0�B��f�x������� ��S������,�� �������ϼ�ޯ���� �����ʿ'�9�K�]� oߒ�ߥ߷�������8��SM%y� {�U�ό������� ����
��.�@�c����v������������z �%�7�I�K�8�\ n���k���� �3�FXj|�����a��7 /M*/</N/`/ r/9�/�/�/�/��/ �/?&?8?J?\?�m? ���?�//�?�?O "O4O�/XOjO|O�O�O �?EO�O�O�O__0_ w?�?�?�?�O�_�?�_ �_�_�_o�O,o>oPo boto�_o�o�o�o�o �oK_]_o_L�o�_ �o�����o� � �$�6�Y�Y�~���𢏴�ƏZ�_ERR� w3�я�PDUSIZ  g��^�p���>�W�RD ?r�Cq��  guestb�Q�c�u��������`�SCDMN�GRP 2xr�;���H�g��\�b�K� 	P01.00 8`��   � ��   B  ���� ���_H���L��L�}�L�����O8�`����l�����a4�U  �Ȥ� �8����\���)�`�;��������d�.�@�R�ɛ_GWROUېy������	ӑ���QU�PD  ?u�����İTYg�����TTP_AUT�H 1z�� <�!iPenda�n��-�l���!�KAREL:*8-�6�H�KC]�m���U�VISION SET���ϴ�!�����R�0�� H�Bߏ�f�x��ߜ߮����CTRL {�����g�
&�?FFF9E3��At�FRS:DEF�AULT;�F�ANUC Web Server;� )����9�K��ܭ����������߄WR_�CONFIG �|ߛ ;��I�DL_CPU_P5CZ�g�B�I�y�w BH_�MINj��)�}�GNR_IO���g���a�NPT?_SIM_D_������STAL_S�CRN�� ���T�PMODNTOL8������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMAST�E��ɾeSLAV�E ~��c�O�_CFGٱBU�O�O@CYCL�En>T�_ASG� 1ߗ+�
  ����//+/=/ O/a/s/�/�/�/�/���NUM��
�@IPCH�^R?TRY_CNZ��@�@��������1 @kI�+E��z?E�a�P_MEMBERS 2�ߙ�� $���2����ݰ7�?�9a�SDT�_ISOLC  �����$J23�_DSM+�3J?OBPROCN���JOG��1�+��d8�?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSRE�QO��KANJI_����a[�MONG ����b�yN_ goyo�o�o�o�Y�`3	�<� ��e�_ִ���_L���"?`EY�LOGGINL�E�������$L�ANGUAGE Y��<T� {q��LGa2�	�b����g�xP��  *��g�'��b����>�MC:�\RSCH\00�\<�XpN_DISP �+G�H��O��O߃LOCp�D�z���AsOGB?OOK ����`��󑧱����X� ����Ϗ����a�*��	p������!�m��!���=p_B�UFF 1�p��2F幟���՟�D� Collaborativǖ ���F�=�O�a�s��� ����֯ͯ߯����B�9�K���DCS ��z� =��� '�f��?ɿۿ���H@�{�IO 1��# ~?9Ø��9�I� [�mρϑϣϵ����� �����!�3�E�Y�i� {ߍߡ߱��������-E��TMNd�_B� T�f�x�������� ������,�>�P�b��t�������L��SE�VD0��TYPN1�$6���Q�RS"0&��<2FLg 1�"�J0��� �����G�TP:pOF�NGNAM1D�mr�t7UPS�GI"5�a�O5�_LOAD�N@G %�%DF_MOTN�y��� MAXUAL�RM�'���(��_PR"4F0d��1��B_PNP� V �2�C	MD_R0771ߕ�B�L"8063%�@ �_#?�ߒ|/�C��z�6��/��z�/Po@P 2��+W �ɖ	T ?	t  ��/�% W?B?{?�k?�?g? �?�?�?O�?*OONO `OCO�OoO�O�O�O�O �O_�O&_8__\_G_ �_�_u_�_�_�_�_�_ o�_4ooXojoMo�o yo�o�o�o�o�o�o 0B%fQ�u� �������>� )�b�M�����{����� ���Տ��:�%�^��p�S�������D_LDXDISAp�B�MEMO_A�PjE ?C
 �,�(�:�L��^�p������ISCw 1�C ��� �4�������4���X���C_MSTR� ���w�SCD 1���L�ƿH� �տ���2��/�h� Sό�wϰϛ��Ͽ��� 
���.��R�=�v�a� �߅ߗ��߻������ �<�'�L�r�]��� ������������8� #�\�G���k������� ��������"F1 jUg����� ��B-fQ��u���h�MK?CFG ����/~�#LTARM_��7"0�0�N/V$� METPUlᐒ3����ND� ADCOLp%A {.oCMNT�/ �%� ����.E#>!��/4�%POSCFz�'�.PRPM�/�9ST� 1���� 4@��<#�
 1�5�?�7{?�?�? �?�?�?�?)OOO_O AOSO�OwO�O�O�O�O�_�A�!SING_�CHK  �/$_MODAQ,#�����.;UDEV }	��	MC:o\�HSIZEᝢ���;UTASK %���%$123456789 �_�U9WTRIG 1���l3%%��9o��"ocoFo5#�VYP�QNe���:SEM_INF� 1�3' �`)AT&�FV0E0po�m)��aE0V1&A�3&B1&D2&�S0&C1S0=>�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o'�� K�������я :�L�3�p�#�5���Y� k�}������$�[�H� ��~�9�����Ưد ��������ӟ�V�	� z�������c�Կ���� 
��.���d��)� ;��Ͼ�q������� ˿<���`�G߄ߖ�I� ��m�ϑϣ����8� J��n�!ߒ�M���������h_NITOR�� G ?�[   �	EXEC1T�/�25�35�45�Q55��P7�75�85�9�0�Қ�4�� @��L��X��d�� p��|�������U2��2��2��2��U2��2��2��2��U223��3���3@�;QR_GRP�_SV 1��k� (�A?��?IܿI���pW�Q_D��^�P�L_NAME �!3%,�!D�efault P�ersonali�ty (from� FD) �RR�2� 1�L6�(L?�,0	l d����� ���//(/:/L/ ^/p/�/�/�/�/�/�/�/ZX2u?0?B?T?�f?x?�?�?�?�?\R< ?�?�?O O2ODOVO�hOzO�O�O�OZZ%`\R�?�N
�O_\TP�O:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHo_)_~o�o�o �o�o�o�o�o 2 DVhz�[omo� ���
��.�@�R� d�v���������Џ�� Ef  F?b� F7��� �  ��!��d ��@�R�6�t���� ��l���ʝ����� ݘ����"� @�F�d���� "𩯹�>ݐA�  ϩU�[�$n�B��E ��~ � @D�  �?�� �?�@��A�@�;f��FH� �;�	l,�	 �|��j�s�d��>��� ��� K�(��Kd$2K� ��J7w�KYJ˷�Ϝ�J�	�ܿ�� @I����_f�@�;z��f�γ��N��� ��	�Xl��������S�ĽÔ�¾X�����5��  ����A?oi#�;��A���� ���l� �Ϫ�-���ܛ�G�G�Ѳ��@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=�����в@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj�a�Be�Ci��@#��Bи�L K� ,ee��^^ȹBР��P�����̠�����ADz ՟�n�3��C�i�@��R�R�Yщ��  ��@� ��Ż���?�ff������n� ɠ#ѱy 9G
(���I�(�@u�P~����t�t���>�����;�Cd;���.<߈<��g�<F+<L �������,�d�,��̠?fff?��?�&&��@��@�x��@�N�@���@T�H �ِ�!-�ȹ�|� �
`������� //</'/`/r/]/�/��eF���/�/�/��/m?��/J?�(E��G�#�� FY�T?�?P?�?�?�? �?�?O�?/OO?OeO k���O�IQOG�?�O 1?�OmO_0_B_T_������A_�_	_��_�_�_ o��A��A0n0 bФ/o C�_Uo8�_�Op��؃o�o��o�o���W����v�oC�E� q�H�d��؜a@q���e�F�BµWB]��NB2�(A���@�u\?��D�������b��0�|�uR�����
x~�ؽ���Bu*C��$�)`�$� ���GC#����rAU�����1�e�G�D�I�mH��� I:�I��6[F���C��I��J��:\IT�H
?~QF�y��p��*J�/ I�8Y�I��KFjʻCe�o��s� ����Џ���ߏ�*� �N�9�r�]������� �����۟���8�#� \�G�����}�����گ ů���"���X�C� |�g�����Ŀ����� ��	�B�-�f�Qϊ� uχ��ϫ�������� ,��P�b�M߆�qߪ� ���߹�������(�� L�7�p�[����������s(���3�:����$���3Ï��d�,�4���@�R��񴲚�xl�~�wa���e��<��wa4 �{�������(L:ueP�P~�A�O�������	����G2W}h ������/�@��O�O7/m/[(d=� s/U/�/�/�/�/�/?��/1??U?C?y?�= � 2 Ef9gF[b��77�9fB)a,a)`C9A`�&`w`@-o�?9de�O-O?OQOpn�?�?�O�O�OD�O9c?�0�A7ht4�w`w`!w`xn
 �O9_K_]_ o_�_�_�_�_�_�_�_��_o#ozzQ ���h��G���$M�R_CABLE �2�h t�a�T� @@�0`�Ae��a�a�a��`ɺ�0�`C�`�aO8��tB�n���yA�aE�M�E��#�o�f�#���0��0�DO���By`��޾*���bE�E��c,��o�g8  ����C�07�d�4
v��d����b��E�ZD&�l�`y`
qC�p�bHE�
v���5D�_)D��)�z�lҠ`��0�q��p�b0�
u�ԋ��b?]�E;h��u/o�c-� �4tH�\�?�9�K�]� o�ԏϏ��
�ɏۏ@����?��eo ��a���������b����� �����`�	 ����@�������% �*�0��6 ��ݐ�����`���	����@�������*,� ,�-�\cO�M �ii���3� �A���%% 2345678901i�B{� f����������j�1����
���`�not sGent3�����;��TESTF�ECSALGR  egfJ�1iqiqš-
:�� �DCb�S�Q�c�u��� 9�UD1:\mai�ntenances.xml��ֿq�� =��DEFAULT-���4\bGRP 2��M�  =��a��{p  �%�Force�so�r check ) ���b�z��p����h5-[ �ϻ�������ϖ�D�%!1st� cleanin�g of con�t. v�ilation��}�Rߗ+��[�ߔߦ߸�ݽ�mech�c�al`����p��0��h5k�@�R��d�v�����(�rol�le_Ƶ�����/���(�:�����Basic quarterly�������,����������M��M��:@�"GpP�a�b`�4��������#C ���M"��{P�bt���Su�ppq�greas!e���?/�&/8/J/\/��C+ g}e��. batn�!y`/��/h5	/�/��/�/? ?_�ѷe�n'�v��/�/��/���?�?�?�?�?�QG=?O�qp"CrB1O��0�/`OrO�O�O`�O�t$��Lf��C!-m��A�O:�OO$_�6_H_Z_l_�t*cgabl�Om���S!<m��Q�_:�
_�_ �_oo0oo)(Ӂ/�_�_���_�o�o�o�o��o�O@haul1�l�2r xm�<qC:��op�������Repla�W�fUȼ2�:�.�_4�F�X�j�|�m�$ %���o�������#��� 
��.�@���d���ŏ ׏����П����U� *�y�����r������� ��	�q��?�߯c�8� J�\�n���ϯ����� ڿ)����"�4�Fϕ� jϹ�˿��������� ���[�0�ϑ�fߵ� �ߜ߮�����!���E� W�,�{�P�b�t��� �߼�����A��(� :�L�^��������� ����� $s�H ������q���� �9]o�Vh z���U�#� G/./@/R/d/��/ �/��//�/�/?? *?y/N?�/�/�?�/�? �?�?�?�???Oc?u? JO�?nO�O�O�O�O+J�r	 H�O�O__ 6M2_@OBE:_p_>_P_ �_�_�_�_�_ o�_�_ oHoo(oZo�o^opo �o�o�o�o�o �o �:z �bA?� ; @�q _� ��Fw�� �Hw* �** @q >v�p2T�f�x�:���8����ҏ��eO^C 7�Տ#�5�G�	�k�}� ��ُ���c����� W��C�U�g���ß)� ����ӯ���	��-� w�����9�������m�@Ͽ��=�O�E	A��$MR_HIS�T 2�>uN��� 
 \�$Force �sensor c�heck  12�34567890�q�3����ß�߉N}SB� �-319.8 h�ours RUN� 9.�Y�!1s�t cleani�ng of co�nt. ventilation0�P�ϖϨ�-�Y����mech��cal�i�%Ό4��o�oDN�t��95���1����rollAeh�+�=�O��Y��Basic q�uarterly ߒߤ߶�
O4�F�� (�����b�t��� ��������M�_�����:�����p���:�S�KCFMAP  ]>uQ��r�5�������ON�REL  .��3���EXCFEN��:
��Q�FNCXJJOG_OVLIM8dN�\� ��KEY8�=�_PAN7�P���������SFSPDTYP8xC��SIG�:>��T1MOT�G���_CE_GRoP 1�>u\�D�����/� ���/�/U// y/0/n/�/f/�/�/�/ 	?�/???�/c??\? �?P?�?�?�?�?�?O�)OOMO,���QZ_�EDIT5 )T�COM_CFG 1���[�O�O�O� 
�ASI ��y3�
__+[_O_��>O�_bH�T_ARC_U�քT_MN_M�ODE5�	U?AP_CPL�_g�NOCHECK {?�� �� o.o@oRodovo�o �o�o�o�o�o�o�*!NO_WAI�T_L4~GiNTƑA���EUwT_7ERRs2���3���ƱJ�����X>_)��|MO�s��}�x:EB�  B4�  �r�x���8�?����� |�~�rPARAM�r]�����r_��:H5�5�G� =  r�b�t�s�X����� �������֟�0��:G�b�t�����S�UM_RSPAC�E�����Aѯۤ�$?ODRDSP�S7�cOFFSET_�CARt@�_�DI�S��PEN_FILE:�7�AF��PTION_IO���q�M_PRGw %��%$*�����M�WORK ��yf ���춍���� � ɂ������	 ч�����It���RG_DSBL'  ��C�{u���RIENTTO�7 ��Cn�A ��UT_SIM_EDy���V�?LCT ��}{Bx �٭��_PEX�P�=��RAT�W d�c��UP )���`���e�w�X]ߛߩ��$�2r��L6(L?}���	l d�� ����&�8�J�\�n� �������������@�"�4�F�X���2�� ��������������*�<w�Tfx �������J` �DT��Tz�Pg�� ����/"/4/F/ X/j/|/�/�/�/�� �/�/??0?B?T?f? x?�?�?�?�?�?�?�? �/�/,O>OPObOtO�O �O�O�O�O�O�O__`(_:_��O*��y_�]2ӆ��_�^�_�_ �W^]^]��/ooSog��Hgrohozo�o�o �o�o�oF`�#|G`A�  9y�����OK�1�k������<o�EA�nq? @D�  �q��4��nq?��C��s�q|1� ;�	l���	 |�Q�s<�r�q>��u
���qF`H<zH~��H3k7GL��zHpG��99l7�k_B�T�F`SC4��k�H���t���-�:����k������s��� � �ሏ����EeBVT���dZ�џ���ڏ ���q-�Fk�y�{jFbU���n@}6�  ����z�Fo��;�	'�� � ��I� �  �:p܋=���ڟ웆�@���B�,�D��B���g�:�N����  '|���g���B��p�BӀC�׏����@  #��Bu�&�ee^�^^މB:p 2���>�m�6p�Z���Dz?o}�܏�������׿������Ǒ��� ~f�  � �M�z��*�?�ff�_8�J�ܿ 3pϑ�ñ8�Чϵʖq.·�	(����P���'��s��tL�>��/�;�C�d;��.<���<�g�<F+<L ��^oiΚr�d@��r6p?fff�?�?&��;�@���@x��@��N�@���@T싶�Z���ћtމ �u�߈w	�x��ti�>� )�b�M��q����� ��������:�%�^��������W����E��  G�aF�� Fk��������� 1U@yd�� ����q��	�� {�A��h����D�a��ird��A{�/w/J/5/n/vA�A���":t�/ C�^/�/Z/ ލ?����/�/1??���Wҵ���g��pE�! ~1�?04�0
1ή1@IӀ��B���WB]�NB2��(A��@��u\?��������������b�0�|�uR����
�>��ؽ��B�u*C��$��)`�? ����GC#����rAU�����1�eG���I��mH�� I�:�I�6[Fߍ��C4OI���J�:\IT��H
~QF��y�Ol@�*J��/ I8Y�I���KFjʻC ��-?�O�O__>_)_ b_M_�_�_�_�_�_�_ �_o�_(oo%o^oIo �omo�o�o�o�o�o  �o$H3lW� {������� 2��V�h�S���w��� ��ԏ�������.�� R�=�v�a�������П ����ߟ��<�'�`� K�]���������ޯɯ���&�8�#�\��3(�J���3:a���9���J�3��c4������������1�����ڿ��1����e���14 �{2�2�r�`ϖτ�(�Ϩ��%PR�P���!�h�!�K�6�o��)����u�|ߵ� �����������3�� W�B�{�f�4���������d�A����!�� 1�3�E�{�i��������������  2 �Ef�7Fb�7���6B�!�!� C9� �� �0@�/`r@������#x�@�+=�3?, TV�8v��0�0���0�.
  D�����// %/7/I/[/m//�/�:� ��ֻ�G����$PARAM�_MENU ?�2�� � DEFP�ULSE�+	W�AITTMOUT��+RCV? �SHELL_W�RK.$CUR_oSTYL� 4<�OPTJJ?PTB�_?Y2C/?R_DECSN 0�Ű<�?�? �?�?�?OO?O:OLO�^O�O�O�O�O�O�!S�SREL_ID � .�����EUS�E_PROG �%�*%�O0_�CCC�R0�B���#CW_H�OST !�*!HT�_=ZT��O_�S�h_zQ�S�_<[_TGIME
2�FXU� ?GDEBUG�@�+��CGINP_FLgMSKo5iTRDo�5gPGAb` %l��tkCHCo4hTY+PE�,� �O�O �o#0Bkfx �������� �C�>�P�b������� ��ӏΏ�����(��:�c�^�p�����7eW�ORD ?	�+
? 	RSc`��/PNS��C4�sJOv1��TE�P�COL�է�2�Z�gLP 3������OjTRACEC�TL 1�2���! ��a �Қ�q�DT� Q�2�Ǡ���D � ��:�ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ�@����������� 6�H�Z�l�~ߐߢ�$� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� �������Щ *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 Fl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� x�N�߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�?��?�?�9�$PGT�RACELEN � �1  ����0��6_�UP �����A@�1�����1_CFG ��E�3�1
@�
<D�0<DZO<C�0�uO$BDEFSPD� �/L�1�0���0H_CONF�IG �E�3� �0�0d�D�&�2 �1�APpDsAl�A�0��0IN'@?TRL �/MOA�8pEQPE�E��G�A<D�AIWLID(C�/M	bT�GRP 1ýI� l�1B � �����1A��33FC� F8� E�� @eN	�A�AsA�Y�Y�A�@?� 	 vO�Fg�_ ´8cokB;`baBo,o>oxobo��o�1>о�?B�/�o�o~�o =%<��
 C@yd��"�������  Dz@�I�@A0�q� � ������ˏ���ڏ� ��7�"�4�m�X���|����Ú)ґ
V7�.10beta1�HF @�����Aq��Q�  �?� �B���P�p �C��~&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@p���f������ҡr�R�ܣ�Rљ����1�i�������t<B!CeQKNO?W_M  lE7F�bTSV ĽJ�BoC_�b�t��������������1�]aSM��SŽK ���	�NB�0����ĿK���-�bb��A�RP���`�0�Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1=�K
 4MU�iǨj� K�]�oߠ� �ߥ߷�������2�� #�h�G�Y��}������
������,�2r7�I��1�<t�H��P3^�p�����,�A4��������,�5(:,�6Wi{�,�7����,��8�!3,�MA�D�6 F,�OV_LD  KD��xO.�PARNUM�  �MC/%�S+CH� E
9'!8G)�3Y%UPD/���E�/P�_CMP_0��0@�0'7E�$�ER_CHK�%05H�&�/�+RS����bQ_MO�+?=5_�'?O�_RES_G6��:�I�o�?�?�? �?O�?O7O*O[ONO OrO�O�O�{4]��<�?�Oz5���O__ |3 #_B_G_|3V b_ �_�_|3� �_�_�_|3 � �_�_o|3Oo>o<Co|2V 1�:�k1�!�@c?�=2T?HR_INRc0i!�}�o5d�fMASS6�o Z�gMN�o�c�MON_QUEUE �:�"�j0��UO�N� U1Nv�+DpENDFqd?`y�EXEo`u� BE�npPAsOPTIO�Mwm;DpPROGR�AM %$z%�Cp}o(/BrTASK�_I��~OCFG� �$��K�D�ATA��T���j12/ď֏��� ���+�=�O�a�����������͟��INFO�͘��3t��!� 3�E�W�i�{������� ïկ�����/�A�@S�e�w�����Θ�a '��FJ�a K_N���T��˶ENB�g ڽw1��2��G�N�2�ڻ P(O�=���]�ϸ�@���v� ��u�uɡdƷ_E?DIT �T���|��G�WERFL�x��c)�RGADJ {Ҷ�A�  $Ձ?j00��a�Dqձ���5�?�$�ʨ�<u�)%e��0����FӨ�2�R��+	H;pl�G�b_�u>�pAod�t$��*�/� **:�j0�$�@�5AY�T���^��q�� �b~�L��\�n��� ������������� 4�F�t�j�|������� ������bLB T�x����: ��$,�Pb ���/���� /~/(/:/h/^/p/�/ �/�/�/�/�/V? ?? @?6?H?�?l?~?�?�? �?.O�?�?OO O�O DOVO�OzO�O_�O�O �O�O�Or__._\_R_ d_�_�_�_�_�_�_�f	g�io�pWo�o{d� �o�~o�ozoB�PREF �R��p�p
�IOR�ITY�w[���M�PDSP�q��pwU�T6����ODUC-T3�����;OG��_TG��8���ʯrTOENT �1׶� (!?AF_INE�p,�~7�!tcp7�>_�!udN���?!icmv���֯rXYK�ض���q)� ,�����p��&�	��R�9� v�]�o�����П����@��*��N�`�*�s�K��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE �R��:�w!d��连�2s�9Ks���PORT_N�UM�s�p����_CARTRE�P{p�Ω�SKST�A�w d�LGS6)�ݶ��tӁp�Unothin�g�������{��T?EMP ޾y���'e��_a_seiban�o\��ol� ��}߶ߡ��������� "���X�C�|�g�� ������������	� B�-�f�Q���u����� ��������,< bM�q��������(L�VOERSIyp�w}� disab�ledWSAVE� ߾z	26�00H768S?�!ؿ����/C 	5(�r)og+^/y�e{/�/�/�/�/�*�,/? �p���]_�p 1�Ћ� �����W�h?z?�W*pURGE«�B�p}vgu,�WFF�0DO�vƲ�vW%���4(�C�WRUP_�DELAY ��\κ5R_HOT �%Nf�q׿GO�5R_NORMAL&H��r6O�OZGSEMI�jO�O�O(qQSKI%PF3��W3x=_ 98_J_\_]�_�_{_ �_�_�_�_�_�_	o/o AoSoowoeo�o�o�o �o�o�o�o+= aOq����� ���'��7�]�K��������)E�$RAF{���K/�zĀÁ�_PARAM�A3���K @.�@�`�61�2C<��y��C�6$�B�ÀBTIF�4`�R�CVTMOUu�vc��ÀDCRF3}��I �+Q�5
=ޅ5���3�1.mU_ � �e�W�B=��1�\�k_-_��yS;�Cd;���.<߈<��g�<F+<L����Ѱ��d�u� L�������ϯ�����)�;�M�_���RD�IO_TYPE � M=U�k�EFP�OS1 1�\�
 x4/����� +�$/<��$υ�pϩ� D���h��ό��'��� ���o�
ߓ�.ߤ�R� ��������5���Y� ��i��*�<�v���r� ��������U�@�y� ���8���\������������?��c����2 1�KԿX��T�x��3 1����nY�>S4 1�'9�K�/�'/�S5 1���/�/��/�/:/S6 1� Q/c/u/�/-??Q?�/S7 1��/�/
?�D?�?�?�?d?S8 1�{?�?�?�?WOBO�{O�?SMASK �1L��O�D�GX�NO���F&�^��M�OTEZ�Ż��Q_�ǁ�%]pA݂��P?L_RANG!Q]��_QOWER ��ŵ�P1VSM_D�RYPRG %�ź%"O�_�UTAR�T �^�ZUME_PRO�_�_4o���_EXEC_E�NB  J�e�GSPD`O`WhՅjbgTDBro�jRM�o��hINGVERS�ION Ź�#o�)I_AIR7PURhP �O(.�MMT_�@T�P#_�ÀOBOT_I/SOLC�NTV@Az'qhuNAME�l���o�JOB_OR�D_NUM ?��X#qH7�68  j1Zc�@�r�rV��s��r�?��r?�r�pÀP?C_TIMEu�a��xÀS232>R1��� LT�EACH PEN�DANw�:GX��!O Main�tenance /Consj2�����"��No UseB�׏������p1�C�y�V�NPO�P\@�YQ�cS�oCH_L`�%^� �	ő��!U�D1:럒�R�@VGAIL�q@�Ӏ�J��QSPACE1 ;2�ż ��YR s�i�@Ct�YRԀ'{~��8�?�� ˯����"���7�2� c�u�����G���߯ѿ 򿵿�(��u�AC� c�u�����Ͻ�߿�� �ϵ��(��=�_�q� �ϕ�C߹������߱� �$��9�[�m�ߑ� ��Q������߭��� � ��	�W�i�{���M� ������5���. S�e�w�����I���� ���*?a s��E���� �/&//;/]o� �����/2/�/? "?�/7?Y/k/}/�/�/ O?�/�/�?�?�?O0O�OKA��*SY�PpM*�8.30�261 yB5/2�1/2018 gA �WPfG|�H��_TX`� !$�COMME��$USAp �$ENABLE=DԀ$INN`QpgIOR�B�@RY�E?_SIGN_�`�A�P�AIT�C�BWR�K�BD<�_TYP<�CRINDXS�@�W�@%VFRI{�_�GRPԀ$UF�RAM�rSRTOO}L\VMYHOL�A�$LENGTH�_VTEBTIRS�T�T  $S�ECLP�XUFIN�V_POS�@�$MARGI�A�$WAIT�`�ZX�2�\�VG2�GG1��AI�@�S�Q	g�`_�WR�BNO_USE�_DI�BuQ_RE�Q�BC�C]S$CUR_TCQP�R"a�^f �GP_ST�ATUS�A @� �A3`�BLk�HE$zc1�h�P@���@}_�FX �@�E_MLT_CTf�CH_�J�`CO�@�OL�E�CGQQ$�W�@w�b#tDE�ADLOCKuD�ELAY_CNT��a3qGt�a$wf _2 R1[�1$X<�2[2�{3[3$Zwy�q%Y�y�q`%V�@�c�@�b$V�`�RV�UV3oh>b�@ � �d�0ar'MSKJ�LgWaZ��C`NRK�PS_RATE�0$���S
`�Q�TAC��PRDH���e�S*��a4�At�0�DG�A 0�P��flp bquS2�ppI�#`
`�P �
�S\`  }�A�R_ENBQ� �$RUN?NER_AXI�<`�ALPL�Q�RU�TH�ICQ$FLI�P7��DTFERE�N��R�IF_CH�SU�IW��%V)�G!1����$PřA�Q�P�ݖ_JF�PR�_P�	�RV_D�ATA�A  {$�ETIM����$VALU$��	�OP_  � �A  2� �SC*��	� �$ITPa_!�SQ]PNPOU}��o�TOTL�o�DS}P��JOGLIb�N�PE_PKpc�Of�ji��PX]PTAS��$KEPT_M#IR��¤"`M�b�APq�aE�@�y�`q�g@١c�q�PG��BRK6�x���L�I��  ?�SJ�q��P�ADEz�ܠBS{OCz�MOTNv�DUMMY16Ӂ�$SV�`DE_�OP��SFSPDO_OVR
���@�LD����OR��T-P8�LE��F����6��OV��SF��F����bF�d�ƣ&c)��fQc�LCHDLY>��RECOV���`���W�PM��gŢ�R�O������_F�?�� @v�S �NVE�R�@�`OFS�PC,�CSWDٱc�ձ��X�B����TRG�š��`E_FDO��MOB_CM}���B���BLQ�¢	�Q�̄V�za�BUP�g��G
��AM���@`K�̊�e�_M!�d�AMxf�Q��T$CA����DF���HBKXd�v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�3�A��ATIO�0��͠��US����WaAB��R+c�`tá`xDؾA��_AUXw�?SUBCPUP���S�`����3Եжc���3�FLA�B�HW_Cwp"�Ns&�]s�Aa��$UNI�TS�M�F�ATT�RIz�Z�CYC=L�CNECA����FLTR_2_F�I��TARTUP`Jp����A��LP�������_SCT*cF�_F�F_P���b�FqS��+�K�CHA/Q���*�d�RSD���Q����Q���_T�H�PROr���հE#MPJ���G�T�� �Q�DI��@y�RAILAC4/�bMX�LOf�xS��ځ���拁���+PR#�S`app��C� 	��F�UNC���RIN�`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ng�DAQ�B�rkL�D�र&q�M�K���TI���j���$�@RIA_S�W��AF��Pñ�#��%%�p9r1��MsOIQ���DF_~P�(�PD"LM-�F�A�PHRDY�DORG�H; _QP�>s%MULSE~Pz�T��*�� J��Jײ���FAN_AL�MLVG��!WRN�%HARDP��Uc�O�� K2$SHADOW]�kp�a02���� STOf�+�_,^�w�AU{`R��eP_SBR�z5����:F�� �3MPINF?�\�4��3gREGV/1DG�b+cVm �C�CFL(��?�DAiP��ҌZ`�� �����Z�	� �P(Q$�A�$Z�Q V�@�[�
o� ��EG��o���kAAR���㌵�2�axG��AXEROB��RED���W�QD�_�Mh�S�YA��AF��FS�GW�RI�P~F&�STRP����E�˰EH�)�$�D�a\2kPB6P��t=V��Dv�OTO�19)���ARYL�tR0�v�3���FI&�ͣ?$LINKb!\�J�Q�_3S���E���QXYZ2�Z5N�VOFF���R�RJ�XxPB��d0s�G�cFI�03g��������_J ��'�ɲ�S&qR0LTV[6���aTBja�"�b�C���DU�F7.�TUR� X��eĂQ�2XP�ЊgFL��E���x@�`�U9Z8����� 1	)�K��Mw��F9��劂����ORQj��G;W3���#�Ґd ���uz����1�tOVE�q_�M��ё?C�uEC �uKB�v'0�x-�wH� �t���& `��qڠ �B�ё�u�q�wh�EC�h����ER��K	B�EP����AT�K�6e9e�W����AXs�'��v�/� �R ����!�� � �P��`��`�3p�Yp�1�p�� ��  �� (�� 8�� H��  X�� h�� x�� ����ޙ�DEBU�$�%3�I��·RAB����ٱ�sV��� 
d�J、��@� ��������Q���a�� �a��3q��Yq+$�`%"\<�cLAB0b�u�'�GRO���b<��B_s��"Tҳ *`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθ0uݸ��PNT0��?�SERVE �Z@� $`EAV�!�PO����nP�!�P@�$!Y@ � $>�TRQ"�b
=��BG�K�%"�2\��� _ � l��5�D6ER)RVb(�I��V0`;�N��TOQ:�7�L�@P
�R��e G�%�Q��� <�50F� ,h�`�z�>�RA�? 2 d!�����S�  M��p0xU ����OCuG��  ��CO�UNT6Q��FZN�_CFGF� 4#��6��TG4�_�=������Î�VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@H�EL�0��� 5b`B_BASN��RSR�6�C�SH����1�Ǌ�2���3��4��5��6ʭ�7��8��}�ROaO����P�PNLEAƭcAB)ë ��AC-Ku�INO�T��(B�$UR0� =�_P�U��!0��OU+�P�d�8j��� V��T�PFWD_KAR���� ��RE(ĉ P��P�>QUE�:RAO�p�`r0P1I� �x�j�P�f��6�QSCEM��0��� A��7STYL�SO j�DIX�&�����S!�_TMCMANR�Q��PENDIt�$KEYSWIT�CH���kHE��`BEATM83PE{@LE��>]���U��F��SpD_O_HOM# O�6@�EF�pPRaB(�A#PY�C� O�!���OV_M|b<0 �IOCM�dFQ�'�h�HKYA �D�Q�7��UF2��M����p�cFORC.�3WAR�"��k��OM|@  @�S�#o0U)SP�@1*�2&3&4E��*T�O��L���8OUNLOv�D4K$�EDU1  �S�Y�HDDNF� �M�BLOB  �p�SNPX_;AS�� 0@�0|��81$SIZ�1�$VA{���MU/LTIP-��# �A� � A$��� /4`�BS���0�C���&FRIF�BO�S���3� N=F�ODBUP߰��%@3;9(����Z@� x��SI��TE�s�r�cSGL�1T�Rp&�Н3B��@�0OSTMTq�3Pg@�VBW�p�4SHO�W�5@�SV��_�G�� 3p$PC�J�PИ���FB�PHSP AW�EP@�VD�0WC� ���A00��PB �XG XG XG$ XG5�VI6VI7VI8VI9
VIAVIBVI�XG�YF�0XGFVH��XbIU1oI1|I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1Y1Y2UI2bIU2oI2|I2�I2�I@�`�X�I2p�X�I2�IU2�I2�I2�I2Y�2Y�p�hbI3oI3�|I3�I3�I3�I3��I3�I3�I3�I3��I3�I3�I3Y3�Y4�i4bI4oI4�|I4�I4�I4�I4��I4�I4�I4�I4��I4�I4�I4Y4�Y5�i5bI5oI5�|I5�I5�I5�I5��I5�I5�I5�I5��I5�I5�I5Y5�Y6�i6bI6oI6�|I6�I6�I6�I6��I6�I6�I6�I6��I6�I6�I6Y6�Y7�i7bI7oI7�|I7�I7�I7�I7��I7�I7�I7�I7��I7�I7�I7Y7�T�VP� UD�y"ՠ��
<A62���t�R��CM)D� ��M5�Rv�]��Q_h�R���e�8���<�YSL���  � �%\2�׀+4�'��W�BVALU��b��'���=FH�ID_L����HI��I���LE1_��㴦�$0C��SAC�! h ��VE_BLC�K��1%�D_CPU5ɧ 5ɛ ������C�� ��R "? � PWj��l#0��LA�1SB���ì���RUN_FLG�Ś����ĳ ����������H���м����TBC2��#/ � @ B��e ��S�8=�FTD	C����V���3dՆQ�THF�����R��L�ESERVE9��F��3�2�E�|�Н�X -$��LEN9��F��f�cRA��W"G�W_5��b�1��д2�MO$-�T%S60U�Ik�0�`ܱF����[�DEk�21LACEi0�CqCS#0�� _MA� pj��z��TCV����z�T�������.B i�'A�z�'AJh�#E�M5���J��@@i�V�z���2Q �0&@�o�h��JK��VK�9��{���щ�J0l����JJ��JJ��AAL���������e4��5�ӕ N1��P����.�LD�_�1�
�CF�"% =`�GROU���1��AN4�C�#m R�EQUIR��E�BU�#��6�$Tk�2$���zя �#�& \�APP�R� C� 0�
$O�PEN�CLOSD�St��	i�
�.�&' �MfЩ�8��W"-_MG߱7�CB@�A���BB{RK@NOLD@>�0RTMO_5ӆ$p1J��P��� ������������6��1�@ %�Р�#�(� ������'��+#PATH''@!6#@!��<#� � '��1SCaA���6IN�ңUCJ�[1� C0@UM�(Y ��#�"������*���*��� PAYwLOA~J2LؠOR_AN^�3L���91�)1AR_F�2LSHg2B4LO�4�!F7�#T7�#ACRL_�%�0�'�$r��H��.�$HA^�2FLEX��J!�) P�2�D��߽���0��* :����z�FG]D��`��z���%�F1]A �E�G4�F�X�j�|���BE���������� ��(��X�T*�A���@�XI�[�m�\At�T$g�QX<�=��2TX ���emX���������� ��������+	�J>+ �-�K]o|�٠AT�F�4�CELFPѪs�J� �*� JEmCTR��!�ATN�vzH�AND_VB.���1��$, $8`Fi2Av���SWu��-� $$M*0.�]W�l g��PZ����A��� 1����:AK��]AkAz��LN�]UDkDzPZ G���C�ST_K�lK�N}DY��� A���� 0��<7]A<7W1�'��d�@g`�P��������"Os"�. M�2D%"��H�����ASYMj%0��� j&-��-W1�/_ �{8� �$�����/�/�/�/ 3J<�:p9�/�89�D_VI��v����V_UN!I�ӛ��cD1J���� ╴�W<��n5Ŵ�w=�4��9��?�?<�uc$�4�3�%�H����/�j��0�DI�zuO��;�k�>S0 �`��I��A���#���@ģ���@���HQl� 1 � -/�ME.Qp��49�ơT}�PT�;pG �+ /� ����'��T�0 $DUMMY1���$PS_�@RF��@  G b�'FLA@ YP(c|��$GLB_TP� ŗ���9 P�q���2 X� z!ST�9�� SBRM M�21_V�T$S/V_ER*0O�p�Ӧ��CL����AGPOl��f�GL~�EW>��3 4H �$Y
rZrW@�x�A1+��A���"��"�U&�4� 8`NZ�"�$�GI�p}$&� �-� �Y�>�5 L�H {��}$F�E^��NEAR(PN�CyF��%PTANC�BΚ�JOG�@� �6Mp$JOIN�Twa' d�MSET.>�7  x�E��HQ�tpS{r��up>�8׼ �pU.Q?��� LOCK_FOxV06���BGLV�s�GLt�TEST_sXM� 3�EMP�����_�$U&@%�w`24� Y��5��2�d��3��C�E- ���� $KA�R�QM��TPDRqA)�����VECn@���IU��6��H=Ef�TOOL�C2�V�DRE IS3�ER6��@ACH� 7?Ox �Q��29Z�H I� � @$RAIL_�BOXEwa�R�OBO��?��HOWWAR�1�_�zROLMj��:q�w�jq� �@ O_=Fkp! d�l�>�9�� �R OB8B: �@�c�KOU�;�Һ�3ơ��r�q_�$PIP��N&`H�l�@���#@CORDED�d�p >f�fpO�� �< D ��OB⁴sd���Kӕи��qSYS�A�DR�qf��TCH�t� = ,8`E�No��1Ak�_{��-$CqKuPVWVA~��> �  �&��PREV_R�T�$EDIT�r&VSHWRkqP�֑ &R:�v�D���JA�$�a$HECAD�6�� �z#�KE:�E�CPSP]D�&JMP�L~�2�0R*P��?��1�%&I��S�rC�pN�E; �q�wTICKğC��MJq3�3HN��@ @� 1Gu��!_GPp6��0S3TY'"xLO��:��2l2?�A t 
�m G3%%$R!{�=:��S�`!$��w`����ճ���Pˠp6S�QU��E��u�TEsRC�0��TSUtB ����hw&`gw�Q)�pO����@�IZ��{��^�P�R�kюB1XPU����E_DO��, XuS�K~�AXI�@���UR�pGS�r � ^0�&��p_) ��ET�BPm��o���0Fo��0A|����Rԍ��a��S=R�Cl>@P� �b_�yUr��Y��yU�� yS��yS���UЇ�U�� �U���U�]��Ul[��Y�bXk�]Cm������YRSC�� 7D h�DS~0��fQ�SP���eATހ��A]0,2N�AD�DRES<B} S�HIF{s��_2C�H�p�I��=q�+TVsrI��E"����a�Ce�
��
��V8W�A��F \��qA��0l|\A@�rC��_B"R{zp�ҩq�T�XSCREE�Gzv��1TINA����t{����A�b?�H T1�ЂB��р��I��A��BE�y RRO������ B��Dv��UE4I �g��!p�S��RSM<]0�GUNEX(@~���j�S_S�ӆ��Á։񇣣�ACY�0�o 2H�pUE;��J�����@GMTJ��Lֱ�A��O	�/BBL_| W8��ЧK ��0s�OM���LE/r��� TO�!�s�RIGH��B�RD
�%qCKGR8л�TEX�@����WIDTH�� �Bh[�|�<��I_��}Hi� L 8K�B��_�!=r���R:�@_��Yґ��O6qJ�Mg0紐U��rh�Rm��LUMh��FpERVw �QP���`�N��&�/GEUR��FP)�M)� LP��(RE%@�a)ק�a�!��f ��5�6�7�8 Ǣ#B�É@���tP�f�W�S@M�U{SR&�O <�����U�Qs�FOC\)��PRI;Qm� �:���TRIP�Om�UN����Pv��0��f%��'���@��0 Q����AG �0T� �a>q�OS�%�RPo���8�R/�A�H�L�q4$����U¡�SU�g�p�¢p5��OFF���T�}�O�� G1R�����S�GUN��6�B�_SUB?���,�SRTN�`TUg2���mCOR| D�RAU�rPE�TZ�#'�VC�C��	3V AC?36MFB1f$c�{PG �W (#�.�ASTEM����L�0PE��T3G��X �\ ��MOV1Ez�<���AN�� ����M���LIM_X��2��2��7�,������ı�
��VF@�`E�+�~��04Y�F�IB�7���5S���_Rp� 2��� WİGp+@��}���P��3�Zx ���3���A�rݠCZ�DRID�����Vy08�90� D~e�MY_UBYd�@��6��@��!��X��P_S��3��mL�KBM,�$+07DEY(#EX`������UM_MU� X����ȀUS�� �z��G0`PACI�� �а@��:��:,�:����RE/�3qL�+���:[��TA�RG��P�r��R<�\ d`��A���$�	��AR��SWH2 ��-��@Oz��%qA7p�yREU�Uh�01�,�HK�2]g0�qP� N�� �EAM0GWORx���MRCV3�W^ ���O�0M��C�s	���|�REF_���x(�+T � ���������3_RCH4(a �P�І�hrj�NA�5��0�_ ��2����L@4��n�@@OU~7w�p6���Z��a2[ư�RE�p�@;0\��c�a'2K�@SUL���]��C��0�^��� NT��L�3��@(6I�(6q�(3� L��@Q5��Q5I�]7q�}�)Tg`4D`�0.`0ПAP_HUC�5S]A��CMPz�F�6(�5�5�0_�aR��a��1I\!X�9��G�FS��ad †M��0p�UF_`x��B� �ʼ,RO���Q��'����UR�3GR�`.�3IDp���)�D�;��A��~�IN��H{D���V@��J���S͓UW�mi=�����TYL�O*�5����bot +�cPA�{ �cCACH� vR�UvQ��Y��p�#�CF�I0sFR�XT8���Vn+$HO����P!A3�XBf�(01 ���$�`VPy� �^b_SZ313he6K3he12J�eh chlG�chWA�UMP�j���IMG9uPAyD�iiIMRE�$^�b_SIZ�$P�����0 ��ASYNB{UF��VRTD)u�5tqΓOLE_2�DJ�Qu5R��C��U���vPQuECCUlVEMV �U�r��WVIRC�aIuVTPG���rv1s��5qMPLAqa��v����0�cm� CKLAS�	�Q�"���d  �ѧ%ӑӠ@�}¾�$�Q���Ue A|�0!�rSr�T�# 0! �r�iI��ml�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f �� >֦3�@Sp�SgLOW>�RO��ACCE���!� 9��VR�#���p:���A1D�����PAV�j��� D����M_B8"���^�JMPG ���g:�#E$SSC@��x&�vPq��hݲ�vQS�`qVN��L;EXc�i T`�s�r���Q�FLD �DEsFI�3�0p2���:��VP2�V�j� �A��V|�4[`MV_PIs���t���A�@��F	I��|�Z��Ȥ����`�A���A��~�GAߥ�1 LOO��1 JC�B���Xc��^`TcP�LANE��R��1F@�c�����pr�M� [`�噴��S����f� ���Af��R�Aw�״t9U��pRKE��d�VANC������ k���ϲϡ�wR_AA� l���2� ��p�#Hć�m h�@��O K�$����2��kЍ0OU&A�"eA�
p�pSK�T�M@FVIEM 2l� ��P=���n �<<��dK�UMM�YK1P��`D6T`ȡ�CU��#A�U��o $��T�IT�$PR�����OP���V�SHIF�r�p`J�Q���fOxE[$� _R�`UTc ����s��q������ G�"G�޵'�T�$��SCO{D7�CNT Q i�l�>a�-�a�;� a�H�a�V���1�+�2u1��D���� w � SMO�U�q��a�JQ���%��a_�R[�r�n׍*@LIQ�AA/`��XVR��s�n�T�L���ZABC��t�t�c�
L�Z�IP��u���LV�bcLn"���MPkCFx�v:�$��� ���DMY_L�N�������@y�w �Ђ(a�u� MCM��@CbcCART_��DPN� $J71D��=N�Gg0Sg0�BUXW|� ��UXEUL|ByX���	������x P	���m�YH�Db  y 80���0�EIGH�3n�?(�� H����$z a���|�����$B� �Kd'��_��L3�R�VS�F`���OVC�2'�$|�>P&���
q���5D�T�R�@ �Vc��SP9HX��!{ ,� �*<�$R�B2 �2 ���C!��  � V-L�b*c%g!)`+g"�`V*�,?8�?�V+�/ V.�/�/?�/�/V(7%3@/R/d/v/�/6?�/ �/�?�?�?O4OOION;4]?o?�?�?�?SO �?�?�O_�O0_Q_8_f_N;5zO�O�O�O�O p_�O_o8o�_MonoUo�oN;6�_�_�_�_ �_�oo%o4Uj�r�N;7�o�o�o �o�o� BQ�r�5� ��������N;8�� ���Ǐ=�_�n����R���ş��ڟN;G ;� џ�
����?���W�i� {�������ï�.��@�����A��dW� <�N�|�������Ŀֿ �ޯ���0�B�_� R�d�꿤϶������� ������*�L�^�� rτ�
������������&�8�J�l�~�; `ҟ @���@���ߩ��-��� �&�,���9�{��� ��a������������� ��A'Y�� �������a#1�
��N;�_MODE  ���S ��[�Y�B���
/\/�*	|/�/R4CWO�RK_AD�	�{�T1R  ����� �/� _INOTVAL�+$���R_OPTION�6 �q@V_�DATA_GRPg 27���D��P�/~?�/�?�9��? �?�?�?OO;O)OKO MO_O�O�O�O�O�O�O _�O_7_%_[_I__ m_�_�_�_�_�_�_�_ !ooEo3oioWoyo�o �o�o�o�o�o�o /eS�w�� �����+��O� =�s�a�������͏�� �ߏ��9�'�I�o��]�����$SAF�_DO_PULS�� �~������CAN_TIM������ SCR ��Ƙ�" 5�;#U!P"�1!��� �?E�W�i� {�����.�ïկ���X��'(~�T"2F���dR�I�Y��2�o+@a얿�����)�u��� k0ϴ���_ ��  �T� � �2�D�)�T D��Q�zό� �ϰ���������
�� .�@�R�d�v߈ߚ�/<V凷������߽��R�;��o �W�p��
�?t��Diz$�~ �0 � �T" 1!�������� ����������*�<� N�`�r����������� ����&8J\ n���������"4FX �� ࿁������ �/`4�=/O/a/s/ �/�/�/�/�/�/�!!/ �0޲k�ݵu�0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ ok $o6oHoZolo~o�o�o �o�o1/�o�o 2 DVhz�/5?�� ������&�8� J�\�n���������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u��� ���`Ò�ϯ ����)�;�M�_� q���������˿ݿ�� ����3� ����&2,��	12345678v��h!B!�U�h�Ch���0� �ϵ����������!� 3�9ѻ�\�n߀ߒߤ� �����������"�4� F�X�j�|�h�K߰��� ������
��.�@�R� d�v������������� ��*<N`r ������� &��J\n�� ������/"/ 4/F/X/j/|/;�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �/�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_�?L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o=_�o �o�o�o�o�o 2 DVhz�����h������u�o�.�@�R���Cz � B��   ����2&� � �_�
���  	�_�2�Տ���,�_�p������ďi�{�������ß ՟�����/�A�S� e�w���������N�� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�_�����<v�_��$SC�R_GRP 1
�� �� �t ��� ���	 ��������� �������_�����Ϝ)�a����&�DE� DW8���l��&�G�CR-3�5iA 9012�34567890���M-20��8~��CR35 ��F:�
��������������:֦�Ӧ��G���&������	���]�o����:���H���>�����������&���ݯ:��j����g�X�����B�t�����������A����  1@����@� (' ?�=��Ht�P�
��F@ F�`z�y����� � �$H���Gs^p��B� �7��/�0// -/f/Q/�/u/�/�/�/�8���P�� 7%?�����"?W?-2?<���]? H�1�?t�ȭ7�������?-4A, �&E@�<�I@G�B-1 3OZOlO-:HA�H�O�O.|O P�B(�B�O��O_��EL_DE�FAULT  ~���-0�SHOTSTR�#]JA7RMIPOWERFL  i�z/UYTWFDO$V� /URRVENT 1�����NU L!DU�M_EIP_-8��j!AF_IN�E#P�_-4!FT$�_->�_;o!��`o� �*o�o!RPC_MAIN�o�jh�vo�o�cVIS�oii��o!TMPpPU�Yd�k!
PMON_�PROXYl�Ve Z�2r��]f���!RDM_SR�V��Yg�O�!�R��k��Xh>���!%
�`M��\i����!RLSYNC��-98֏3�!gROS�_-<�4"���!
CE4pMT'COM���Vkn�˟{!	��CONS̟��Wl���!��WOASRC��Vm�vc�!��USBd��XnR���Noӯ��� ����!��E��i�0����WRVICE_�KL ?%�[ �(%SVCPR#G1��-:Ƶ2ܿ�"˰3�	�˰4,�1�"˰5T�Y�˰6|ρ�˰7�ϩ�˰�����	9����ȴf�!�˱ οI�˱��q�˱ϙ� ˱F���˱n���˱�� �˱��9�˱��a�˱ ߉��7߱��_��� �����)���� Q����y��'��� O����w����� ����˰��İd �c������ =(as^�� ����/�/9/ $/]/H/�/l/�/�/�/ �/�/�/�/#??G?2? k?V?}?�?�?�?�?�? �?O�?1OCO.OgORO �OvO�O�O�O�O�O	_��O-_��_DEV ��Y�MC�:5X�`GTG�RP 2SV5P���bx 	� 
+ ,�P5P5_�_ �T�_�_�_o�_'o9o  o]oDo�ohozo�o�o �o�o�o�o5{�_ g������ ����?�&�c�u� \�������Ϗ���J \)���M�4�q���j� ����˟ݟğ��%� ��[�B��f����� �ٯ�������3�� W�i�P���t���ÿ�� �ο���A�(�e� L�ί��RϿ��ϸ��� ��� ��O�6�s�Z� �ߩߐ��ߴ������ '�~ϐ�]���h�� ������������5� �Y�@�R���v����� ����@�	��?& cu\����� ���;M4q X�������/ �%//I/[/B//f/ �/�/�/�/�/�/�/�/ 3??W?�L?�?D?�? �?�?�?�?O�?/OAO (OeOLO�O�O�O�O�O��O�O�O_"Ud ��NLy�6 *� 		S=>���+c"_VU@Tn_Y_B����B�2�7J�j~Q´~_g_��_�Q%JOGGGING�_�^7T(?VjZ�Rf��Y���/e�_%o7e�Tt�]/o�o{m�_�o �m?Qi�o�o;)Kq%��o�}o s������9� {`��)���%���ɏ ���ۏ�S�8�w�� k�Y���}���ş��� +��O�ٟC�1�g�U� ��y�������'��� �	�?�-�c�Q���ɯ ����w���s���� ;�)�_ϡ���ſOϹ� ����������7�y� ^ߝ�'ߑ�ߵߣ��� �����Q�6�u���i� W��{������=� �M���A�/�e�S��� w������������ =+aO���� ��u���9 ']���M�� ����/5/w\/ �%/�/}/�/�/�/�/ �/=/"?4?�/?�/U? �?y?�?�?�??�?9? �?-OO=O?OQO�OuO �O�?�OO�O_�O)_ _9_;_M_�_�O�_�O s_�_�_o�_%oo5o �_�_�o�_[o�o�o�o �o�o�o!coH�o {������ ; �_�S�A�w�e� ������я���7��� +��O�=�s�a����� �П�����'�� K�9�o�������_��� [�ɯ���#��G��� n���7���������ſ ����a�Fυ��y� gϝϋϭϯ�����9� �]���Q�?�u�cߙ� �ߩ���%���5���)� �M�;�q�_���߼� �߅������%��I� 7�m������]����� ������!E��l ��5������ �_D�we �����%
// ���=/s/a/�/�/ �/��/!/�/??%? '?9?o?]?�?�/�?�/ �?�?�?O�?!O#O5O kO�?�O�?[O�O�O�O �O_�O_sO�Oj_�O C_�_�_�_�_�_�_	o K_0oo_�_co�_so�o �o�o�o�o#oGo�o ;)_Mo��� �o����7�%� [�I�k��������� �ُ���3�!�W��� ~���G�i�C����՟ ���/�q�V������ w��������ѯ�I� .�m���a�O���s��� ����߿!��E�Ͽ9� '�]�Kρ�oϑ��� ��Ϸ����5�#�Y� G�}߿Ϥ���m���i� �����1��U��|� ��E���������	� ��-�o�T������u� ����������G�, k���_M�q�� �����% [Im���	 ���//!/W/E/ {/��/�k/�/�/�/ �/	???S?�/z?�/ C?�?�?�?�?�?�?O [?�?RO�?+O�OsO�O �O�O�O�O3O_WO�O K_�O[_�_o_�_�_�_ _�_/_�_#ooGo5o Wo}oko�o�_�oo�o �o�oC1Sy �o��oi���� �	�?��f�x�/�Q� +���Ϗ�����Y� >�}��q�_������� ˟���1��U�ߟI� 7�m�[�}����ǯ	� �-���!��E�3�i� W�y�ϯ��ƿ����� ���A�/�eϧ��� ˿UϿ�Q�������� �=��dߣ�-ߗ߅� �ߩ��������W�<� {��o�]����� ����/��S���G�5� k�Y���}��������� ������C1gU ������{��� �	?-c��� S������/ ;/}b/�+/�/�/�/ �/�/�/�/C/i/:?y/ ?m?[?�??�?�?�? ? O??�?3O�?COiO WO�O{O�O�?�OO�O _�O/__?_e_S_�_ �O�_�Oy_�_�_o�_ +oo;oao�_�o�_Qo �o�o�o�o�o'io N`9��� ���A&�e�Y� G�i�k�}�����׏� ��=�Ǐ1��U�C�e� g�y����֟���	� ��-��Q�?�a���ݟ ��퟇��ϯ��)� �M���t���=���9� ��ݿ˿��%�g�L� ����mϣϑϳ��� ����?�$�c���W�E� {�iߟߍ߯������ ;���/��S�A�w�e� ������������� +��O�=�s������ c�����������' K��r��;��� ����#eJ� }k����� +Q"/a�U/C/y/ g/�/�/�//�/'/�/ ?�/+?Q???u?c?�? �/�?�/�?�?�?OO 'OMO;OqO�?�O�?aO �O�O�O�O__#_I_ �Op_�O9_�_�_�_�_ �_�_oQ_6oHo�_!o �_io�o�o�o�o�o)o Mo�oA/QSe�����%{,p��$SERV_M�AIL  +u�!���q�OUTP�UT�$�@��RV 2�v  $� (�q�}���SAVE7�(�TOP10 2W�� d 6 	*_�π(_����� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ�ݷ��YP��'�FZ�N_CFG N�u$�~���~�GRP 2��D� ,B   �A[�~�D;� B}\��  B4~��RB21��H7ELL��u���j�k�2�����%RSR�������
� C�.�g�Rߋ�v߈��� ������	���-�?�Q��  �_�%@Q���_���,p1����ޖ�g��2,pd����HKw 1�� �� E�@�R�d��������� ��������*<�e`r���OMM� �����FT?OV_ENB�_����HOW_REG�_UI�(�IMI_OFWDL� ��^�)WAIT� ��$V1�^�NwTIM����VA�_)_UNcIT����LC�TRYB�
�M�B_HDDN 2W� 2�:% 0 �pQ/�qL/^/�/�/��/�/�/�/�/�"!O�N_ALIAS k?e�	f�he� A?S?e?w?�:/?�?�? �?�?�?OO&O8OJO �?nO�O�O�O�OaO�O �O�O_"_�OF_X_j_ |_'_�_�_�_�_�_�_ oo0oBoTo�_xo�o �o�o�oko�o�o ,�oPbt�1� ������(�:� L�^�	���������ʏ u�� ��$�Ϗ5�Z� l�~���;���Ɵ؟� ���� �2�D�V�h�� ������¯ԯ���
� �.�ٯR�d�v����� E���п���ϱ�*� <�N�`�r�ϖϨϺ� ��w�����&�8��� \�n߀ߒߤ�O����� ������4�F�X�j� |�'���������� ��0�B���f�x��� ����Y������� ��>Pbt�� ����(: L�p����c �� //$/�H/Z/ l/~/)/�/�/�/�/�/��/? ?2?D?V?]3��$SMON_DE�FPRO ����1� *SYST�EM*0m6RECALL ?}9� ( �}9c�opy frs:�orderfil�.dat vir�t:\tmpba�ck\=>147�.87.149.�40:17680� 98 �6517�2]?O+M}0�2m?db:*.*�?�?� �?O�O�O8C4x�4:\HO�@ZOuAtO��O_)_ }5�Ea �O�OpF�O_�_�_�? �?XOsO�_o(o;O�_ _O�_o�o�o�OL_^_ �O�o$7_�o�om_ �o���_�_Po�_} � �3oEo�io��� ���o�oV�oy�
�� /Aҏe��+���� ��_�u����*�=� ؟a���������N� [�񏃯�&�9�ʯܯ o��������ɟR�� ��"�5�G��k��� �Ϡϳ�ůX��{�� �1�C���g��ϊߜ� ����ӿa�w߫��-� ?���c������� P�]��υ��(�;��� ��q����������T� �߁�$7�I���m� ������H�Z���}  3�E��i����1
<��Lout�put\test�_server.�pcC : o� �_6279142?4:3597y
/ /������aw+/�/ -?Z/cu/�/?*? �P�/�?�?�?; L?^?q�?O&O9/K/ �/o/O�O�O�/�/dO �/O_"_5?�?�?k? �O�_�_�?�?V_�?{_ oo�����_�o �o/OAOSO�_�_�o �O�O�o�O�o����$SNPX_A�SG 2�����q� �P 0 '%�R[1]@1.Y1��y?��s%� !��E�(�:�{�^��� ����Տ��ʏ��� A�$�e�H�Z���~��� џ����؟�+��5� a�D���h�z�����ů �ԯ���
�K�.�U� ��d�������ۿ��� ���5��*�k�N�u� �τ��ϨϺ������ 1��U�8�Jߋ�nߕ� �ߤ����������%� Q�4�u�X�j���� ���������;��E� q�T���x��������� ��%[>e �t������ !E(:{^� �����/�/ A/$/e/H/Z/�/~/�/ �/�/�/�/�/+??5? a?D?�?h?z?�?�?�? �?�?O�?
OKO.OUO �OdO�O�O�O�O�O�O _�O5__*_k_N_u_ �_�_�_�_�_�_�_o 1ooUo8oJo�ono�o��o�d�tPARAM� �u�q ��	��jP�d�9p�ht��pO�FT_KB_CF�G  �c�u�sO�PIN_SIM  �{vn���p�pRVQSTP/_DSBW~r"t|�HtSR Zy� � & R�OB195_SE�RV M����vTOP_ON_?ERR  uCy~8�PTN Zu�k�A4�R?ING_PR�D���`VCNT_GOP 2Zuq�!px 	r��ɍ����׏��wVD��RP' 1�i p�y ��K�]�o��������� ɟ۟����#�5�G� Y���}�������ůׯ �����F�C�U�g� y���������ӿ�� 	��-�?�Q�c�uχ� �ϫ����������� )�;�M�_�qߘߕߧ� ����������%�7� ^�[�m������� ������$�!�3�E�W� i�{������������� ��/ASew ������� +=Ovs�� �����//</ 9/K/]/o/�/�/�/�/ �/�/?�/?#?5?G? Y?k?}?�?�?�?�?�?��?�?OO)�PRG�_COUNT8vq�k�GuKBENB���FEMpC:t}O_UP�D 1�{T  
4O�B�O�O�O_ _!_3_\_W_i_{_�_ �_�_�_�_�_�_o4o /oAoSo|owo�o�o�o �o�o�o+T Oas����� ���,�'�9�K�t� o���������ɏۏ� ���#�L�G�Y�k��� ������ܟן���$� �1�C�l�g�y����� ����ӯ����	��D� ?�Q�c���������Կ Ͽ����)�;�d��_�q�=L_INFO� 1�E�@ �2@����������� ��B�  ?B4 �4*�@HYSDEBUGU@ʶ@���d�If�SP�_PASSUEB�?x�LOG  *���C��Qؑ��  ��A��U�D1:\��Uߦ�_MPC�ݵE&�8�A���V� �A�SAV !������ҶX���SVZ�T�EM_TIME �1"���@ 01@$X��X�E������$T1SVGgUNS�@VE'�E���ASK_OPTIONU@�E�A�A+�_DI��qOG��BC2_GRP �2#�I�����@��  C���<Ko�C�FG %z��� 1�����`��	� .>dO�s� ������* N9r]���� ���/�8/#/\/n/v$Y,�/Z/�/�/ H/�/?�/'??K?]� k?=�@0s?�?�?�?�? �?�?O�?OO)O_O MO�OqO�O�O�O�O�O _�O%__I_7_m_[_ }__�_�_�X� �_�_ oo/o�_SoAoco�o wo�o�o�o�o�o�o =+MOa�� �������9� '�]�K���o������� ��ɏ���#��_;�M� k�}��������ß� ן��1���U�C�y� g�������������� �	�?�-�c�Q�s��� �������Ͽ��� �)�_�Mσ�9��ϭ� ������m���#�I� 7�m�ߑ�_ߵߣ��� ��������!�W�E� {�i���������� ����A�/�e�S�u� w������������� +=O��sa�� �����9 ']Kmo��� ����#//3/Y/ G/}/k/�/�/�/�/�/ �/�/??C?��[?m? �?�?�?-?�?�?�?	O �?-O?OQOOuOcO�O �O�O�O�O�O�O__ ;_)___M_�_q_�_�_ �_�_�_o�_%oo5o 7oIoomo�oY?�o�o �o�o�o3!Ci W������ ���-�/�A�w�e� ���������я�� �=�+�a�O���s��� ����ߟ͟��o�-� K�]�o�ퟓ�����ɯ��צ��$TB�CSG_GRP �2&ץ��  �� 
 ?�  6�H�2� l�V���z���ƿ��������(�d׊E+�?�	 �HC���>���G����C�  �A�.�e�q�C��N>ǳ33��S�/]���Y��=Ȑ� C\�  Bȹ��B���>����P���KB�Y�z��L�H�0�$����J�\�n�����@�Ҿ����� ����=�Z�%�7��鈴�?3�����	�V3.00.�	�cr35��	*����
�������Ƈ� 3��4�  7 {�CT�v�,}��J2�)��������CFG +�ץ'� *�������I����.<
�<b M�q����� ��(L7p[ ������/ �6/!/Z/E/W/�/{/ �/�/�/�/.�H��/? ?�/L?7?\?�?m?�? �?�?�?�? OO$O�? HO3OlOWO|O�O��� �Oӯ�O�O�O!__E_ 3_i_W_�_{_�_�_�_ �_�_o�_/oo?oAo So�owo�o�o�o�o�o �o+O=s� E���Y���� �9�'�]�K�m����� ��u�Ǐɏۏ���5� G�Y�k�%���}����� ßşן���1��U� C�y�g�������ӯ�� ����	�+�-�?�u� c����������Ͽ� ��/�A�S�����q� �ϕϧ��������%� 7�I�[���mߣߑ� �������߷��3�!� W�E�{�i����� ��������A�/�e� S�u������������� ��+aO� s��e����� 'K9o]� ������#// G/5/k/}/�/�/[/�/ �/�/�/�/??C?1? g?U?�?y?�?�?�?�? �?	O�?-OOQO?OaO �OuO�O�O�O�O�O�O ___M_�e_w_�_ 3_�_�_�_�_�_oo 7o%o[omoo�oOo�o �o�o�o�o!3�o �oiW�{��� ����/��S�A� w�e�������я���� ���=�+�M�s�a� ��������ߟ�_	� ��_ן]�K���o��� ����ۯɯ���#�� �Y�G�}�k�����ſ ׿��������U� C�y�gϝϋ��ϯ��� �����	�?�-�c�Q� s�u߇߽߫������ ��)��9�_�M���� /����i������%� �I�7�m�[������� ������������E Wi{5���� ����A/e S�w����� /�+//O/=/_/a/ s/�/�/�/�/�/�/? '?��??Q?c??�?�? �?�?�?�?�?O�?5O GOYOkO)O�O}O�O�O��O�N  �@S� V_R�$T�BJOP_GRP� 2,�E�  ?�Vi	-R4S.;\��@�|u0{SPU �>��UT� @�@LR	 ��C� �Vf  �C���ULQLQ>�33�U�R�����U�Y?�@=�Z�C��P��ͥR�>�P  B��W$o�/gC��@g�d�Db�^����eeao�P&ff�e=��7LC/kaB� o�o�P��P�ef�b-C�p��^�g`�d�o�PL�Pt<�eVC\  �Q�@�'p�`�  �A�oL`�_wC�BrD�S�^��]�_�S�`<P�B��P�anaa`C�;�`L�w�aQo�xp�x�p:���XB$'tMP@�PCAHS��n���=�P𥅡�trd<M�g E�2pb����X�	� �1��)�W���c�� ����������󟭟�7�Q�;�I�w���;d��Vɡ�U	V3�.00RScr35QT*�QT�A��� E�'�E�i�FV#�F"wqF>���FZ� Fv�R�F�~MF����F���F��=�F���F�ъ�F��3F����F�{G
�GdG��G#
�D���E'
EMK�E���E����E�ۘE����E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F���vF�u�<#�_
<t���ٵ�=�_��V� �R�p�V9� ]E_STPARtp�H�FP*SHR\�ABL/E 1/;[%�S�G�� �W�G�BG�G� WQG�	G�E
G�GȖ�QG��G�G�ܱv�RD	I~�EQ�ϧϹ�������W�O_�q�{ߍߐ�߱���w�S]�CS  !ڄ���������� ��&�8�J�\�n��� ���������� ]\�`� ��	��(�:������
��.�@�w�NUoM  �EEQ�P	P ۰ܰw�_CFG 0���)r-PIMEBF_TTb��CSo�,GVERڳ-B,�R 11;[ 8I��R�@� �@&  ����� ��//)/;/M/_/ q/�/�/�/�/�/?�/ ?J?%?7?M?[?m?> �@�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_l�_�Y@cY�M�I_CHAN8 �c cDBGLVĂ�:cX�	`ET�HERAD ?*f�\`��?�_�uo�oQ�	`ROUT6V!	
!�d�o~�lSNMASKQh|cba255.u�ߣ'9ߣY�OOLOFS_DIb���U;iORQCT�RL 2		�Ϸ~T����� #�5�G�Y�k�}����� ��ŏ׏�����.���R�V�PE_DE�TAI/h|zPGL�_CONFIG �8�	���/�cell/$CID$/grp1V�@̟ޟ����Ӏ�o ?�Q�c�u�����(��� ϯ������;�M� _�q�����$�6�˿ݿ ���%ϴ�I�[�m� ϑϣ�2��������� �!߰���W�i�{ߍ��߱�%}F�������/�A�C�i�H� Eߞ����������?� �.�@�R�d�v���� ������������* <N`r��� ����&8J \n��!��� ��/�4/F/X/j/ |/�//�/�/�/�/�/ ??�/B?T?f?x?�? �?+?�?�?�?�?OO �?>OPObOtO�O�O�O����User� View ��}�}1234567890�O�O�O_#_`5_=T�P��]_���I2�I:O�_�_�_�_�_�_X_j_�B3�_GoYo�ko}o�o�o o�op^4 6o�o1CU�ovp^5�o���� �	�h*�p^6�c� u����������ޏp^7R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3� �OM�_�q��������y  e��Yz���	�� -�?�Q���uχϙ�俀����������>�� e�5i��c�u߇ߙ߫� ��d������P�)�;� M�_�q��*�<��i� ��������)���M� _�q������������ ����<�û��=Oa s��>����* '9K]f� Q�������/ �%/7/I/�m//�/ �/�/�/n<��^/? %?7?I?[?m?/�?�? �? ?�?�?�?O!O3O �/<׹��?O�O�O�O �O�O�?�O_!_lOE_�W_i_{_�_�_FOXG9 +_�_�_oo(o:o�O Kopo�o)_�o�o�o�oP�o ��	g�0�o M_q���No� ���o�%�7�I�[� m�&l�n��Ə؏ ���� ��D�V�h� ��������ԟ柍� g�ڻ}�2�D�V�h�z� ��3���¯ԯ���
� �.�@�R���3uF�� ����¿Կ������ .�@ϋ�d�vψϚϬ� ��e�w���U�
��.� @�R�d�ψߚ߬��� ��������*���w� ��v������� w�����c�<�N�`� r�����=�w��-��� ��*<��`r ����������  ��1C Ugy�����<��    -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_��  
��(  }�%( 	 y_ �_�_�_�_�_�_o	o +o-o?ouoco�o�o�o:�Z* �Q &�J\n�� ����o���9� (�:�L�^�p������ ���܏� ��$�6� }�Z�l�~�ŏ����Ɵ ؟���C�U�2�D�V� ��z�������¯ԯ� ��
��c�@�R�d�v� ����᯾�п�)�� �*�<�N�`ϧ����� �Ϻ��������&� 8��\�n߀��Ϥ߶� ��������E�"�4�F� ��j�|������� �����e�B�T�f� x�������������+� ,>Pb��� ������� (o�^p��� ���� /G$/6/ H/�l/~/�/�/�/�/ /�/�/?U/2?D?V?�h?z?�?�/�`@  �2�?�?�?�3�7�P���!frh:\�tpgl\rob�ots\m20i�a\cr35ia.xml�?;OMO_O qO�O�O�O�O�O�O�O ���O_(_:_L_ ^_p_�_�_�_�_�_�_ �O�_o$o6oHoZolo ~o�o�o�o�o�o�_�o  2DVhz� �����o�
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ �ݟ��&�8�J�\� n���������ȯߟٯ ���"�4�F�X�j�|�@������Ŀ־�8.1� �?@88�?�ֻ�ֿ� 3�5�G�iϓ�}ϟ��� ���������5��A��k�U�wߡ߿��$T�PGL_OUTP�UT ;�!�!/ ������ ��,�>�P�b�t�� ������������ (�:�L�^�p�������������2345678901������ ���"��BT fx��4�����
}$L^ p��,>���  //$/�2/Z/l/~/ �/�/:/�/�/�/�/?  ?�/�/V?h?z?�?�? �?H?�?�?�?
OO.O �?<OdOvO�O�O�ODO VO�O�O__*_<_�O J_r_�_�_�_�_R_�_ �_oo&o8o�_�_no �o�o�o�o�o`o�o�o "4F�oT|� ���\��}���@��0�B�T�e�@�������� ( 	 ��Џ����� �<�*�L�N�`����� ����ޟ̟���8� &�\�J���n�������@��ȯ���"������ �*�X�j�F�����|� ¿Կ��C���ϱ�3� E�#�i�{�忇ϱ�S� ���������/ߙ�S� e�߉ߛ�y߿���;� ������=�O�-�s� ���ߩ��]������� �'����]�o���� ��������E����� 5G%W}����� �g���1� Ug	w�{�� =O	//�?/Q/// u/�/��/�/_/�/�/ �/�/)?;?�/_?q?? �?�?�?�?�?G?�?O �?OIO[O9OO�O�? �O�OiO�O�O�O!_3_ �O_i_{__�_�_�_��_�_�R�$TPOFF_LIM >�|op:��mq�bN_SV`  �l�jP_MOoN <6�d�opop2l�aST�RTCHK =�6�f� bVTCOMPAT-h�af�VWVAR >rMm�h1d �o� �oop`ba_�DEFPROG �%|j%ROB�195_SERV�	�j_DISPL�AY`|n"rINST_MSK  t|w ^zINUGp��odtLCK�|}{QUICKMEN��dtSCRE�p�6��btpsc@dt�q��b*�_.��ST�jiRACE_CFG ?Mi��d`	�d
?��u�HNL 2@"|i����k r͏ ߏ���'�9�K�]��w�ITEM 2A��� �%$12�34567890<����  =<��П<��  !���p��=��c��^� ���������.���R� �v�"�H�ί��Я� �����*�ֿ���r� 2ϖ�����4�޿�ϰ� ��&���J�\�n���@� ��d�v��ς������ 4���X��*��@�� ���ߨ������� T���x������l� �������,�>�P��� ����FX��d���� ��:�p" ��o����� F6HZt~�� N/t/�/��// /2/ �/V/?(?:?�/F?�/ �/�/j?�??�?�?R? �?v?�?QO�?lO�?�O �OO�O*O|O_`O _ �O0_V_h_�Ot_�O_ _�_8_�_
oo�_@o �_�_�_Lodo�_�o�o 4o�oXojo3�oN�o r��o��s��S�B���z� 3 h��z ��C�:y
 P�v�]���~�UD1:\������qR_GRP� 1C��� 	 @Cp���@$��H�6�l�Z��|� ����f���˟���ڕ?�  
���<� *�`�N���r������� ޯ̯��&��J�8�Z���	�u�����s�SCB 2D� �����(�:��L�^�pς��|V_C�ONFIG E��� ��~����Ϝ�OUTPUT� F���� ��5�G�Y�k�}ߏߡ� �������������#� 6�H�Z�l�~���� ����������%�9� K�]�o����������� ������"�5GY k}������ �1CUgy �������	/ ,?/Q/c/u/�/�/ �/�/�/�/�/??(/ ;?M?_?q?�?�?�?�? �?�?�?OO$?7OIO [OmOO�O�O�O�O�O �O�O_ O2OE_W_i_ {_�_�_�_�_�_�_�_ oo._AoSoeowo�o �o�o�o�o�o�o ������!�6oew� �������� +�=�0oa�s������� ��͏ߏ���'�9� J�]�o���������ɟ ۟����#�5�F�X� k�}�������ůׯ� ����1�C�T�g�y� ��������ӿ���	� �-�?�P�c�uχϙ� �Ͻ���������)� ;�L�^�q߃ߕߧ߹� ��������%�7�I� Z�m��������� �����!�3�E�V�i� {��������������� /AR�d�w� �������+=O2u���k}gV�Kv� ���////A/S/ e/w/�/�/�/`�/�/ �/�/??1?C?U?g? y?�?�?�?`�?�?�? 	OO-O?OQOcOuO�O �O�O�?�O�O�O__ )_;_M___q_�_�_�_ �O�O�_�_oo%o7o Io[omoo�o�o�o�_ �o�o�o!3EW i{����o�� ���/�A�S�e�w� ������������ �+�=�O�a�s����� ����̏ߟ���'� 9�K�]�o��������� ȟۯ����#�5�G��Y�k�}�������ž��$TX_SCRE�EN 1G�g�}i�pnl/��gen.htmſ�*�<��N�`ϽPan�el setupd�}�dϥϷ����������ω�6�H�Z� l�~ߐ�ߴ�+����� ��� �2�߻�h�z� ������9�g�]�
� �.�@�R�d������ ����������}��� <N`r��; 1��&8� \��������QȾUALRM_�MSG ?��� �Ȫ-/?/p/ c/�/�/�/�/�/�/�/�??6?)?Z?%SEoV  -�6�"ECFG Iv��  ȥ�@�  A�1  w B�Ȥ
 [? ϣ��?OO%O7OIO�[OmOO�O�O�G�1G�RP 2J�; 0Ȧ	 �?�O �I_BBL_NO�TE K�:T?��lϢ��ѡ�0RDEFP�RO %+ (%N?u_Ѡc_�_�_�_ �_�_�_o�_o>o)o�boMo�o\INUSER  R]�O�o�I_MENHIS�T 1L�9  �( _P��'�/SOFTPAR�T/GENLIN�K?curren�t=menupage,69,1�opBTfx �(
~253/������p)�~381,23�L�^�p��	#�71�̏ޏ�����q0��uedi�t(rROB195t0RV��Y�k�}����(�7H�ԟ���
����)q10X�j� |�����/���4H�ܯ � ��5R�`q|oB� T�f�x������1�ƿ ؿ���� ϯ�D�V� h�zόϞ�-������� ��
�߫Ͻ�R�d�v� �ߚ߬�;�������� �*��N�`�r��� ��7�I�������&� 8�#�\�n��������� ��������"4F ��j|����S ��0BT� x�����a� //,/>/P/�t/�/ �/�/�/�/�/o/?? (?:?L?^?I��?�?�? �?�?�?�?�/O$O6O HOZOlO�?�O�O�O�O �O�OyO_ _2_D_V_ h_z_	_�_�_�_�_�_ �_�_o.o@oRodovo o�o�o�o�o�o�o �o*<N`r�o? ������ 8�J�\�n�����!��� ȏڏ��������F� X�j�|�����/�ğ֟ �������B�T�f� x�����+�=�ү��� ��,���P�b�t���������z�$UI_�PANEDATA 1N���ڱ�  	��}/frh/�cgtp/wid�edev.stm� ?_fonts?ize=14��!��3�E�W� )pr�imYς�  } } �itree�� �Ͼ�������[��)� �M�4�q߃�jߧߎ� ���������%�7���[�7��� �   V{v��flex���6e���������J�ual��"��ϧ�X� j�|�����G������� ����BT;x _������i� ݰܳ7�-?Q cu����0�� ��/!/3/�E/i/ P/�/t/�/�/�/�/�/ ???A?(?e?w?^? �? �?�?�?OO +O~?OOaO��O�O�O �O�O�OFO_�O'_9_  _]_D_�_�_z_�_�_ �_�_�_o�_5o�?�? Eo}o�o�o�o�o�o*o �onO1CUgy �o������� 	�-��Q�8�u���n� ����Ϗ�Tofo�)� ;�M�_�q�ď���� ˟ݟ���z�%�I� 0�m�T�������ǯ�� ����!��E�W�>� {�� ���ÿտ��� �^�/�Aϴ�e�wω� �ϭϿ�&�������  �=�$�a�s�Zߗ�~� �ߢ��������� %�]�o�����
� ��N����#�5�G�Y� ��}���v��������� ����1UgN@�r��4�F���@�"4FX)� }��l����� /j'//K/2/D/�/ h/�/�/�/�/�/�/�/�#?5??Y?��C�=���$UI_POST�YPE  C��� 	 �e?�?�2QUICK�MEN  �;��?�?�0RESTO�RE 1OC��  ��*defaul�t�;  REE�VIEW:LDU�AL�?mmen�upage,107,1fO�O�O�O�O�rDozF381,26,22�O_ _2_D_ mF_j_|_�_ �_�_EAL?�_�_G_�_ "o4oFoXojoo�o�o �o�o�oyo�o0 B�_Oas�o�� �����,�>�P� b�t��������Ώ�� �������L�^�p� ����7���ʟܟ� � ��$�6�H�Z�l��!� ����������� � 2�կV�h�z�����A��¿Կ���
��=SC�K@N ?�=�u1sc+@uU2K�3K�4K�5Kĕ6K�7K�8K��2U�SER-�2�D�ksTMì�3��4��5�ĕ6��7��8���0N�DO_CFG �P�;� ��0PDA�TE ����None�2��_INFO 1QC�@��10%�[��� Iߊ�m߮��ߣ����� �����>�P�3�t���i���<-�OFFS_ET T�=�� ��$@������1�^� U�g������������ ����$-ZQcu���?�
�����UFRAME  �����*�RTO?L_ABRT	(��!ENB*GR�P 1UI�1Cz  A��~��@~���������0UJ�9MSK  M@�;-N%8�%��/��2VCCM��V��ͣ#RG�#Y�9����/����D�BeH�p71C����3711?�C0�$MRf2_�*S��괰	���~XC56 *�?�6�Y��1$�5����A@3C��. 	��8�?��OO KOx1FOsO�5�51ⴰ_O�O�� B����A2�DWO �O7O_�O8_#_\_G_ �_k_}_�__�_�_�_��_"o�OFoXo�%TCC�#`mI1�i���u��� GFS�»2aZ; �| 2�345678901�o�b�����o@��!5a�4BwB�`�56 311:�o=L�Br5v1�1~1�2 ��}/��o�a��# �GYk}�p�� �����ُ�1�C� U�6�H���5�~���ߏ����	���4�dSEGLEC)M!v1b3��VIRTSYN�C�� ���%�SIONTMOU�������F��#b������(�u FR:\�H�\�A\�� ��� MC��L�OG��   U�D1��EX����'� B@ �����̡m��̡  �OBCL�1�H�� �  =	 �1- n6 � -������[�,xS�A�`=��͗���ˢ��TRA�IN⯞b�a1l�
�0d�$j�T2cZ; (aE2ϖ�i�� ;�)�_�M�g�qσϕ� ���������	��F�STAT dmB~2@�zߌ�*j$i�\���_GE�#eZ;7�`0�
� 0}2��HOMIN� �f������ ~�����БC�g��X���JMPERR� 2gZ;
   ��*jl�V�7������ ��������
��2�@��q�d�v�B�_ߠREr� hWޠ$LEX�ԹiZ;�a1-e��V�MPHASE  �5��c�!OF�F/�F�P2n�jJ�0�㜳E1�@��0ϒE1!1?s#33�����ak/�@kxk䜣!W�m[�䦲�[����o3;� [ i{���� /�O�?/M/_/q/ ��/��//�/'/9/ �/=?7?I?s?�/�?�/ �/�?�??Om?O%O 3OEO�?�?�O�?�O�O �?�O�O�O__gO\_ �OE_�O�_�O�O/_�_ �_�_oQ_Fou_�_|o �o�_�oo�o�o�o�o ;oMo?qof-�oI �����7� [P��������� ˏ��!�3�(�:�i��[�ŏg�}������TD_FILTEW��n�� �ֲ:���@���+�=�O�a� s���������֯� ����0�B�T�f�x����SHIFTME�NU 1o[�<��%��ֿ����ڿ� ���I� �2��V�h� ���Ϟϰ�������3��
�	LIVE/�SNAP'�vs�fliv��E�����ION * U<b�h�menu~߃������ߣ���p����	����E�.ォ50�s�P�@� �Z�AɠB8z�z�!�}��x�~�P���  ���MERb���<�0���kMO��q���z��WAITDINE�ND������O9K1�OUT���SD��TIM����o�G���#����C���b������RELEASE������TM�������_�ACT[�����_DATA r�%L����xRD�ISb�E�$X�VR�s���$Z�ABC_GRP �1t�Q�,#�r0�2���ZIP�u'�&����[�MPCF_G 1	v�Q�0�/� �w�ɤ� 	|�Z/  85�`�/�/H/�/l$?��+ �/�/�/?�/�/???|r?�?  �D0 �?�?�?�?�?�;����x�]hYLI�ND֑y� ���� ,(  * VOgM.�SO�OwO�O�M i?�O�O^PO1_ �OU_<_N_�_�O�_�_ �__�_�_x_-ooQo�8o�_�o�oY&#2z� ���oC� e?a?>N|�oq��햋qA�$DSPH�ERE 2{6M� �_�;o���!�io |W�i��_��,��Ï ���Ώ@��/�v��� e�؏��p�����������ZZ�� � N