��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA �� �FT�{ @� LOG_8	�CMO>$D?NLD_FI:��SUBDIRCA�P�v� �8 .� 4� H�AD_DRTYP�H �NGTH����z +LS�&�$ROBOT2P�EER2� MAS�K4MRU~OM�GDEV�� R�CM+ �;$Z ��QSI�Z�X�� TAT�USWMAILS�ERV $PL�AN� <$LI}N<$CLU����<$TO�P$�CC�&FR�&�J�EC�!�%ENB{ � ALARl!�B�TP�3�V�8 S��$VAR9M ON
6��
6oAPPL
6PA� 85B 	7POR��#�_�!�"ALERT��&�2URL }}�3ATTAC���0ERR_THRO�3US�9z!�800�CH- Y�4MAXvNS_�1�A�MOD�AI� �$B� (APW7D  � LA �0v�NDATRYQFDELA_C@y'>A�ERSI�A�'R]OtICLK�HMR0��'� XML+ :3S/GFRM�3T� X�OU�3PING_�_COPA1�Fe3�A�'C�25�B_AU��� k 6R,2COU|�!H!UMMY1RW�2?�RDM*�� $DIS�.� SMB�	"�BCJ@"CI2�AIP6EXPS��!�PAR��TC�L�
 <(C<�0�SPTM�E� GPWR��X�V�Ro l5��!��"%�7�ICC�%H� kfR�0leP� O_DLV��YNo�3 <oNbX_��P~#Z_INDE�
C�`OFF� ~U�R�iD��c�  ? t �!�`'MON�%sD�&rHOU�#EWA,vSqx;vSqJvLOCA� �Y$N�0H_H-E���@I"/ }3 $ARPz&4�1F�W_\ �2I!F�`;FA�Dk0�1#�HO_� IN�FO�sEL	% �P K  !k0W�O` $ACCE� LVZk�2�H#ICE�L��  �$�s# �S��k���
��
`�rK`SQi�]���5|�I�0AL`h�z�'0 ��
����F����]��܅��$� 2ċ ��w������� č��!r�Z���4����Ċ!147�.87.224.�20h�S���96�����܁܁3�_{p_�  ċ� ?bfh.ch̟� 1�C�U�g�y����������ӯ^�� _FLT�R  ��π *��������n�ndxč2n��rSH�P�D 1ĉ � P!
robs?tation֯՚!k�.�Q�ſ ��������޿?�� c�&χ�JϫϽπ��� �����)���M��"� ��Fߧ�j��ߎ��߲� ��%���I��m�0�� T��x�������� 3���W��{���P��� t������������� Sw:�^�� ����= ah$Zׯ$ _L�A�1��x!1.��ğP�1�Q�255.%�S	���2��E �//*/<&3F/��  l/~/�/�/<&4�/�@50�/�/??<&56?���0\?n?�?�?<&6 �?�%@�?�?�?
O1��?P��MY� MY��c���� Q� �VN<�O�O_�O+_@=_O_"_s_�_NPd_ �_�_�_�_�_o!o3o �_Woio{oVNLoM ��o�l�oAo
.�@U}iRCo�nnect: i�rc\t//alertsE���� Pu����1�C��UуP_R8�d��H�~�������Ə؏ ���� �2�D�V�S$���8�(p����o ͟ߟ��QA8�	�d�A�B4��j�h�9�Q+��@DM_�A+��SMB 	X�8%ğVO���߯���_CLNTw 2
X� 4C�ɯ0��l�c�B�T� ��x���Ͽ������ )�;��_�q�Pϕ���MTP_CTRL ��%���ϙd c���ߋ��?�*�c�d�l��N���@{��Vߵ�Ƥ��������ѓC��USTOOM {���}�@ }�DTCP+IPu�{��h�E.�TEL�{��A=���H!Ta�t��çroblo�lr�  ���!KCL���F�>�!CRT����������!CO#NS&����n+���