��   u��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����UI_CON�FIG_T  �� A$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�62�ODE�
3�CFOCA �4VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�;�  &USTOM~0 t $} RT_SPID�r,DC4D*PAG� �?^DEVIC�EPISCREuE�F��IGN�@$/FLAG�@C��1  h 	$P�WD_ACCES� E �8��C��!�%)$LABE�� $Tz jа@�3�B�	CUS�RVI 1  < `�B*�B��A7PRI�m� t1�RPTRIP�"m��$$CLA�@ O���sQ��R��RhP\ SI�qW�  �5�QIRTs1q_�P'�2 L3hL3!�pR	� ,��$?����R�P�S�S��Q�� , ��  o��
� ��)/SOF{TP.@/GEN�1�?current�=menupag�e,1133,1�8o�o�o�o��Mo_o,1388vo/NA �'�o�n9�o������ocmc4�80|�%�7�I� �zQa�s��������� ͏\����'�9�K� ڏo���������ɟX� ����#�5�G�Y�� }�������ůׯf������1�C�U��� TPTX���y�򨑿o� s ��o���$/so�ftpart/g�enlink?h�elp=/md/;tpia.dgd�����"�4��r&ɿۻpwd꿁ϓϥϷ�� �������#�5���Y� k�}ߏߡ߳�B�T��������1�C�����zQ'f	oC ($ �ߕ���������i  zQ�Q�c�SHj�n������
)���Q(a��*������  ��P����@��n���8��P#`  �V������SB 1�XR_ \ }�%`REG V�ED�� wh�olemod.h�tm4	singl�Edoub\�triptbrows�@�! ����/A�S|�/Adev.sJl�o�1�	t���w �G/Y/k/5/�/�/�/8�/�/ ?� �P? *?<?N?`?r?�?�?�? �?�6�@?�?�?�? O 2ODOE	�/�/wO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_��_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?? z������� 
��O@�R�!�3��� ��QOcOI�ݏ�� *�%�7�I�r�m���� ����ǟٟ�����_ /�)�W�i�{������� ïկ�����/�A� S�e�w�����iֿ� ����0�B�T�f�x� s��Ϯ�}Ϗ����ϭ� ����>�9�K�]߆߁� �ߥ����������� #�5�^�Y�k�9���� ������������1� C�U�g�y��������� ������ſ2DVh z�������� 
��@R	�� �������/ */%/7/I/r/m//�/ �/�/�/���/�/?!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SO!�O�O�O�O�O�O �O__0_+T_f_5_�G_�_�_�Z�$UI�_TOPMENU� 1�P�QR 
d�Q�fA)*defa�ultqOZM*�level0 *\K	 o� So��_Qocbtpio�[23]�(tpst[1�heo�ouo�3oEo�-
h58e?01.gif�(?	menu5&yp�Hq13&zGr%zEt4M{4�a����� ����eB�C�U��g�y�����,�pr�im=Hqpage,1422,1�� ݏ���%�0�I�[��m������2���c?lass,5��០���)�4���130�f�x�������5���53ʏ����( �2�5���8ٯm� �������4�ٿ����!�3�^I�P�Q�_ k�m]��a[ϕ�ϝf�ty�m�o�amf[�0�o��	��c[1364�g.�59�h�a���k�Ax2uK}�� azmWw%{�ߩsK�]� 6�H�Z�l�~�ɿ��� ��������� �2�D� V�h�z�	���2���� ������	��ʟ?Q cu�(T��� ����Ѥ1$�N�`r�����ainedic�����//�con�fig=sing�le&��wintpĀ /`/r/�/�/E��W��/{���gl[4@7��ow�?���!8��B� 6�i.?h?>82ڀ�??�?�?z\rLz\r4s&x�? OVx `�6O��O�O�O�O�O �O��O_#_5_G_Y_ k_�O�_�_�_�_�_�_z,$;4$doub?%�o��13ؠ&du�ali38#�,4�_Pobo�_9o,n'o 9ato�o�o�o}_, >Pbt��� ��������o4�F� X�j�|������ď֏���=J�/,�wω� ����YOw���s�͔����ϡ�u��l�V�ȟ�.��?RO<��߬ߚ�6��u7��� ���� �/�A���e�w����� ����N������+�(=�O�."$13�� �ϭϿ���ܿ���� +�=�O���s߅ߗߩ� ������"���'�9�K�]�����6d���`������,$۬74�@�/�A�S�e�C�����?�	TPTX[G209�,���2�(��������1I8��(
����0P2���10_�1�Y�tv���H���0�
�1�
�ïqC:4$treeOviewA#.f3�~�m381,26=o ���l����/ /+/�O/a/s/�/�/�/�_B�5$oq� ?)?;?F/_?q?�?�? �?�?H?�?�?OO%O�7O�/�/�1�/r2pV��O�O�O �6XO�edit2azO�O _._@_�?���OS L_�_�_�_~��_�_G� o}o�CoUogoyo �o�o�o�o/o�o�o	 -?Qduӥ� �������?2� D�V�h�z������ ԏ���
����@�R� d�v�����)���П� ������<�N�`�r� ����%���̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� �_�_X�o|��o��� �����������ߋ� )�S�e�x߉ߛ߭߿� �ߓ��,�>�P�b� t￿���������� ���(�:�L�^�p��� ������������ �� $6HZl~� ������ 2 DVhz��� ���
/�./@/R/ d/v/�/7�IϾ/m��/ I���??)?;?M?`? q?�?�/�?�?�?�?�? OO%O7O��nO�O�O �O�O�O�O%/�O_"_ 4_F_X_�O|_�_�_�_ �_�_e_�_oo0oBo Tofo�_�o�o�o�o�o �oso,>Pb �o������� ��(�:�L�^�p�� ������ʏ܏/�/ $��/H��?MOk�}��� ����ş؟�W���� 1�C�U�h�y�����_O ԯ���
��.�y�@� d�v���������M�� ����*�<�˿`�r� �ϖϨϺ�I������ �&�8�J���n߀ߒ� �߶���W������"� 4�F���X�|���� ����e�����0�B��T���*def�aulta�2�*?level8��������{� t?pst[1]���ytpio[#23��u�������	menu_7.gif�
�13�	�5�
��
�4�u6�
ʯ? Qcu����� ��//�;/M/_/�q/�/�/�/6"pr�im=�page,74,1�/�/�/�??+?6"�&cl?ass,130?f?@x?�?�?�?=?O25�?@�?�?O O2O5#D< �?lO~O�O�O�O�/�"18�/�O__'_9_DON26@_u_�_�_�_��_��$UI_U�SERVIEW �1��R 
���_>��_
o�m(oQoco uo�o�o<o�o�o�o�o �o);M_qo ~������ %��I�[�m������ F�Ǐُ������ .�@���{�������ß f������/�ҟS��e�w�����F�*z�oom��ZOOM��W�I��$�6�H� Z���~�������ƿi������ �2�DϦ�m�axresH�MAXRES߯E�� �Ͼ������ϗ��*� <�N�`�߄ߖߨߺ� ��w�������o�%�J� \�n���5������ �����"�4�F�X�j� �w������������ ��BTfx� �?������ '=�t��� �_��//(/� L/^/p/�/�/?�/�/ �/7/�/?$?6?H?Z? �/~?�?�?�?�?i?�? �?O O2O�/?OUOcO �?�O�O�O�O�O�O
_ _._@_R_d__�_�_ �_�_�_sQ