��  I��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT  &2�*� � ��  �$$CLA�SS  ���������� V�ERSION��� �5�IRTUAL��' � 1 � T����CR-�35iA���  �aiS12/4000 80H�
H1 DSP�1-S1��	P�01.00W, � 	� ��
]�  ��# �:�������� {�F�2�r9  ��9����� HH� � ����� ���Ϋ C ��Z �
t
t������ ��s� 1�2��?��u�|��u3�	8�����&��<
=� ^ ����� J���hI�����; 2 �� ����H�a����~#��	�  �� !� �� �:?8����'by��c/�/�/�/?���?;?;(X?j?|?��1��3C(  �b����I�I2.���>�����wm"�܎?�?"4��<N`6i2�|2��� �����׶���{����4	����� @l�� 
����n�m �'!�!%F���� 34���=��!�	����;�	':+�J V W
��R UV$jO�������z's��-   ���(�%c	�	`�� �#
��%z�'� �
B _�_�_�_�_$?�_��3�_o+o=o��4����<���.���L.��m5�����;7�����; 	EFođo���c�?S%b8gw3|b�@ORK �&��m��ptG�p����S�8gHB\P�@��.��+ I'7�A7�a#����2�B+�0�����+;= ��x":+�� ����� �X"�|�o�� ��Z2Xw�����)�(w)B�"� d�#�c A��#=:rY:q�K� ]�o����_�� oɏۏ ����#�5�G��&�Bt�oR�b4/5!A4�k4|4�ov�����ϓH�X��!2�D��K�99~��5
� �������l�� ���w�0��%'���S@A�S�u� ����� 5V$��b�(S ��z#�V@��� �cXR7 (��t Zֲ#=rY�!���@�'�9���]���fd� ��������ѿ�����6d�Nb�iSR1C��x5�|}���˚p��`�M�����tG���������"�� D@�r��X��$�  �b*�<���#  z�  V$�rA�? ���Y���P�B�����`��(�%��ZP2Σ� Au��$�rZT�C� ��������L��p�9� K�]�o��������;" �R@�r6�|�h�zό̜`R=�V����Ϻ����� ����Ͻ���>U`� ��x�V$y����C|�Cz#�� ��O���;�(|ߎߠ�i {���������/ASew�����xPTa��Ng�	�,����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?P<�P?t?�?�?�?�?�? �?�?OO(O0C�� FO����O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o ^?&o8oJo\ono�o�o �o�o�o�o6OhOZO# ~O�OXj|��� ������0�B� T�f�x�������
o�� �����,�>�P�b� t������o����*< N�(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�ȏ���� ��ƿؿ���� �2� D�V�ҟğn����� ������
��.�@�R� d�v߈ߚ߬߾����� ����*N�`�r� ������������ ^ϐς�K��ϸπ��� ������������" 4FXj|��� ��2��0B Tfx����� ��R�d�v�>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?��?�?�?�? OO $O6OHOZOlO~O�� �O/"/4/�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo �?vo�o�o�o�o�o�o �o*�O�O�Os �O�O������ �&�8�J�\�n����� ����ȏڏ���Zo� 4�F�X�j�|������� ğ֟�D� �z� �f�x���������ү �����,�>�P�b� t������������ ��(�:�L�^�pς� �Ϧ�"����8�J�\� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z�ֿ����� ������
��.�@�R� �����ϛ�������� ��*<N`r ������� &��8\n�� ������/l� 5/(/�������/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?@OO,O>OPObO tO�O�O�O�O�OJ/</ �O`/r/�/L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �?�o�o�o�o 2 DVhz�O_�O� _0_�
��.�@�R� d�v���������Џ� ���*�<�N��o`� ��������̟ޟ�� �&�8��]�P��� ���ȯگ����"� 4�F�X�j�|������� Ŀֿ����h�0�B� T�f�xϊϜϮ����� ����r�d�߈����� t߆ߘߪ߼������� ��(�:�L�^�p�� ������&��� �� $�6�H�Z�l�~����� ��0�"���F�X� 2 DVhz���� ���
.@R dv������ �//*/</N/`/�� �/x/���/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4O�XOjO|O�O�O�O �O�O�O�O__�/�/ 6_�/�/�/�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o NO(:L^p� ����&_X_J_� n_�_H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������o�� ԟ���
��.�@�R� d�v���������,� >���*�<�N�`�r� ��������̿޿�� �&�8�J�\ϸ��ϒ� �϶����������"� 4�F�¯��^�د��� ����������0�B� T�f�x�������� ������v�>�P�b� t��������������� N߀�r�;�ߨ�p� ������  $6HZl~�� ��"���/ /2/ D/V/h/z/�/�/�/ �/�/BTf.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O��O�O�O�O�O_ _&_8_J_\_n_�/�/ �_ ??$?�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B �Ofx����� ����v_�_�_c� �_�_������Ώ��� ��(�:�L�^�p��� ������ʟܟ�J � $�6�H�Z�l�~����� ��Ưد4����j�|� ��V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬ������ ����*�<�N�`�r� �ߖ�����(�:�L� �&�8�J�\�n��� ������������"� 4�F�X�j��ώ����� ��������0B �����ߋ������ ��,>Pb t������� //r�(/L/^/p/�/ �/�/�/�/�/�/ ?\ %??���~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O0/�O
__._@_R_ d_v_�_�_�_�_:?,? �_P?b?t?<oNo`oro �o�o�o�o�o�o�o &8J\n�� �O������"� 4�F�X�j��_�_�_�� o o�����0�B� T�f�x���������ҟ �����,�>��P� t���������ί�� ��(���M�@���̏ ޏ����ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������X� �2� D�V�h�zߌߞ߰��� ����b�T���x����� d�v��������� ����*�<�N�`�r� ������������� &8J\n�� �� ���6�H�" 4FXj|��� ����//0/B/ T/f/��x/�/�/�/�/ �/�/??,?>?P?� u?h?���?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O __ $_�/H_Z_l_~_�_�_ �_�_�_�_�_o�?|? &o�?�?�?�o�o�o�o �o�o�o
.@R dv������ >_��*�<�N�`�r� ��������oHo:o� ^opo8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������ į֯�����0�B� T�f�x�ԏ����
�� .�����,�>�P�b� tφϘϪϼ������� ��(�:�Lߨ�p߂� �ߦ߸������� �� $�6ﲿ��N�ȿڿ� ����������� �2� D�V�h�z��������� ������
f�.@R dv������ >�p�b�+���`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/?"? 4?F?X?j?|?�?�?� �?�?2DVO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�/�_�_�_�_�_�_ oo(o:oLo^o�?�? vo�?OO�o�o  $6HZl~�� ������ �2� �_V�h�z������� ԏ���
�fo�o�oS� �o�o��������П� ����*�<�N�`�r� ��������̯ޯ:�� �&�8�J�\�n����� ����ȿ$���Z�l� ~�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ������� ������,�>�P�b� t��������*�<� ��(�:�L�^�p��� ������������  $6HZ��~�� ����� 2 �����{����� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/?b?<?N?`?r? �?�?�?�?�?�?�?L OO���nO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_ ?�_�_oo0oBo Tofoxo�o�o�o*OO �o@OROdO,>Pb t������� ��(�:�L�^�p��� �_����ʏ܏� �� $�6�H�Z��o�o�o�� �o؟���� �2� D�V�h�z�������¯ ԯ���
��.���@� d�v���������п� ����t�=�0Ϫ��� Ο�ϨϺ�������� �&�8�J�\�n߀ߒ� �߶�������H��"� 4�F�X�j�|���� ����R�D���h�zό� T�f�x����������� ����,>Pb t������� (:L^p� �����&�8� // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?�h?�?�?�?�? �?�?�?
OO.O@O� eOXO����O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o op?8oJo\ono�o�o �o�o�o�o�o�ozOlO �O�O�O|��� ������0�B� T�f�x���������ҏ .o����,�>�P�b� t�������8*� N`(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~�ڏ�� ��ƿؿ���� �2� D�V�h�ğ�π���� �����
��.�@�R� d�v߈ߚ߬߾����� ����*�<`�r� ������������ �&��ϔ�>������� ������������" 4FXj|��� ����V�0B Tfx����� .�`�R�/v���P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�? OO $O6OHOZOlO~O�O� �O�O"/4/F/_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo do�?�o�o�o�o�o�o �o*<N�O�O f�O�O_���� �&�8�J�\�n����� ����ȏڏ����"� ~oF�X�j�|������� ğ֟���V�zC� ��x���������ү �����,�>�P�b� t���������ο*�� ��(�:�L�^�pς� �Ϧϸ������J�\� n�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z��述��� ������
��.�@�R� d�v����ώ���,� ��*<N`r ������� &8J��n�� ������/"/ ~�����k/�����/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?RO,O>OPObO tO�O�O�O�O�O�O</ _�Or/�/�/^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �oO�o�o�o 2 DVhz��__ �0_B_T_�.�@�R� d�v���������Џ� ���*�<�N�`�r� �o������̟ޟ�� �&�8�J������ � �ȯگ����"� 4�F�X�j�|������� Ŀֿ�����z�0� T�f�xϊϜϮ����� �����d�-� ߚ��� ���ߘߪ߼������� ��(�:�L�^�p�� ��������8� �� $�6�H�Z�l�~����� ����B�4���X�j�|� DVhz���� ���
.@R dv������ �//*/</N/`/r/ �� ���/(�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFO�XO|O�O�O�O �O�O�O�O__0_�/ U_H_�/�/�/�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o `O(:L^p� ������j_\_ ��_�_�_l�~����� ��Ə؏���� �2� D�V�h�z������� ���
��.�@�R� d�v������(��� >�P��*�<�N�`�r� ��������̿޿�� �&�8�J�\�n�ʟ�� �϶����������"� 4�F�Xߴ�}�p���� ���������0�B� T�f�x�������� ������,���P�b� t��������������� �߄�.�ߺ��� ������  $6HZl~�� ����F�/ /2/ D/V/h/z/�/�/�/�/ PB?fx@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O��O�O�O�O_ _&_8_J_\_n_�_�%��$SBR2 1� 5�P T0 �  C?7 �_�_�_o o2o DoVohozo�o�o�o�o�o�Q�o�_!3 EWi{���� ����o� A�S� e�w���������я� ����+��O�2�s� ��������͟ߟ�� �'�9�K�]�@���d� ����ɯۯ����#� 5�G�Y�k�}���r��� ��׿�����1�C� U�g�yϋϝϯ��Ϥ�~�_�����!�3�E� W�i�{ߍߟ߱����� �������(�:�L�^� p�����������  �����H�Z�l�~� ��������������  2D(�:�z�� �����
. @RdvZ��� ���//*/</N/ `/r/�/�/�/��/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�/�? O"O4OFOXOjO|O�O �O�O�O�O�O�O_�? 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o "_boto�o�o�o�o�o �o�o(:L^ pTo������  ��$�6�H�Z�l�~� �����Ə؏����  �2�D�V�h�z����� ��������
��.� @�R�d�v��������� Я���؟�*�<�N� `�r���������̿޿ ���&�
�4�\�n� �ϒϤ϶��������� �"�4�F�X�<�|ߎ� �߲����������� 0�B�T�f�x��n߮� ����������,�>� P�b�t����������� ����(:L^ p������� ��$6HZl~ �������/  /D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?6/v?�?�?�?�? �?�?�?OO*O<ONO `OrOV?h?�O�O�O�O �O__&_8_J_\_n_ �_�_�_�O�O�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�_�o 0BTfx��� ������o,�>� P�b�t���������Ώ �����(�:��^� p���������ʟܟ�  ��$�6�H�Z�l�P� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� �ϴ�����*�<�N� `�r߄ߖߨߺ����� �����&�8�J�\�n� ������������� �"���X�j�|��� ������������ 0BT8�J���� ����,> Pbt�j��� ��//(/:/L/^/ p/�/�/�/�/��/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�/O  O2ODOVOhOzO�O�O �O�O�O�O�O
__ O @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo 2_ro�o�o�o�o�o�o �o&8J\n �do������ �"�4�F�X�j�|��� �����֏����� 0�B�T�f�x������� ��ҟ��ȏ��,�>� P�b�t���������ί ������:�L�^� p���������ʿܿ�  ��$�6��D�l�~� �Ϣϴ����������  �2�D�V�h�Lόߞ� ����������
��.� @�R�d�v���~߾� ��������*�<�N� `�r������������� ��&8J\n �������� ��"4FXj|� ������// 0/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?F/�?�?�?�?�? �?�?OO(O:OLO^O pO�Of?x?�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�O�O�_�_o  o2oDoVohozo�o�o �o�o�o�o�_�o. @Rdv���� ������o<�N� `�r���������̏ޏ ����&�8�J�.�n� ��������ȟڟ��� �"�4�F�X�j�|�`� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ��Ŀ��(�:�L�^� p߂ߔߦ߸�������  ����6�H�Z�l�~� �������������  �2��(�h�z����� ����������
. @RdH�Z���� ���*<N `r��z��� �//&/8/J/\/n/ �/�/�/�/�/��/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?�/O 0OBOTOfOxO�O�O�O �O�O�O�O__,_O P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o B_�o�o�o�o�o�o�o  $6HZl~ �to������  �2�D�V�h�z����� ������
��.� @�R�d�v��������� П�Ə؏�*�<�N� `�r���������̯ޯ �����
�J�\�n� ��������ȿڿ��� �"�4�F�*�T�|ώ� �ϲ����������� 0�B�T�f�x�\Ϝ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ ������� ��2DVhz�� �����
//./ @/$d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?V/�?�?�?�?�? �?OO&O8OJO\OnO �O�Ov?�?�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�O�O�_oo 0oBoTofoxo�o�o�o �o�o�o�o�_,> Pbt����� ����(�L�^� p���������ʏ܏�  ��$�6�H�Z�l�