��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����DRYRUN�_T   � �$'ENB �4 NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��SAW_� G �%$INIT�	RESUME_/TYPEN &J�_  4 �$($FST_IcDX�P_ICI�0 �MIX_BG�-A
_NAM�c MODc_U�Sd�IFY_TqI�.yMKR-�  $LI�Nc   �_SIZcw� k�. , $USE_FL4 �p�&i*SIMA��Q#QB6'SC�AN�AXS+IN�S*I��_COUN�rRO��_!_TMR_VA�g�h>�i) �'�` ��R��!�+W[AR�$}H�!�{#NPCH���$$CLASS ? ���01���5��5%0VERS��.7  {�@2IRTU� �.?@0'/ l5+5�������Y0B�6m071�5��%71 �?���?
O��}5I2�;.FOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_��%F�W?N8�0 ����_�_�_��@��o { 2�;� 4%L_AN�D_Bt_���QI��%L Jo���:dLmu�%�[o�o7g�1zo�o 
�X�o�o�o�o���p
Oa@ �dvu�S���=�9@Y0ma`�s�1�t�a	l1Y0�>�&�8�J� \�n���������ȏڏ ����6�1��1 �2� D�V�h�z������� ԟ���
�44�6�S!�2�9  �[�m��������ǯ ٯ����!�3� �M� f�x���������ҿ� ����,�>�I�b�t� �ϘϪϼ�������� �(�:�L�W�p߂ߔ� �߸������� ��$� 6�H�S�e�~���� ��������� �2�D� V�a�z����������� ����
.@Rd o�������� *<N`k} ������// &/8/J/\/n/F