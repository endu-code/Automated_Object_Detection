��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV����RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DISc �S�MB�	"�BC�J@"CI2AI<P6EXPS�!��PAR��SCL^�
 <(C�0��SPTM�E� P#WR��X�V�Ro l5��!�"Y%�7�ICC�%� �kfR�0leP� _GDLV��U�QNo�3 <oNbX_��P~#Z_INDE�
C�`OFF� ~U�R�iD��c�  ? t �!�`'MON�%sD�&rHOU�#EWA,vSqx;vSqJvLOCA� �Y$N�0H_H-E���@I"/ }3 $ARPz&4�1F�W_\ �2I!F�`;FA�Dk0�1#�HO_� IN�FO�sEL	% �P K  !k0W�O` $ACCE� LVZk�2�H#ICE�L��  �$�s# �S��k���
��
`�rK`SQi����5|�I�0AL`h�z�'0 ��
����F������܅��$� 2ċ T"�w������� č��!r�Z���4����Ċ!147�.87.224.�20h�S���96�����܁܁3�_{p_�  ċ� ?bfh.ch̟� 1�C�U�g�y����������ӯ^�� _FLT�R  ��π ,��]� ����n�ndxč2n��rSH�P�D 1ĉ � P!
robs?tation֯՚!k�.�Q�ſ ��������޿?�� c�&χ�JϫϽπ��� �����)���M��"� ��Fߧ�j��ߎ��߲� ��%���I��m�0�� T��x�������� 3���W��{���P��� t������������� Sw:�^�� ����= ah$Zׯ$ _L�A�1��x!1.��ğP�1�Q�255.%�S	���2��E �//*/<&3F/��  l/~/�/�/<&4�/�@50�/�/??<&56?���0\?n?�?�?<&6 �?�%@�?�?�?
O1��?P��MY� MY��c���� Q� �VN<�O�O_�O+_@=_O_"_s_�_NPd_ �_�_�_�_�_o!o3o �_Woio{oVNLoM ��o�l�oAo
.�@U}iRCo�nnect: i�rc\t//alertsE���� Pu����1�C��UуP_R8�d��H�~�������Ə؏ ���� �2�D�V�S$���8�(p����o ͟ߟ��QA8�	�d�A�B4��j�h�9�Q+��@DM_�A+��SMB 	X�8%ğVO���߯���_CLNTw 2
X� 4C�ɯ0��l�c�B�T� ��x���Ͽ������ )�;��_�q�Pϕ���MTP_CTRL ��%���ϙd c���ߋ��?�*�c�d�l��N���@{��Vߵ�Ƥ��������ѓC��USTOOM {���}�@ }�DTCP+IPu�{��h�E.�TEL�{��A=���H!Ta�t��çroblo�lr�  ���!KCL���F�>�!CRT����������!CO#NS&����n+���