��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS8?  �DMM�A@�  @ $��AbEREG_OFl�B�BME�HAS�C�1�A �DRE�-   � �0�B{F S{T� �M�DTRS$ST1D6XlQCWFA� 7X �QCW�"YV�"eS/ �A~7   $�@�TINd@�0SkUL� �R_@�  $}@ S�W@�RO�RR�%	 �P�T� Ɔ@JU� �SqFS;4D6
 �2P�0�_@cFOL[d!$FIL� jjEʄP�C�S�aDI~G4RC_SCA���cINTTH�RS_BIdA�dS�MAL�bCOL��bG�`� �� ��_IVTIM��$!0B"�$S?0xCCBDSDN��-qI2wT2w�DEBUdA\!SCHN�"TOfa0�!  � Q0mr<0V� ��;!�rAUTTUuN� TRQaʤuE40N �qFS'3AXG  � 1(eb}t�rI�v%�@�a|gr7 l �!|�3@WEIGH�qV�2 uS_5QF(�MT2�WA� 	pEs?NTERVA�; @- Q�� S!�t�AS0�S�$J-_ST�A�p JQg���1�(���2��3��W����� hqx��"COWG_X�Y�Z�6ҁCM�p?�p<�܂RSLT�4�@�D��D���r_�p9_�q7  �~�b#�0VROUNDCM?VPERIODA�w1PUU3F2D�'�TM1� �Ƒ_D<��GAMMc1^�TRXI�K�5K�K��CLbP�&�O00ADJ�GAVu�UPDB"�rI%0 ,$M"�P30f��� �d�:pG p"��HC�D�GV�#GVY:��Z�JDO5�,q���S��$R��E�_8@{٣�pA�PHBC��$#VF6�P��2L����@IL[����;� ��;�d@���RG����NEW_���r�Qp}���ڡ�5OBOA@�fY�sW2/�G<�	 ����ȴ\�2�E�KP��NUCNPRGO�V����@`d_TWԔc,�G�E^!NV02#C�c0@�WTS�TRL_SKI2!O$SJ�Q��NQp�GW��#��7 �\ ;0FR]b� � CMDC���T0�b���TO?�� � �5گ���_�Ah �0 '��ALARM��_�*�TOT6�F#RZn l�,!Y 3�� X!��mӥ�X �Œ`X P�ʕ�U#��2��2
�8X#Z���FIX�8�ґF�"��IT�`IeB�PN_d��CH��%��_DFL _�B#F2N�ڶ�3����� ��3�"�����ʷ�� ����3��3p
��X��DIA����/#� ���%�����[1��g1�[� ��Z��#��!���%���$0�@
p��7F���D�� HA�pU��5����v�FSIW.6 �2PN@�`uR>!�PHMP�`HCK%���>0G�'�*#e A����pN�T��^H	��HUFARzs3��A��Ugv�Ca�$v0Q �����@p@p ��  SI0�� P�5�I�RTU_��� %S�V 2���  � �6>0]@�]	Q�EF@� �oP�  @p P� �/@/'/9/K/U%@pd@p
m hK�/w/�/�/ �(��$��/� �/�/ ?.8e"�/?J?\?r? 8?�?|?�?�?�?�?�? �?>O4ObOO�OTO�O �OjO|O�O�O�O_�O (__\_f_�_B_�_�_ �_�_ o�_$o�_Ho>o o^b�/�ot��%�/�o��o�k	MC:� 5678  A�fsdt1 78901234qx#5w  	q 6xz.Ops�3'��j l�o�o����������,�5�DMM c�)5�A ���x�������=���O�R 2	Q� "��m��_� tu�B?)D�N�S4D 
FQ�!tY�d�!Ls`|�q`rƈ̀?�l��B𴐠�$ ON�FIG �}(�[ � ������i!�� 2��,
Hand guide���?�3��� � �X��с��ь��g#�=���A��ύ�������p �ݯ�(��L�7�p�x[����m*�� ����ʿܿ� ��$� 6�H�Z�lɌ��ό��� ���������
�C�E�]I 2Q�(�0� -�zՀ�F�M���_`πB��<��d�C�  ��uq�=#�
_aNnk=(��K����̥�@��e��=D�y���_a;�����8I��_aIt�$ �$F�>�s��k"���Q�Fۀ3]儢ѯǯ����!�/�``+��=���.�����_a�$敕��(4$������>�E���B<~w%�_a8�E�y5�;�j�A��Ҝ�Q�>��]�_a?��m���஑����~u1�?�3�3����0�:�o ����0�����LSB��~uq�ӻ���m�S]���/8��� ��� t�	eF|���P]��߯���x�n��;�.��z��3�'	���,��B���4*� 2/V��%D�DGH  *%v�+� �^-��
�/��/u/F~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?�;)�7�?�?�o�?�8J�hq�?�?zyjG�_F?SIW Q��9 ��O�O�Ou�