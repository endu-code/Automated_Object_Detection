��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk" 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&@B4��_sC3���r[R�_p�d`U��@VAD>CMVROU
b�1�PERIO�sF1P���2D-��3%T��1_D��2�Ĥ�3��T����K�9K��K�7CL���0�gADJ����_Udr�YRAUX�@�	 �4�@C�P?a�$� A�&�n@ qUX_AXS��PJF��� 
 h�D�rӠ�Cd��C�t �C�F�@�H�G1P�FOX�p4XAXISU� Tj��D͡�q�E�AP@M@ 	8BQ܀HR
$IDX\P�RV�QSa�GRT��L $F�E�_Uנ���TTOOL�R�p;�A��p�vy1DOf` \�>�0R_PKG�RQ{ BQ NR��PBQS�P[Q G2	hQ�P�S&�P2�Q�Qba�	�1ad��$VFLw0IM�,�LT�r�:a���Tc�6Tb����$�DYG��C$d0JgGUg	�d�4�d�cMPS>WP  �$ @��  ����aڐ@&�@ &�`VE�RSION�h�I@�5�aIRTUAL�o�avS�?�h&�  �aL|J\n� �������� "�4�F�X�j�|����� ��ď֏�����0��B�T�f�x��a+u|P1�1 29{\8�@I@�� ֓Ә~��  ?�a� @�@����A�  �����#���@�3��-�?�Q�?��g�U����  D�  Bp  =���Ϳ�?333?!�a�̠�̤@��ߥ�A ��/  & �G�P ?fffˡ>��ߥ��� ����0�ܙD���̤ˡ ��k�C�Z�[��`��0�����ӿٲ��B�ђǟI�ÿ��;���F@ K���������Dz��l�W�I��ٺ��ܑ�P`��!w���ēV��'�9� K�]�o�5ߓ���_�q� ۿ�������#�9� G�y�7�I�j�߳��� ��������a��!���y�3����ϋ�9� K�]�oρϓϙ���x� ��D���������� �,>�b���0���� ���`�ɤ����ȗ� Đؓ���2/d���@L����^/\�Ϣ�]��ĐW��"�@�"��'B����������/" � $đƚ�$1>B,4_��(����1?��x�?�?�8>����� ��//@/�?T/f/?O �/�/�/�/�/�/�O? ?,?>?P?b?;_�?__ �?�?�?�?�?OO(O �_o^OpO�O�O�O�O �O�O�O __$_�oH_ Z_3~_�W��fx���2�����	���o2�2-�V�h� z�������ԏ��� �����Dqdd�����l ��ߩߩ�b�����o��@��ğ���cd�p@(������qT�@� a>Ho�
}��[��c|�>LŠ���_v���O<#�
�Qsbp|���X��o�C���� a?e?a��3�T`��@  �G_�
�T���_@����x�2bo%{Bta �������1��U�g�k�`>X�ؤ�����^��It$ ��$$�K>�٢
���A���߭�'�����4�+�{��s�.����ރa$敕��(4�$ܛ�S�e�;��=.��>��H�Ճa�5����8M�	Y��;�=���3��a�B�	9�R�=�v�a� �ߡ����������m�����   �b\'������`k�S� K�X�,�w�������/�(����C��Q�??333;�s�<���saD/  C``G�P ?fff/a>$���?_	W�_�� 0��_g�;�5c?� 4'e��u<�j� F@ ��[�� DzI ����w5���y ܃�����/� ��/�/7I�_I/[/ m//�/�/�/�?�?�? �/?!?3?E?W?i?{?@�?kO}O�?�?�L�O q�O������ �O���O�O�_
__._ @_R_d_o�_�_,o�_ o�_�_oobo%``&/ $.(��? ��>�"��o����}� �o��E+̰�B��+� �ȴC��8�����{j 4�~gĠ{t��"�������$�3t7�q��<���>���3t� cu������� ���)�W���_�q� ����������ݏ�ȯ �%�7�I�k�%���� j���ǟٟ���Ϳ 3�E�W�i�{�a����� ��կ�L�o0��������2Q/�A�S�e�v�	Uώ�2�߲����� ������0�B�T�[ Ru���������7M ;	;	/�DO*GT�V�  �M�D�i���Op������Ѱ����A>��a��f��B�BH����>L! H���g�<'#�
�ϲp��w�p�E�v������A@��7������@\A �b�f��D?B,�� 7J���_���Bб�� �Z{�p��N���>�4_�U�/��It$ //$��>%�5
/a'A��a/�	/�/-/?&��+��=��%.����%���$敕�%(4$���%�/�+;��.�#5>��H/5��5���?58M�YK5��= g5��8�x?�+	�/�?�?�?�7? �?O$O6OHOZO�o�|GnlG  ;� �`�X���E�E�� �A��O�O�O	_�2 _�^����`=�e?333���B������D/  C��GÿP ?fff��> ���e�Y�Q�iȌO Vb�m����W�i�]o oo�o��k��_wo�o�`F@ uawU�`Dz�P$to��o�j"���� � �_�_oo'o�KoU �)��o�oﯥ�� ���1���"�Y� k�}�������ŏ׏� ǟٟX�1��̸k��o C��o'9KQ� ��0�B���f�x����� ����z�������l� >�P�b�t���lu�ς0\�nπϊx�O��� ����4�����C� <���R(����c� $�C� ���׺�� ڷ  �Ę�~Jk���_V�؏��/�?�Q�]�>�����]�� ��������+��O� a�s߅߳�U������� ������9�K�$o� ����������� �#�5�G�u�k�)�� ������������ 1ǼZό�/0/B/X%�2�l�/�/�/�/�-��"2�/? ?2?D? V?h?z?�?�?�?�d�n �>�GYGZ<���Y �Y�������ijO|O�O�O�FK �GLOP^Ib!W�#�> ��'_����4U>�L}PdQ�.B�<#�
K+p4_�B�8t�FB���� �SU�RkU@��lT ��o�δ���ζ��0o��eB,TUPo �o�o�o�o��P�>a�T�O�OrICI�t$ �$�&>��R
k�wAHD�e����v�@+��̞+�.���7��A$�敕G�(4$�xS���;��.��>��H���A5{����8M�Y���==dPÅ�B�ԏ�{	�
���.��g�Y� n���������%o�=��>ȗ  B� �R�T_b�P#��J� �X/�A�S�e��|�j��B�	��S��?3�33�E+��D7IcaD�/  CG�P_ ?fff�A>�Q 8D����O=X蟲� �M�O���o��˿ ���?Y�ӿ-�Kl�F@ _�k�ӥbl�Dz���k�]�/�p�~!^/P) �;� M�_�q���Iߧ���s� ����K��%�7� M�[ߍ�K�]�~���� �������!�3�u�#�5����Sl���)ϟ� M�_�qσϕϧϭ�GR ����X��������
 �@R�v�� �����/�ϸ����ȫ��  viڗ�N.k_=C��/ o�㢄`s���U�"�d �Q�f�PcEci3�/6 |P3$�ښ�$E>�Us��(��)o�<�?�8>�����:/-/ ?/Q/c/u/�/`O�/�/ �/�/?�O?)?;?M? _?q?J_�?�?�_�?�? �?O#O�_7OIO"omO O�O�O�O�O�o�O�O _!_3_oW_i_B�_�{���z���u2@	�����.�F�2A�j�|������� ď֏�����
�-� Xqxd�����l���� �b�����Ɵ؟���!�wd�p<�����(�qh�T�_a>\���}z�o� s��>L�٠�� o��y<#�	
�Q�bp��/�l��o.�c���_aSeWa��G�h`ǥ@�Ȥ[ s��T���_�V�ꌿFbo9{B�a����π3�E�(�i�{�.k�>�l�����ϥ�Itk$ ��$8�>��	
���A�����;�x����H�+��̇��.�����G�$�{����(4$ܯռg�y�;��.��>���H��G�5�=���8M�Y�O��=���G��a0�V�	 M�f�Q��u��ߵ��� ���� ����'��$�  �bp;� �����g�_�l�@� ��������C�����c���e��S?33�3O���P���ñD/�  Ct`G�P /?fffO�>8��� Ss	k�_!xD�s {�O�IwS�'H�;e#��/��j� F@ ��/o�� Dz] ����I8�q��y ܗ� ����//�/�/ K]�_]/o/�/�/�/ �/�/�?�?�??#?5? G?Y?k?}?�?�?O�OO�?g|�#O��O� ����/	_���O �O�__0_B_T_f_x_ 2o�_�_@o�_$o�_o o,ovo$%t:/&8B(�OPp\cҹ 6��o�~ǯ���o��E ?��BPp?��ܴW� ��L������jH��gؠ �tPq6�#������8��GtK߅���	��>���Gt�w�� ��������+� =�k��s��������� ͏����ܯ'�9�K� ]��9�����~�ɟ۟ ���-�#��G�Y�k� }���u���ů���l@D�������2e C�U�g�yߊ�iϢ�2����������� � 2�D�V�h�of��� Դ������KMO	O	C� XO>Gh�j"�4�a�X�}�ӴИ��������p�>�a��z�p�B�B\���>L5 �\���{�<#�
��p�����E,ϊ�����p������İ#@pA$�b� z�B�SB@�KJ���s���B�n�@������t >��Hs�i�*/�It$� C/$��>�I
#/u'A �u//�/A/�S&��+����%.�����%��$�=��%(4$�5�/��+;��.75>���HC5��5���S58M�Y_5��=@ {5��L��?�+	�/ �?�?�?�7?O&O8O�JO\OnO}K�$CC�SCH_GRP1�2 2�����A&� �\��Xo��  O��`�lt  �E�E���A�__,_�>_�2U_C^����`<Q�e?333��R�����#D/  C�аG�P ?fff��>���e�Y�Q �}��Ojb�m����W �i��o�o�o���2o�o�E`F@ `8uDa�U�E`Dz�P YtDo6�j6��� �o&o8oJo\o "��o�L�^��o�o� ����&�4�f�$� 6�W�������ď֏� ���N������f����x�&8J\ n�����e�w�1��� ����ѯ������+� ��O���s�������󿀡u�Ϸ�ϣϵϿxȄ���ٳ.��i�'� #��x�q�H��R<L� �����8�W� � ����4 ����J@���sLV�����/��t���>��� �Ē�����*�<�N� `�9��ߖߨߺ��ߊ� ����&�8�J�#n� ��Y��������� �"��F�X�j�|��� ��^��������� 0B/f�����S/e/w/�%2�l�/�/�/$�/=�22?C? U?g?y?�?�?�?�?�? �?�d�nN1!Q|Y|Z qȝ�Y�Y�՟�����i�O�O�O�O�FP�� W�O�I�!AW-3�>5�\_�S�H��iU>L�P�Q�cB��<#�
�`p�i_RE��V<B���,0�U bA�U@푡T4�Lo��В��fȚeo��B a�U�o�oBT�P>Ea�T�O�O��~CIt$ �$�6>��R
��wA�}D�����v!P+����`�.����l� Q$敕|�(�4$܈�@�R�;�{�.��>��H��� Q5��Ѕ8M�Y܅(M=�P�� R�	�/�	&�?�*�c� N���������ǟٟ��Zo Mؾ��  �I�b�T�b�PX� @�8JE�hd�v�����P�����<B�>��S,�?333(U`�)T|lI�aD/  CM�G�P ?fff(Q>amD,�L�D�� ���L�TM(_"�P� ,� �!��?���xbπ��F@ ��0���Hb��Dz6��Ā����d�"ʳ!�/�) �p���������~� ܿ�Ϩߺ�$�6π6� H�Z�l߂ߐ��߀�� ������� �2�D�V�h��X�j������� ��^����ϔϦϸ��� ����|R�������	 -?Qu� �����O���M/���/�� ��) 5�i���.�_ nC��/����`��)  e�"�d0a�f%`�E�i h!?k�Ph$)!��$ z>�U��8 $$�^ox�<�?�8>��� $ �:P/b/t/�/�/�/�/ �O�/�/??D?�OL? ^?p?�?�?�?_�?�? �_ OO$O6OXOolO ~OWo�O�O�O�O_�O �o _2_D_V_h_No�_ �_w�_l�/����u2>��.�@�R�c�B{�2v����� ÏՏ�����/�A� H�?�b��q�dةت�l $�(�(�r1��AC�@���:�1�V��d�p@q�ݟ��q����Ia>���S}���5sť>L���5o��TyO<#�
�Q�bpů�d���c������Ia�e�a�|��`��@ I������Sd,�o@۶$���{bLon{B�a ��G�h�z�]Ϟϰ�ckM�>��!�L�B��^ړIt$ �$m�K>�"�
��N�Aٔ�N���p��,�}�+�{�̼�.������|�$敕��(4�$��՜߮�;��=.�>��H�|��5��,�8M�	Y8儝=��T�|�%qe��	�ߛ���� �������#�5�G����\�4Y�   (r�p�E��M����� ����u���������x�(������*��?333����ș���D/  C�`G�P ?fff��>m�ɔ��	��_Vx y�C�����~��� J\}peX��d�<�j� F@ ��d��� Dz� $����~���y �����/8 B/??���_�/�/ �/�/�/�/?�?�?O F?X?j?|?�?�?�?�?@O�O�OEOO�L�XO �0_��//&/8/ >_آ_/_�_S_e_w_ �_�_�_go�_�_uoo Yo+o=oOoao�oY%�`o/I[mw(�<O �p�c�k�!�~��Γ 0)� Ut�R�pt� P�Č�0Ɓ������j }��g��t�qk�X�֎L�m�|t�ߺ�,�<>�J�>���|tJ� �������� <�N�`�r���B����� ̏ޏ���ۯ&�8�� \�n�������n�ȟڟ �����"�4�b�X�� |�������į����� ���p�Gy��/�E�2�xߊߜ߮߿�	����2������ 1�C�U�g�y��� �����	�4	4
)̀M �	�	xOsG�ϟW� i��������8����9�K�O����� Q>��a��R R��!�>Lj Q����<'#�
8��p!��p�EaϿ����� Q@��@���X@�A Y�b��w��Bu�7 �Jײ����B�A =�����/��� >�}����_/6�It$ x/$��>%�~
X/�'A5��/�R/�/v/�&��+��=�5.���$5���$敕45(4$��@5�/
;;��.�l5>��Hx5��5����58M�Y�5��=Q �5����?�+	�/�?�?OGT? FO[OmOO�O�O��|�n�G  �� p��L� U�E�� �A�_._@_R_�2i_�W^����`��e?333��R��$�X�D/  C�GÿP ?fff��> �-��ei�Q<����O �b}����Wy��o �o�o̵��Fo�o8�Y`F@ LuXa�U Y`Dz�PmtXoJ��jk�K�=� � (o:oLo^opo6��o� `�r��o�o8�� �� $�:�H�z�8�J�k��� ��Ə؏���� �b� �"���z�4���� ��:L^p���� 4y���E�����ӯ� ��	�ÿ-�?�ѿc��� ��������ϵu��0�Ϸ����xȘ��� �c�G}�;�X&�� ��\��Rq`������ m��� P�P ��� #�i  ����J��2�`V�����/�����>����Ħ�� �,�>�P�b�t�M��� �߼����ߞ���(� :�L�^�7���m�� ��������$�6� Z�l�~�������r�� ���� DV// z�����g/y/�/�%�2�l�/�/�/
?=�322.?W?i?{?�? �?�?�?�?�?�? t�n NE!e�Y�Z�ܝ�Y �Y��ϗ��i�O�O�O�OVd� )W�OP�I�!UWA3L>I��p_-g�\��}U>�L�P�Q�wB)<#�
�tp}_RY�8�VPB��L@ D�U4bU�U@��T H�`o/����fܚyo3&+Bu�U�o �o 2Vh`�>Ya�T_�O��CI�t$ �$%6>��R
��A�D���(���v5P+��̞t�.�����4Q$�敕��(4$�x��T�f�;��.ȅ�>��Hԅ4Q5{���8M�Y��<M=�P�4R��C�	:�S�>�w�b����� ��ɟ۟���noM�>�  �]� (b�T�b`l�T�LJY� -hx�������0�ů���PB�R��S@�?3�33<Ut�=T�I�aD�/  CaG�P_ ?fff<Q>%a �D@�`�X��(1��� `�hM<_6�d�@�� 5�(O���vϔ��F@ �Ŵ��\b��DzJ��Ĵ���x�p6��!�/�) ܄� ������̿����ϼ� ��8�JϔJ�\�n߀� �ߤ��ߔ������� "�4�F�X�j�|��l�~��������r��� �ϨϺ����������R �����/AS e��-�� �c�a/'�//%//����= I �i#���.�_~C��/ ��,��`��= ,e2�d Da�f9`�E�i|5? �P|$=!#�4�>e��%84$8�ro�<�?H>���4$Jd/v/ �/�/�/�/�/�O�/? ?*?X?�O`?r?�?�? �?�?�_�?�?�_O&O 8OJOlO&o�O�Oko�O �O�O�O__�o4_F_ X_j_|_bo�_�_��_�(l�1/����u2@R�0�B�T�f�w�V��2����ŏ׏��� ��1�C�U�\�S�v� �q�d���l8�<�<� 0rE�+�UW��!�N�E�j��d�p����(�����]a>�̯�g}���Is٥>L�"�	�IoӒhy<#�	
�Q�bpٯx���w�����]a�e�a�����`�@]��� ��g/d@�-o�8�տ�b`o�{B�a����[π|ώ�qϲ���wka�>���5�`�V���Itk$ 0�$��>�6�	
�b�A�b�
߄�x.�@֑�+������.����Ր�$�{����(4$��ռ����;��.$�>���H0吡5�=�@�8M�YL嘝�=	�h吢9qy��	 �߯����������%�7�I�[�j��$C�CSCH_GRP�13 2������&� �\�~E�y  <r���Y�� a�����������@+��B0����y>��?333�����ܙ�D/  �C�`G�P ?fff��>��ᔜ�	 ��_jx��W�ĝ�� �������el�����j2F@� %%1���2Dz � F$1#/��#���y �%7 I?mw/9?K?�� �_�/�/�/�/?!?S? O#ODO{?�?�?�?�? �?�?�?;O�O�OzOSO\��O�e_/%/7/ I/[/m/s_�R_d_o �_�_�_�_�_�_�oo o�o<o�o`oro�o�o �o�%��/~���(�qO�p�cɠ�V ��ޓe^�5U�)� 9R�p����%Ġ�Dƕ� ���j���g!��t�q������`�9���t���οa�s��>����t�����)� ;�M�&�q�������Տ w�ݏ���%�7�� [�m�F�������ǟ� ������3�E�W�i� ����Kϱ�ïկ��� ߿�/��S���|�@�R�d�z�2��߿�H���������2� 0�B�T�f�x���� ���������>�i	 i
^̵M�	�	���O�G �������������=�m�n�����.�ڱ>"qI��@R5R��V>L� �ƿ<P���<#�
m�MpV��2U����)���ڱ��u.��@�A�!r9�Ϭ� �B��l�JR�ݿ��BN�vr��/�//A/��� >2���x���/k�It$ �/-$��>��
�/�'Aj��/�/?�/�& �+���M5.��y�Y5$敕i5�(4$�u5-??;;���.�5>��H��55���58'M�Y�5�=� �5���?;	?,OO PO;G�?{O�O�O�O�O��OG���n�G  ��6p���  EU-U%�2QQ_c_u_��_	B�_�^)��+p<�u?333MR�Y��D/  C�:�G�P ?fff>�Z�u9i1a q���
_�b9}A�g =y/�o�o���{o��oOmʎ`F@ `�u�a�U5�`Dz#` �t�oQz�р�r� �]ooo�o�o�o k��o�����#m� #�5�G�Y�o�}���m� ���׏�����1� C�U���E�W�֟��i���K��o��� ��ϯi����z�� ����,�>���b�t� Ϙ�꿼�ο��<π�u:� ���������͟�"Ø�G��p� �W��Ϻߑ�b��� ��Ң��� �U��XǞ U���J@��g���V���?�K������>��� ���=�O�a�s߅ߗ� �߂��������1��� 9�K�]�o���l�� �������#�E�� Y�k�D���������� ���1CU; y�d/���
ߜ/�/�/�%2+|	??-?$??P=//h22c?�? �?�?�?�?�?�?
OO .O5t,~ONz!��Y�Z ��ii	"��./�0y�O�O'__CV��� ^W�O�I�!�Wv3��>~��_@-����"#�U>L�P�Q"�B�A)<#�
��p��_QR���PV�B����uy�Uib��U@6��T}o@/���f��oh9[+B ��U�o4UgJ��P:`>�ad9_/_���CIt$ 	�$�Z6>�b
�;�A��D;��]���jP+���̩�.������iQ$敕Ņ(�4$�х����;�{�.��>��H	��iQ5���8M�Y%�qM=�PA�iR!R�x�	o���s��� ���ן����"�4��oIM!�F�  "��]b2d�b:`�� ���J��bh����ѯ�Pe���讅B���cu�?333qU��rT|�I�aD/  C��G�P ?fffqQ>Za�Duŕ���� C(f�0͝Mq_k��� u7�I�j�]EO׿Q�x����F@ ��0�Q��b�Dz��Ā��ϭ�k��!�/�) ܹ�˿ݿ���� %�/����m���� �ߣߵ���������� ��3�E�W�i�{��������2����� E����������� %�+�R
�@R dv��T��b �F*<N�F���/\�6/H/Z/d�� )�r ~�iX�/�.�_ �C/?��a�p��r  ae=2�dyavn`�E�i �j?��P�$r!X�E4 �>9e�Z8i$m��oxL+O7H>���i$ 7J�/�/�/�/�/�/? �O)?;?M?_?�?/_�? �?�?�?�?�?�_O%O �_IO[OmOO�O[o�O �O�o�O�O_!_O_E_ i_{_�_�_�_�o�_ �_�o]l4/f/�
��2�2��e�w��������Ă2����� ��0�B�T�f�x��� �ĈΫ��q�d!�!�| m�q�q�erz�`����@D�V���z����d%�@��&�8�<��҃��>���}����~s�>LW�>�~o��yO<#�
%arp�ୢ��N���������e�a-�Ų�`E�@ ��F���ddu�bo@$�m�
��b�o�{Bq .�*ϐϱ��Ϧ������k��>�j�����L�^#�It$ e�$��K>�k�
Eߗ�A"����?߹�c�u�Ơ+�{���.�����š$敕!�(4�$�-�����;��=.Y�>��He�š�5��u�8M�	Y��͝=>���Ţnq����	��������� A�3�H�Z�l�~��������}��   qr�����9����� ݚ��	-?��(VD���s��?333ͥΤ��E�D/  C�`G�P ?fff͡>�����	�)o�x ������ͯ���� ����e��3�/<%zFF@ 9%E��FDz� Z$E�7/	/�X�8�*� �'9K]#?� �/M?_?��%o�/�/ �/?'?5?g?%O7OXO �?�?�?�?�?�?�?O@OO�O_�OgO!\��O /y_'/9/K/]/o/�/ �_!�f_x_2o�_�_�_ �_�_�_�oo,o�oPo �oto�o�o�o�o�%�`�/����(ȅO �p�cPɴ�j(�E�� yr�IU�^�MR�p�� ��Z�ձy�ʰ=�=�z ƏwV���q�������M���t���u�<����>����t�� ���+�=�O�a�:� ��������鏋��� �'�9�K�$�o���Z� ����ɟ۟�����#� ��G�Y�k�}�����_� ůׯ�����1�C� �g�����T�f�x���2����������	�� �2�D�V�h� z����������� ��2�R�}	}
r��M �	�	���O�G����� ��������Q����������B.�9�>�6q]��TRIR��j�>L� �ڿd���<'#�
��a�pj	pFU��=���9�@-�1��!B��@�A �5rM�����B��� �Jf ���Bb�� ��///C/U/�� >F������/�It$ �/$�>%��
�/�'A~��/��/?�/�&" +��=�a5.���m5!�$敕}5(4$�܉5A?S;;��.��5>��H�5!5����58M�Y�5)�=� �5!��
O0;	'?@O+OdOOG�? �O�O�O�O�O�O[�|�n�G  �� Jp��� YUAU9� FQe_w_�_�_B�_��^=��?p�-u?333)aR*m���D/  CN�GÿP ?fff)> n�-uMiEa����_ �bM}U�)#gQy-/�o "���o	c���`F@ �u�a	eI�`Dz7`�t�o��e#z�є߆� � qo�o�o�o�o��o� ����%7��7�I�[� m�����Ï������� ���!�3�E�W�i��� Y�k��ß}����_ կ������� }¯ԯ����
��.� @�R��v���Ϭ��� п����P��uN��0�� �����*� 6ìW�τޡk��� �ߥ�b���*��� �1�&���i�"� lǲ i�*�Z��{���V�!�%?_������>���!���Q� c�u߇ߙ߽߫ߖ��� ����E���M�_�q� ��������� �%�7�Y�m��X �����������! 3EWiO��x/ ���߰/�/�/�%�2?|?/?A?S?d=C/|22w?�?�?�?�? �?�?OO0OBOIt@~ cN�!��Y�Z�%�)i )i"2��B/Dy�O_;_2_WV�� rW�OP�I�!�W�3J>����_T-����6#�U>�L`�Q6�BU)<#�
��p�_eR��8/dV�B��J� ��U}b��U@J��T �©oT/-��f%��o|Mo+B��U�o Hi{^��dN`�>�a"dM_C_��CI�t$ �$n6>�#b
�O�A�DO���q��-�~P+��̞��.���Ʌ}Q$�敕م(4$�x兝���;��.��>��H�}Q5{��-�8M�Y9��M=�PU�}R&!f���	�������������� ��$�6�H�W��$�CCSCH_GR�P14 2����y�&�� \m.2�p)  )"��qbFd �bN`֥���Jávh⯀����y�/���B���+c��?333��Uޢ�T�I�aD/ � C�G�P ?fff�Q>na�D�� ʹ±�W(��D©ͱM �_���ɉl�~ϟ�q�YOφ�����F�@ �����b�Dz��3����Ϡ�1�/�) �� �� $�6���Z�d�&�8�� ����������� �� @����1�h�z��� ��������(�����g�@����z���R �� $�6�H�Z�`�R?Q u������ ��){M_q ��{ժ/��k/}/�/���^�� �y�� C/>�_�CR/K?"�� p&� uer2t�a1v �`�E�i��?�`�$ �!��z4�>Me&��8�$����oNL`OlH>����$lJ�/�/�/? ?(?:?_^?p?�?�? �?d_�?�?�? OO$O �_HOZO3o~O�O�O�O �O�o�O�O�o _2_D_ V_�_z_8�_�_�_�_ �_�o
oo�@o�li/ �/-�?�Q�g�2�̚������Џ����2 ��/�A�S�e�w��� �������Ľ����+t V�V�K|�������r�� �����y�������Ԧ*tZ��[�m�q��
��a>!6��}-8"�sC�>L��s�x�o=��y<#�
Za:rpC��������au
qb���pz�@��{�"&�� �d��oYƢ�?��b�o�{B;qc�_������� ���.��k˰>����ʯ����X�It$ Z��$�>���
z���AW���t��ߘߪ����+���:�.����F���$敕V�(4$�b��,��;��.��>��yH����5����O8M�Y���=s� �����q��	�	 �� �=�(�v�h�}����������4�ڝ���  �r# �ôn� ˰2��>P@bt��y�� y��%?333��:�F�z�D/  �C'pG�P ?fff�>�G�%& ^o�x���&-.�� �*)�����e֟�h�</Zz{F@� n%z�"�{Dz �$zl/>/���m�_� �J\n� �X?��/�?�?�/ Zo?"?4?F?\?j?�? ZOlO�O�?�?�?�?O O0OBO�O2_D_�O�OV\��O8/�_\/n/�/ �/�/�/�_V��_�_go �_�_�_oo+o�oOo ao�o�o�o�o�o�o�o )�%'��/����(ȺO�s����� ]�z�H����~U��� �R��΂��
����� r�r�Bz��Ew��B�����քT�ʵ���t���8Ϫ���Ș>����tȚ*�<�N�`�r� ����o���̏ޏ��� ��&�8�J�\�n���Y� ������ڟ����2� �F�X�1�|������� �֯������0�B� (�f�x�Qߜ�����ߛ߭���2,���H�,�=��U�2P� y������������ 	��"$.<�gчĲ	 �
���M��_�G �)����0����K������wc�#�>kq�-݉R~Rӟ>L� ��<��.�<#�
���p�>{U��=r���#�b�f��Vw��@#Q�jr�-��� R��J�U�&�H�B����!/B/T/7/x/�/=�'>{�&x�/��It$ �/-$G�>��
�/(7A��(?�/J?�/6W �+��̖5.��y��5V$敕�5�(4$ܾ5v?�;;���.�5>��H��5V5��E8'M�YE^�=� .EV��?Oe;	\?uO`O �O�G�?�O�O�O�O_�!_�6�~3W  �pJ�' �UvUn�{QO�_�_�_��_RB�_�^r��tp<bu?333^�R�_���D/  C���G�P ?fff^>G��bu�iza ��0�S_r�}��^Xg �yb/$6WJ�2��o�>����`F@ `�u�a>e~�`Dzl` �t�o��Xz���߻� ܦo�o�o�o�o ���ޏ��Zl�� l�~�������Ə���� ȟ� �2�D�V�h�z� ����������������2��
�����  ������	�ÿ-� ?�Q�c�u���Aϫ��� O��3���)�;υπ3���I�#�5�G�Q���_�k��EW�Ϲ� ���
��ڥNb�ޢ _�N*��f
&[�� ���W��� ��_�EZ@2��&�VG�V�Z?���$�>��� V�$��ߘߪ߼����� �����(�:�L�z� ��������� � ��6�H�Z�l���H �����������< 2�Vhz��� ���/�J!�S��/�/	?52t|R?d?v?$�?�=x/�22�?�? �?�?OO/OAOSOeO wO~tu~�N�!�ij ,Z�^i^iR"g�M�w/�yy1_C_p_g_�V��0�W_%Y)1�W�3>���_�-�ڢk#�U>LD`+ak�B��)<#�
�p��_�Rץ;/�V�B����e�b�2e@�3d���o�/Qb��OvZ��o���+B �e}�������`>�aWd�_x_�9�SIt$ R�$��6>�Xb
2���A�T��,���P�b��P+�����.�������Q$敕�(�4$��ҏ�;�{�.F�>��HR�޲Q5��b�8M�Yn��M=+`���R[!����	��џ���� ��.� �5�G�Y�k�}���o�MjΏ�  ^"���b{d&r�`� ҥ�Jס�h����,�P��C�1��B���`c��?333�U�T|�I2qD/  C��G�P ?fff�Q>�a�D��޹ֱ �(��y����M�_���� ��ϒϳϦ�O Ϛ�x��*3�F@ &�02����b3�DzȰGԀ2�$��ϴ�E1%?9 ���&�8�J�� n�x�:�L������ �������"�T��$� E�|������������<�����{�T�� ����f�&�8�J�\� n�tbSe�� ������ =�as�������/��/�/�/��� r�� �=y��W/>2o �Cf/_?6��Kp:�  �e�2Gt�afv�`*U*y ��?�C`�$�!���4 N�e:��8�$���oxbLtO�H>����$ �J�/�/??*?<?N? '_r?�?�?�?�?x_�? �?OO&O8Oo\OnO Go�O�O�O�O�O�o�O _�o4_F_X_j_�_�_ L�_�_�_�_�_�oo 0o	�To�l}/�/A�S�e�{�2�̮���ҏ�����2�1�C� U�g�y���������ӟ �������?tj�j�_| �������r�������@����̯ï�>tn�@�o�����/���a>#!J��}A6�sW�>L�����oQ��yO<#�
naNrpW����3���*�����auqv��/p��@ ��"":���d��o@mƶ�S�r�o �BOq w�s��������0�B��k߰>3���ޯԯ��^l�It$ ��$��K>���
����Ak���߈��߾��+�{��N�.���Z���$敕j�(4�$�v�.�@�;��=.��>��H����5����8M�	Y���=������q���	�-��Q�<� ��|�����������H������   �r7 �״��߰F. &�3�Rdv�
�(��*��, ��%?333�N�Z����D/  C;pG�P ?fff�>��[�%:2ro�x �:-B��>)� ��/u�|�P/<nz�F@ �%��6Dz$�$���/R/*����s� �^p���l?� �/�?�?/$/no$?6? H?Z?p?~?�?nO�O�O �?�?�?O O2ODOVO@�OF_X_�O�Oj\��O L/�_p/�/�/�/�/�/ �_j��_�_{o�_�_	o o-o?o�ocouo�o �o�o�o�o�o=�%;�`?���	8��O �#s�����q���`� ����U���R�� ₣���������Vz �Yw��V�����h�޵�����LϾ�<Пܘ>����ܚ >�P�b�t��������� Ώ����2�ԯ:�L� ^�p�����m���ʟ�� � ��$�F� �Z�l� Eϐ�����Ư��ꯨ� � �2�D�V�<�z��� e߰�����߯�����2,,
��.�@�Q�	0�i�2d���� ����������/�6$ -.P�{ћ��	�
��] 
�_W/�1)�� ��(D����_������ыw�7�>�q�AݝR�R#ӳ�>L� �#ϭ�B�<'#�
ʱ��p�Rp�U��Q����7�@v�z��j���@7Q �~r�A�	�R�� Z�i�:�\�B��� �5/V/h/K/�/�/Q�;>�:0�/��It$ 
?$[�>%�
�/<7A��<?��/^??6k +��=̪5.����5j�$敕�5(4$���5�?�;;��.��5>��H
Ej5���E8M�Y&Er�=� BEj�SOy;	p?�OtO�O�G�?��O�O�O_#_5_D[��$CCSCH_G�RP15 2����fQ&� \Z�]�  ғp^ 3�;�U�U���Qc �_�_�_ofBo
n�����pvu?33�3r�Rs���D/�  C��G�P /?fffr>[�� vu�i�aοD؈_1r�} ��r�g�yv/Yk��^�F��os���pF@ �uqse�pDz�` ����z8������ ��o�o �o#�GQ��%� ��ʿ����ŏ׏� ��-�����U�g�y� ��������ӟ�ïկT�-�笸g��?�� ��#�5�G�M��,� >���b�t��������� v�����h�:�L� ^�pϺ�h���~�X�j�|߆��K��Р�� zW0������?�8�� �b ���b_��z &o����ʌ����  �Ԕ�zZg���:f|肋�n?�;�M�Y�>�����Y������� ����'� K�]�o� ���Q���������� ��5�G� k�}��� ����}����� 1Cqg%/��� ����	�/-@V߈�?,?>?T52�| �?�?�?�?�=�/�22�?
OO.O@OROdO vO�O�O�O�t�~�N�! $CiCj8,���i�i�" �����/�yf_x_�_�_�V$G0�WH_ZY^1g�3�>��#o�-p���#0e>Ly`�`a�*R�)<#�
G'"p0o�R�p/�VR�����Oe�b ge@��hd�� �/����Fv��,���+B(!PeL��@��	����`>q��d�_�_n�ESIt$� ��$�6>��b
g���ADT��a�ۏ������P+���'�.����3��Q$�=�C�(4$�O����;��.{�>���H���Q5�����8M�Y���M=@``���R�!П��	� ��*��c�U�j�|��������!�M��ħ  �"��b�d [r�`���J��h+��=�O�a��x�f�R����c��?333��U'��T3YgqD/ � C G�P ?fff�Q>�a4T�� ��K�(䯮��] �_������������OU���)�G*h�F�@ [�g�ϵrh�Dz��|�g�Y�+���z1Z?L9 �7�I�[� m��E�ϭ�o���� ��G���!�3�I�W� ��G�Y�z��������� ����/�q�1����C���%ߛI�[� m�ߑߣߩCb�� T����� <N�r���� �/��?�ߴ/�/�/��ȧ�� �ry֧ �/J>go1S�/�?k߲ �po� �e�2|t�a�v �`_U_y/*�?2'x`/4 �!֪�4AN�eo��8�$��%�L�O�H>����$�J?)?;?M? _?q?�?\_�?�?�?�? O�_O%O7OIO[OmO Fo�O�O|o�O�O�O�O _�o3_E_i_{_�_ �_�_�_��_�_oo /oSoeo>��o�l�/ �/v�������2�㏐����*�	�B�2 =�f�x���������ҟ ������)�T�tt �����|�����r�� ���
�¯ԯ����st��8�������d�
P�q>X!��v8k�s��>Lհ��x�o���<#�
�a�rp��+�h�*�_���qOuSq��C�dpõ@ĴW"o�� �d���o������Br5�B�q�����/�A� $�e�w�*{�>h����	��ߡ�It$ Z��$4�>��
���A����7������D�+��̃�.������C�$敕��(4$ܫ�c�u��;��.��>��yH��C�5����O8M�Y��K�=�� �C��q,�R�	I�b� M���q�������������}�#��   �rl 7�ķ� �{c[�h<ȇ�@��?���_��a y�O%?333K���L�����D/  �CppG�P ?fffK�>4���O%o g�o�@
"o-w�K� Es)O�/#/D/7u��+/�/�z�F@� �%�+k��Dz Y�$��/�/E*ց���� ܓ��� ��?�	?�?�?G/Y/ �oY?k?}?�?�?�?�? �O�O�OOO1OCOUO gOyO�O�O{_�__�O�\�_�/�_�/�/�/ �/�/�/o���_�_�o o,o>oPoboto.�o �o<�o �o( r 5p�6?�"�4�>8�_L�Xs��2� ��ÿ������U;�� �RL�;����S���H� ���ɋzD��w԰��L��2
�����4�C��G�����>���C��s��������� ͏ߏ����'�9�g� 	�o���������ɟ�� ���ؿ#�5�G�Y�{� 5Ϗ���z�ůׯ��� )����C�U�g�y��� qϯ������7��@��������2a,?�Q�Hc�u��eߞ�2�� ��������
��.�@� R�d�k$b.�������	 �
��G]KK?�T_:W d�f)0]Ty���Д 	����l�>�q�v��R�RX��>L1X�<��w�<#�
���p���U(߆����l��ů����@lQ �r�v�>� OR<��GZ���oϑ�B��/j/�/�/�/�/�/��p>�Doxe&?��It$ ??-$��>�E
?q7A��q??�?=?O6� �+����5.��y��5�$敕�5�(4$�E�?�;;���.3E>��H�?E�5��OE8'M�Y[E��=wE�HшO�;	�?�O�O �O�GO_"_4_F_X_�j_��W~|W  K��p�h"p �U�U���Q��_�_o�o�B0on����p<M�u?333��R����!D/  C���G�P ?fff�>����u�i�a �y؜_fr�}����g �y�/m���{������ pF@ `�q�e� pDz�` 4����z2��� ��o%7 ��[e�'�9����� ��Ǐُ���A��� �2�i�{�������ß ՟�)�ׯ�h�A����{��S���%�7� I�[�a��@�R��v� ��������п����� ��*�|�N�`�rτ��π|��ߒ�l�~ߐߚ��_��д�*)�WD�� ��S�L�#��b8 '� �Зs�4$�S&� )�ʠ���0�ԨюZ@{���o'f����?��O�a�m�>��� ��m���������)� ;�_�q�����e ��������%��I� [�4���������� �����!3EW� {9/������ �/A�jߜ�.?@?R?h52�|�?�?�?$�?�=�/�22�?O 0OBOTOfOxO�O�O�O �O�t�~�N1,$WiWj L,���i�i�"�����/��yz_�_�_�_�V+$�[0�W\_nYr1gC�>�7o�-.�#��#De>L�`ta�>R��)<#�
[;"p�Do�R ��/�VR���%!ce�b {e@ȡ|d�'�/�����Zv��@���+B <!de`�����/���`> q�d�_�_���YSIt$ ��$��6>��b
{�͇A�XT͏u�����P+����;�.����G��Q$敕W�(�4$�c��-�;�{�.��>��H����Q5����8M�Y��]=t`ӕ�R�!�
�	���>� )�w�i�~�������Ư�5�M��ا  �"$��b�dor�`3� �Z ��h?�Q�c�u�P����z�R���c�?333e;�d|GY{qD/  C( �G�P ?fffa>�aHT�'��_ �(����'�/]o��+� ���������Oi���x=�[*|�F@ o�0{��#r|�Dz��Ԁ{�m�?��ʎ1n?`9 �K�]�oρϓ�Y� ���߃�����[� #�5�G�]�k��[�m� ������������1��C���3E����W� ��9߯]�o߁ߓߥ� �߽Wb��h�� �,�Pb� ������*/���(?���/�/�/��� ��0#�yꧠ/^>{o ES�/�?�p�0 �e�2�tq�v psUsy C*�?F'�`C41��4 UN�e���8�$��9x�L�O�H>����$ �J+?=?O?a?s?�?�? p_�?�?�?�?O�_'O 9OKO]OoO�OZo�O�O �o�O�O�O_3_�oG_ Y_2}_�_�_�_�_�_ ��_oo1oCo)go yoR��o�l�/�/������ą2���	��-�>��V�2Q�z��� ����ԟ���
�� #��=�h��t�����| �����r����@֯���1��t��@L���ʩ΁x�d�$q>l!��.�����>L�б��/�O<#�
�a�rp���?�|�>�s����$qcugq��W�xp׵@ $شk"��.��d�o@������Vr'I�B�q ����"�C�U�8�yߋ�>{(�>|���'����^��It$ ��$H�K>���
��)�A���)���K����X�+�{�̗�.������W�$敕��(4�$ܿ�w��;��=.��>��H��W��5���8M�	Y�_�=а/�W� �@�f�	]�v�a����� ����������"1��$CCSCH_�GRP16 2����S?&� \G�/>J�  ��  K� ���(���o�� Pȼ���S�	��s��u �c%?3�33_��`�����D�/  C�pG�P_ ?fff_�>H� ��c%���o1�u" �-��_�z�)c�F/X/ y/Ku3��`/�/�z�F@ �%�`��Dz�4��/�/pz*�ʏ�� �� ���/�?4/>? O O|/�/�o�?�?�?�? �?�?O�O�O_BOTO fOxO�O�O�O�O_�_�_A__�\�T_�/,o �/�/�/?"?4?:o�� o+o�oOoaoso�o�o �oc�o�oqU' 9K]�U5��k?E�W�i�s8�8_���s ��g�ێ׿��,�%� �Up�� b��O�L��� g��\�ϥ���zy��w �����g
T�Ҟ'� i�x�[��(�:�F�>���x�F����� ̏ޏ�����8�J� \�n���>�����ȟڟ ���׿"�4��X�j� |�����j�į֯���� ��0�^�T��x��� �������������πl�C�u���+�A�2@�,t���������2����	��-�?� Q�c�u������$�.�� ���00%�|]�� t҉_oW�ߛ)Se����4��5G	(K������>�q��b�R��>L�fM����<#�	
4��p��U]������������<���T@�QU�r  /��sĄRq�3&|Z/�¤���B�=9/�/��/�/�/�/?�˥>��y��[?2Itk$ t?$��>�z	
T?�7A1�?N?�?xr?�6� +���E�.��� E�$�{��0E(4$�<E��?K;��.hE>���HtE�5�=��E8M�Y�E���=M�E�}ѽO�;	 �?�O�O_WPOB_W_ i_{_�_�_/���~�W  ���p� �H"�e�U���Q� o*o<oNo�BeoSn�����p��u?33�3�b� 	T!D/�  C�G�P /?fff�>�! �u y�a8Ϯ��_�r � ��g��/�����Ű�B��4�UpF@ H�Tq�e�UpDz�`i�TF���z8g�G�9� �$6 HZl2����\�n� ��4����� �6� D�v�4�F�g����� ԟ���
��^�����v�0�������6� H�Z�l�~�����0u� ��Aϫ���Ͽ��� ��)�;���_ϱσϕ� �Ϲ�߱��Ǐ�߳���ψȔ�����_) �Wy�7�T�߁�X� �bm \������i$� �&�LL)����e ����Z��.��\f�����?/������>����Ԣ���(� :�L�^�p�I���� ���� ��$�6�H� Z�3~���i������ ��� 2/Vh z���n/��� 
/@R+?v�@����c?u?�?�52�| �?�?�?OM�//B2*OSOeOwO�O�O�O �O�O�O�O�t�~^A1 a$�i�j�,ح�i�i�" �˧�/�y�_�_�_�_
f`$�0%g�_�Y�1Qg=C�>E�lo=pc�X��#ye>L�`�a�sR9<#�
�p"pyobU��/fLR���<%@!�e0rQ �e@���dD�\ ?����vتu/" /";Bq!�e���@.��R�d�+p>Uq��d o�_���SIt$� Џ$!F>��b
���A�T���$�Ώ���1`+���p�.����|�0a$�=���(4$ܘ�P��b�;��.ĕ>���HЕ0a5�����8M�Y�8]=@�`�0b�!�?�	6� O�:�s�^�������ů�ׯ���j]���  �"Y�$r�d �rph�P�HZU�)xt��������,�����LR��N��c<�?333�8ep�9d|Y�qD/ � C] G�P ?fff8a>!q}T<� \�T��
8-���\�d] 8o2�`�<����1�$%�_���rߐ*��F�@ �հ��Xr��DzF��԰Ϣ�t�2��1�?�9 ܀ϒϤ� ���ώ����߸���4� FߐF�X�j�|��� �����������0� B�T�f�x���hz������n���ߤ� ����������b�� �+=Oa/ ��)/�/��/ /_/�]?#��/?!?+����90E#�y� �/�>�ozS�/�?�(� �p�90(uB�t@q�v 5p�U�yx*1O{'�`x4 91�D�N u��!H04�4�n�L�O�H>���04�J`?r?�?�? �?�?�?�_�?OO&O TO�_\OnO�O�O�O�O �o�O�O�o_"_4_F_ h_"|_�_g�_�_�_ �_oo�0oBoTofo xo^�o�o���o$|�/ -?��я���2N�,��>�P�b�s�R���2 ������ӟ���	�� -�?�Q�X�O�r����t ���|48�8�,�A 'Q�S���J�A�f��t쀁�������
��Yq>�!ȿc��8�E�յ>L��xEϢd�<#�
�a�rpտt���s�����Yq�u�q�����p�@YĠ"��c� +t<)��4
�ϋr\~�B�q����W�xߊ� m߮���s{]�>��1��\�R���It$ Z,�$}�>�2�
�^�A�^���*�<�ލ�+�����.�����匱$敕��(4$������;��. �>��yH,���5��<�O8M�YH���=� d���5�u���	��� ���������!3�EW��l�D.i  8�� ��U� � ]����������@������� y:Ø%?333������ة�D/  �C�pG�P ?fff��>}�٤�%� ��of��S"�-���� ��)��Z/l/�/�uh���t/�/�z F@�  5!t�� Dz �!4/�/�/�*���� ��� // $/�?H/R?O&O�/�/ �o�?�?�?�?�?�?.O �O�O_VOhOzO�O�O �O�O�O_�_�_U_._�\�h_�/@o�/ ?? $?6?H?No�-o?o�o couo�o�o�o�ow�o �o�i;M_q �i5��?Y�k�}��8�L_���s�{1� ��֣@�9�e�%� b����`�!Ԝ�@֑� ���z���w�Ԅ���{
h��\�}��������<�N�Z�>�����Z���Ώ���� �(��L�^�p����� R���ʟܟ� ��� 6�H�!�l�~�����į ~�د���� �2�D� r�h�&ߌ�����¿Կ ����
���.π�W����-�?�U�2�,���H���������2�� ��/�A�S�e�w��� �����$�.�����D D9ܐ]���ҝ_�W �߯)gy����H��I[	_�	����>�q$��bb��1>Lza��<+��<#�
H�(ҁp1�eq����������P�	�h@�Qi�r/�߇� �R��G&�Z-/�¸���B)�QM/�/�/�/�/
??�˹>!��x�o?FIt$ �?-$��>��
h?�7AE�?b?�?�?�6� �+���(E.��y�4E�$敕DE�(4$�PEOK;���.|E>��H��E�5���E8'M�Y�E��=a�E����O�;	�?_�O +_WdOV_k_}_�_�_�_"/���~�W  �����\"�  ee 
a�,o>oPo�bo�Byogn��<��u?333�(b��4	h!D/  C��G�P ?fff�>�5�uyq L����_�r���g ��/�������V��*�H�ipF@ `\�hq�e"ipDz�` }�hZ�,��z{�[�M� �8J\n� F����p�����H� ���"�4�J�X���H� Z�{���ğ֟���� �0�r� �2�����D��į&���J�\�n��� ������D����UϿ� ѿ�������=�O� ��s��ϗϩϻ���߀Ņ�ۏ�������Ȩ�����s)�W��K� h2�ߕ�l��b� p� �����}$��&�` `)0���3�y0����Z@��B��pf�����?�&/������>��� �Զ��*�<�N�`�r� ��]��������� �&�8�J�\�n�G�� ��}�������� � 4F/j|��� ��/��0/ Tf??������w?�?�?�52��?�?O$O+M
?CB2>OgO yO�O�O�O�O�O�O�O 	_��*^U1u$�i�j �,��i�i�"��ߧ	?���_�_o�_ft$��09g�_�Y�1egQC!>Yрo=w�l��#�e>L�`�a��R�9<#�
��"p��o,bi��/+f`R��!P%T!�eDre �e@��dX�p?������v쪉C"/6;B �!�e��0�B�%�f�x�++p>iq�do
o�ˏ�SIt$ �$�5F>��b
ď�A��T���8���E`+���̄�.������Da$敕��(�4$ܬ�d�v�;�{�.ؕ>��H��Da5����8M�Y �L]=�`�Db�!-�S�	J�c�N��� r�����ǯٯ�������$CCSCH�_GRP17 2����@�&� \4>|��79  �" m�8rt�rp����\Z ��=x����Ϳ߿@�����`R�b��cP�?333Le��Md�Y�q�D/  Cq GÿP ?fffLa> 5q�TPՑɉ��8b� �p�x]Log�t�P�3� E�f�8% _��Mߧߤ*��F@ ����M�lr��Dz{���������g��1�?�9 � ������������!�+� ����i�{ߤ{��� �������������/� A�S�e�w��������� ��.��A�� ���������!�' �b�<N`r ��P/��^/�B/ /&/8/J/�/B�q?X�02?D?V?`��%n0 z#�yT�
?�>�o�S? O�]��p�n0<u9B �tTq�vIp�U�y�*fO �'�`�4n1T�AD�Nu�VHe4H��\'_3X>���e43Z�? �?�?�?�?�?O�_%O 7OIO[O�O+o�O�O�O �O�O�O�o_!_�oE_ W_i_{_�_W�_�_� �_�_ooKoAo�eo wo�o�o�o��o�o�� Y|0?b?���.��2��a�s�����������2������� ,�>�P�b�t����Ԅ� ��ҁ�t���im� m�a�v\����@�R��v����t!���"�P4�8��Γ�q>�!�������z�
�>�LS�:�z���<#�
!q�p
ϩ��8J���ݢ���q�u �q)����pA�@�B� �"�Ϙ�`tq^ �i
��r���B�*�&� �߭߿ߢ����ߨ{���>��fđ���H��I�t$ a�$��>�g�
A��A���;���_�q�°+��̞�.������$�敕�(4$�x)�����;��.U��>��Ha���5{��q�8M�Y}�ɭ=:�����j�����	��������=�/�DVhz���$�CCSCH_GR�P18 2�����&�� \��v/��  m�� �� 5Ғ�٪��&�8J\��saݢ��� o��%?333�ɵ"ʴ�A�D/ � C�pG�P ?fffɱ>����% )!%����"�-�� ɿ��)�߰/�/�/�u���P/�/$?!�c F�@ V5b!���c Dz�w4b/T?&?�*T�4�&� �2/D/V/ h/z/@O�/�?jO|O�/ �/!�?
OO.ODORO �OB_T_u_�O�O�O�O �O__*_l_o,o�_�_>l��_ ?�oD?V? h?z?�?�?�oo�o O�o�o�o�o� 7I�m���� ���5��?����ӏ�8Ȣ_��sL�� ��E�A������fe� Z�jb뀹Ŷ�V���u� ��9�9�*��-�R�*� ��
��<���jӘ�����ϒ�����>���ℰ��$�6�H� Z�l�~�W�����Ɵ؟ ���� �2�D�V�h� Aό���w�¯ԯ��� ���.�@��d�v��� ��ȿ��|������ *��N�`�9���̭� ߏq����2 <������%��=�2 8�a�s����������� ����
4>$O�o� �����]�����_ �W�9����n���3��	��_
K��>S�z�qb8fb�Ӈ>L��x�ρ�<#�
��~�p�&ce��%Z���J�NѦ>"_о@a�R�j/� ���R�ϝ&�Z�/=��0�Bѧ�/	?*?<? ?`?r?%� >c!���?�It$ Z�?$/�>��
�?GA�O�?2O�?�6�?+���~E.�����E>$敕�E(4$ܦE^OpK�;��.�E>��yH�E>5���EO8M�Y�EF=� U>��'_MK	DO]_ H_�_lW�O�_�_�_�_��_	ok�$CCS�CH_GRP19 2���:a�&� �\.��1�  ��g�2"$�" �e eV
�a7(�o�o�o�oP:R�o�nZ�\��J�?333F�bG|�	�!D/  Ck��G�P ?fffF>/!�J��y�q�� �\o�j�rFawn� J?-�?�`�2��G�x�����pF@ Ӆ0�qGuf"�pDzup��я��a����� ܯ������ �%����c�u���u� ��������ϟ���ѯ �)�;�M�_�q��������鯗���(����� ;������ӏ���	� �!Ϛ ����6�H� Z�l�~ϐ�Jߴ���X� ��<�� �2�Dߎ�<��k�R�,�>�P�Z�� �h�t��)Ng��� ����Wr� �h� 6%3��$N!�&C ��) ��`������h�Nj;� ��%�fP�_�BO|/x!->���_� -
������������ ��1�C�U���%�� �����������	 �?Qcu�Q/� ��/��E; �/_q����/� ��?/S,*�\��? OO(E2}�[OmOO�O�M�?�B2�O�O�O __&_8_J_\_n_�_ ��~��^�1�$yz< c�gygy[2p�V��?��@:oLoyopo�f�$@@�go.i2A�g�C�!>���o�=��t3u>LMp4qt/�R�9O<#�
!�"p�b�D?�f�R����!�%�!#u�r� ;u@ ��<t����?Z$k�X/@�c� ��"�/�;B�! $u ���������ݏ��+�p>�q`t�o�oB�^cIt$ [�$�FK>�ar
;���Ad���5���Y�k��`+�{����.����޻a$敕�(4�$�#�۟�;��=.O�>��H[��a�5��k�8M�	Yw��]=4p���bd1��ʛ	��گů��� 7�)�>�P�b�t�������$CCSCH_�GRP1A 2������?&� \�>p�>�9  g2�� �r�t/��p����Z� �x �2�D�VϷ�m�[���R���is��?3�33�e��di;�D�/  C� G�P_ ?fff�a>�q d��� �/�8ٿ�� ���]�o����Ǐ�߼� �߯%�_J����:]�F@ P�\����r]�Dz��q�\�N� �p��NA.O I �,� >�P�b�t�:��ߢ�d� v�����/����(� >�L�~�<No���� ������ $f&�~8��� >�P�b�t���r }�I/����� /�/1/C/�/g/�/�/ �/�/�/?���?��?�?�?��Ȝ�0�# F�˷�??N;c�?�O `��T�d�0�u�BP� �qo��p3e3�$:�O'7 Lp$D�1˺�D6^�ud��H�4����\�_�X>����4�ZOO 0OBOTOfOxOQo�O�O �O�O _�o__,_>_ P_b_;�_�_q�_�_ �_�_o�(o:o�^o po�o�o�o�ov��o�o  $
�HZ3�~��|�?�?k�}�����2@��؟�������7�22�[�m������ ��ǯٯ������� I�i��ɔʉ������ ؂�����ٷ�ɿ����h���-Ǚ���(��Y�E��>M1t���k`��>L������{��<#�	
�qx�p�� �]���T����D�H���8�Y���@��L2 d���t�����
}�7��*�By��ŝ��$�6��Z�l��	�>�]�������Itk$ ��$)�>���	
��
�A��
���,�x����9�+���x��.�����8�$�{����(4$ܠ��X�j�;��.��>���H��8�5�=���8M�Y��@��=��8��!G�	 >�WB{f���������$C�CSCH_GRP�1B 2����4&� �\(��/+�  �a0,�Ԭ� 	БyP�~1؝�@��4��T��V0y��D5?333@��AĄ���D/  �Ce�G�P ?fff@�>)х�D5�) }!��V�"d=l�@� ['h9D�'?9?Z?,����/A?�?��� F@� �5�!A%`�� Dz o �4�/�?�?[:ˑ���� ܩ/�/�/�/ �/�O?O�O�O]?o? �oO�O�O�O�O�O�O �_�_�_#_5_G_Y_k_ }_�_�_�_�o�o"o�_�l�5o�?�?�?�? �?OO���o� 0BTfx�D�� �R��6���,�>� ��6Ee�LO&�8�J�TH�ob�n���H�� ���ς����eQ"�� �bb�0�-���H���=� ���١�Z�������b��H5�����J�Y��<�v�	��'�>���Y�'���������џ ���ο�+�=�O�}� υ�������ͯ߯�� ����9�K�]�o��� Kߥ�����ۿ���� ?�5���Y�k�}Ϗϡ� �����ϰ���M�$�V������"�2w<U�g�Hy�����{��2�� ������ 2DV hz�4x>�����) *�]ma)a)U�joPg z�|94Fsj����(,������>ʁ����b�bn��>LG .!n�<���<#�
��ҁp���e>����������%�"��5%@�a6$ɂ�/��T� ebR�6]j�/�҅ߧ�B��%?�?�?�?�?�?�?�ۆ >�!Z$�x{<OIt$ UO-$��>�["
5O�GA�O/O�OSOeF��+����E.��y�U�$敕U�(4$�U�O�K;���.IU>��H�UU�5��eU8'M�YqU�=. �U�^�_�K	�O�_�_ �_�W1_#o8oJo\ono��o�k�$CCSC�H_GRP1C �2����a�&� \���j���   a�ހ�"~$)2� u�e �
�a�(,>P�R(gU~��Ӏc#��?333�r��51D/  C��G�P ?fff�>�!����qߏ� �o|�����w��? ����׏�ՑD����<�W�F@ J�V��u�"W�Dz�pk�V��H��؊H�(�� �&�8�J�\�n�4��� ��^�p�ڏ����� �"�8�F�x�6�H�i� ����į֯�����@`�� ϟ�x�2̸�� ���8�J�\�n����� ��"wω�C߭Ͽ��� �������+�=���a� �߅ߗߩ߻�ﳕ��`ɟ�����јȖ� ����@9�g{�9�5/� ���Z��rN0^���% ��J4�!i6� --9� ��!�F ����j��0�%^v�����O�/�<��>�����
 ��*�<�N�`�r�K ����������� &8J\5/��k/ �����/"4 ?Xj|���p? ���//?B/T/ -Ox/�,����eOwO�O�E2��O�O�O_]	�?1R2,_U_g_y_ �_�_�_�_�_�_�_�� ��nCAc4�y�z�<ڽ �y�y�2�ͷ�?���o �o�o�ovb4�@'w��o�i�ASw?S�!>�G�n	Me�Z��3{u�>L�p�q�/ub
I<'#�
�!r2p{rpWŻ?vNb���!@>5B1�u2�S0�u@�� �tF�^�	O�$��/�� ںw�12?$KBs1�u �����0��T�f�;�>W��t�o���c�It$ ҟ$#V>%��r
���A�d�ଟ&�П�3p+��=�r�.���~�2q�$敕��(4$�ܚ�R�d�;��.�ƥ>��Hҥ2q5����8M�Y�:m=�p
�2r�1�A�	8�Q�<�u�`��������ǿٿ������$CCSCH_G�RP1D 2����.�&� \"N��%I  �2[�&� �t�����s�Jjx�+� �ϩϻ���.�����Nb��P��s>�?33�3:u��;t~i��D/�  C_0G�P /?fff:q>#�d >��wі/HP���^� fm:U�b�>�!�3�T�&5o��;��:��F@ ����;�Z���Dzi��������U�8�A�O�I ܣߵ� �����߱������� W�i�/i�{������� �������/A Sew��������/��/�� ���������/�r� /�/*/</N/`/r/�/ >?�/�/L?�/0??? &?8?�?0�_OF� O2ODON��\@h3�� B��?�N�|cO _� K�ˀ�\@*�'RǄB� �7��e���:T_�7�p �D\AB�/T�^���DX�SD6�p�lo!h>���SD!j�O�O�O �O�O�O�O�o_%_7_ I_w__�_�_�_�_ �_��_o�3oEoWo io�oE��o�o���o�o �o9/�Sew ���������G�@OPO�����2q� O�a�s�����u���2��ү�����,� >�P�b�t�{�r�� ���� �W[�[�O� dJt�v�.�@�m�d���߄����"�&��Ǽ�|�>�1�φ�p��h���>LA��(�h�򲇙<#�
��p�ϗ��8���˲��|��������Ѐ/�@|0��2�� ��N�_L��W�߮����B����z��@��������>���T��u�6��It$� O�$��>�U�
/���Aā�)���M��_���+�����.��������$�=�(4$������;��.C>���HO��5���_8M�Yk��=@(Ї��X����	�� ����+2D�Vhz��$CC�SCH_GRP1�E 2�����&� �\��d?��  [��0��x�#�� %�Ǻ���/&/8/�J/�a/O.˲��0<]ӻ5?333��"�����/�D/  C�܀G�P ?fff��>�����5�)�! ����v2�=㽷��' �9��?�?�?����>?�?O�Q0F@ `DEP1�%��Q0Dz�  eDP?BOO�:B�"�� � ?2?D?V?h? ._�?�OX_j_�?�?� �O�O
__2_@_r_0o Boco�_�_�_�_�_�_ ooZo�oro,|��oO�2ODOVOhO zO�O��q�=�� �������%�7� ɏ[��������������Eܟ�O�������HȐoِ�:�u�3� /�����}�Tu�"H�Xr ِ�դ�D��c��'� '��ѯ�@��ّ�@��*��X&��Д����߀�����>��� Д�� ��$�6�H�Z� l�Eϐ�����Ư���� ��� �2�D�V�/�z� ��e߰�¿Կ���� �.��R�d�vψ϶� ��j����������� <�N�'�r��ܛ�͟_�q�����2�<������$��+2&O as������ ��4�>=�]�)�* }��m�)�)���o�g���9����&\����!'����M'9��>A�h/�_rTr��u%>L� �!��o��<#�
��l�p�u/"Qu��&H����8�<�%,2M�%@�a�$@�X?����b��ߋ6�jq?+����B m�%�?�?O*OONO`O�� >Q1�$����O�It$ �O$�>��"
�O�GA���O�O _�O�F- +����lU.����xU,!$敕�U(�4$ܔUL_^[;�{�.�U>��H�U�,!5���U8M�Y�U4=� e,"��o;[	2_Ko6ooo Zg�_�o�o�o�o�o�o�{�$CCSCH�_GRP1F 2����(q&� \�|��  �� U� 2�$�2� �umuD rq%8����(b���~H�J��#8�?3334%�r5$x�1�D/  CY�GÿP ?fff4!> 1y8�y�q����J �X�`4/O�\�8O� -�N� ���5�����΀F@ ��́5�T2΀Dzc��͏�����O������ � ������ӏ叫�	�� կ�Q�c���c�u��� ������ﯭ����� )�;�M�_�q�����׿ �ϗ��￩̸)ϋ� ߯���ӟ���	�� �"�� ߺ�$�6�H�Z� l�~�8�ߴ�F���*� ��� �2�|�*�Y�@�0�,�>�H���V� b�9<w����/v� ����E��0��V�$5! �4<1�610��9��N �� ��V�<z)��%�v>M�0_j?�>���M�}� ������������� 1Cq/y�� ����/�	�/- ?Qc�??���? ���/3/)/�?M/ _/q/�/�/{?�/�/�O �/A<�J��O�O _U�2k�I_[_m__�]oO�R2�_�_�_�_o o&o8oJo\onou�l� �n�A�4���<Q�U� U�IB^�D�nOp�(:g^�v�4	P�w
Py Q�w�Sv1>�����M����bC�u>�L;�"�b?�b�I<#�
	1�2p��r��82O�v�b��v1�5 �1����0)�@v�*� ��Տ�OH4Y�F?�Q�2y?�KB�1�� t�������˟ݟ�;z��>΁N�yo0�sI�t$ I�$�V>�O�
)�{�At{�#��G�Y��p+��̞�.������q$�敕�(4$�x�ɯ۫;��.=��>��HI��q5{��Y�8M�Ye��m="����rRA����	��ȿ���׷%���,�>�P�b�tσ��$�CCSCH_GR�P1G 2������&�� \�N^�I  UB����r� �z�����j����߀ �2�Dߥ�[�I��b����W���?333�u
Ҳt�i)�D/ � C�0G�P ?fff�q>���d�� ����?�H��p����m ����鵟�����5��o8���	JK�F�@ >�J��тK�Dz��_�J�<����<Q_Y ��,�>� P�b�(���Rd�� ��	?����,: l*<]���� �� T//�l&,���~/,�>� P�b�t����/�k/}/ 7?�/�/�/�/�/�/�? ?1?�?U?�?y?�?�? �?�?���O���O�O�O��Ȋ�@�34��� oO-^)��c~Ow_N%�� B�R"�@���R>���]� ��!u!�J�_G:�T �A�ʦT$ny�RֻX�D����zl�o�h>����D�j�O__0_ B_T_f_?�_�_�_�_ �_��_oo,o>oPo )�to�o_��o�o�o�o ��(�L^p ���d���� � ���6�H�!�l����O �OY�k�}���2��Ư�د�����%�2  �I�[�m�������� ǿٿ������7�W� �ق�w������ƒ� ����Ϸ����� �V���ׇϙɝ�G�
3��>;Ab���Y"8N"ߓo�>L�П�xߏi���<#�
��f�po��K%���B����2�6���&�G���@���:BR��� ń�Ï���k�%����Bg��Ջ����$� �H�Z����>K�������ϭ���It$ Z��$�>���
����A�����������'�+���f.����r&�$敕�(4$܎FX�;��.�>��yH�&�5���O8M�Y�.�=�� �&�ϑ5	,E 0iT�������� +�$CCS�CH_GRP1H 2���"!�&� �\��?�  ҒO@��Ԛ���% g%>�l!�/�/�/�/P"�/�.B��D@��2E?333.Շ"/�|rɦ�D/  CS��G�P ?fff.�>�s�2Es9k1��  �D/�2RMZ�.�I7VI 2�O'OHO�ϵ?/Ox�O���0F@ �E0�1/5N��0Dz]0�D��?�O�OIJ������ ܗ?�?�?�?�?�_ O_�_�_KO]O��]_ o_�_�_�_�_�_�o�o �oo#o5oGoYoko}o��o�o��o�|� #�O��O�O�O�O�O _	��������0� B�T�f�x�2�����@� ҏ$�����,�v�$U�S�:_�&�8�BX� P�\���6'쟪��� p������u?2���rP� ����6���+��Ş� ��H����Џ�P�6*#� �����&8�G�*d�x��	��>���G� �w���������ѯ� ����+�=�k��s� ��������Ϳ���� ��'�9�K�]��9�� ��~���������-�#� ��G�Y�k�}ߏ�u�� �ߞ���;��D�������2eLCUgy�i��2��� �� 2DVh oDfN������)�*�� K}O9O9C�X>wh�jI@"/4/a/X/}&�� @�'/)�'�p�>���/z��r�r\��%>L501\��{�O<#�
���p�/��"�u,��&����p���5�2��#5@ pq$4���?z�B�Sr@�@FKz�?��s��B�� 5OnO�O�O�O�O�O��t0>�1H4s/i/*_^#It$ C_$�K>�I2
#_uWA $�u__�_A_SV� +�{���U.����Uޣ!$敕�U(4�$�e�_�[;��=.7e>��HCe�!�5��Se8M�	Y_e�=0{e�"L��o�[	�_�o�o�o�g o&8J\n}{��$CCSCH_�GRP1I 2�����q?&� \��X�>��  O�̐ �2l4Bt0�u�u��q �8��,�>��bU�C�ʿ���Q3��?3�33�%��$�#AD�/  C��G�P_ ?fff�!>�1 �������}��j� ϝ��/Ƈә�O���� ş��2�����E�F@ 8�D����2E�DzڀY�D�6��pƚ6	 �� &�8�J�\�"�����L� ^�ȟڟ�گ���� &�4�f�$�6�Wώ��� ��Ŀֿ����N���ߍ�f� ܸ���x� &�8�J�\�n������" e�w�1�߭߿����� �߯��+��O��s� �����������������Ȅ����� .I�wi�'#?�x�q Hռ�<@L���5�8D �1WF�0%I��� 40��z�s5L�����_�?t��>�������� *<N`9/�� ����/�& 8J#?n�Y?�� ����?/"/�?F/ X/j/|/�/�/^O�/�/ �/�/?�?0?B?_f?��<����S_e_w_�U2@��_�_�_�_m�Ob2oCoUogoyo�o �o�o�o�o�o��~ 1QQD|�|�qL��̉̉ �B�ϻ��O癟����vPD�P���y(�QA�-c�1>5�\���MS�H��Ci�>Lಀ���?cr�I<#�	
�1`Bpi��EթO�<r���1,E0A�� �A@��@����4� L��O�4�½?���e�B�?[BaA����럀���B�T�K�>�E�ń����~sItk$ ��$f>�Ƃ	
���A}t򯚯�x��Ц!�+���`��.���l� �$�{��|�(4$܈��@�R�;��.��>���H�� �5�=�е8M�Yܵ(}�=���� ��A	�/�	 &�?�*�c�Nǜ��ϣ������������$C�CSCH_GRP�1J 2�����&� �\^��Y  �BI��鄔� �y�a�8zf���ߗ�@�߻������<r�>�y΃,�?333(����)�ly��D/  �CM@G�P ?fff(�>�mt,�m� e�?�H>���L�T}(� C�P�,��!�B�E�o��)����J��F@� ����)�H���Dz W��������C��Q�_�Y ܑ����� ������E�W� �?Wi{���� ���/AS ew��y/�/
/��,�/��/������ ������?|��/�/�? ?*?<?N?`?r?,O�? �?:O�?O�?OO&O pOM_4_ _2_<�/JPVC��0��O �^��js�O�_�%9⹐ �"JP�b��0�Ԗ%� �u���JBo�G���TJQ�0�d�n����2hAT�$�^��lx>���ATzq_�_�_�_�_ �_�_�oo%o7oeo �moo�o�o�o�o�� �o�o֏!3EWy 3���x����� '��۟A�S�e�w��� o��������5�_>_Я���
�2_�=�O�Ha�s���c���2�� ��ҿ�����,�>� P�b�i�`��ή�Δ�� ���E-I�I�=�R/8' b�d��.�[�R�w�͔���������ת�j�>�A��t��"�"V���>L/��V�<��u�<#�
��ݒ�p�߅��%&��ֹ���j������⾐�@j!�B��t�<� M":���E*�m���Bޑ��h�����~�������n�>��B�m�xc�$��It$ =-$��>�C�
oA��o�;M���+����.��y����$敕��(4$���;���.1>��H�=��5��M8'M�YY��=�u��F���	��� ��/ /2/D/V/�h/w+�$CCSC�H_GRP1K �2����!�&� \���RO��   I��@��f��n��%�% ���!��??&?8?�(O?=>����@K�E?333���"���ɾ�D/  CʐG�P ?fff��>���ĩE�9�1�w� �/dB�M�ͥ��7�I�� �O�O�O��y�,O�O _<��?@F@ 2U>A�5��?@Dz�0ST>O�0__�J0��� �O O2ODOVOozO �_FoXo�O�O���_�_ �_
o o.o`o0Q �o�o�o�o�o�o�o@H���`��� �Or� _2_D_V_h_z_ ����_�q�+������� ˏݏ��%���I� ��m������ퟛUʯ`�_�������X�~ Ǡӓ(��'c�!���� r�k�B��26�F�Ǡ�� ��2���Q������ ��	�.��ǡ�*���m�F6�������n�<�ό�>������� � ��$�6�H�Z�3� ~�������⿄���� � �2�D��h�z�S� �ϰ������ϰ�
�� ��@�R�d�vߤߚ�X� �����������*�<� `�쉯��M_q�2�L����	��2=Oa s�������D �N .+K�v9v:k��} �9�9����w���I�/ �/�/�/�&J�z 7�{/�)�;7'��>�/�V?��M�B���c5�>L�0�1��]"��<'#�
z�Z�pc?2p?���66"����@&�*�5B;�5@�q �4.�FO�����r��yF �z_O���B[�5 O�O__�O<_N_��0>?A�4�/�/�_x#�It$ �_$>%��2
�_�WAw$�_��_o�_�V0+��=�Ze.���fe1�$敕ve(4$�܂e:oLk;��.��e>��H�e15����e8M�Y�e"-=�0�e2��)k	 o9$]Hw�o ������$[