��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����CCSCB2�_GRP_T � h $CO�MPMATEXP_1  :2F	�RIXU   d?$OFFSEAFGAGEsm;f�z� z_OKRGf � ��P��H FS_TYTS�BFRAMEe�$INIT_TO�L�RANGE2�_Ff�T�F�TRATIOe|� �H_LIMU��LFSOF�ST_S�mUP�S_����	e� O�L_{UDUMM�Y2U�3�N�� �$$CLA�SS  �������I��I�V�ERSION��  �5~�IRTUAL�ܻ' 2 �I�� �  � d����$g�A}נA������VA�.��1��dġ�C0�A,�]�@�����:���
*@��p������+A�A�����U�����A�K��A���C-���A�
��-7���EW\�� ��@��l@�����$6�A����@�u��=��h��@&\��9)��"07��)Hh�����@���@B'���\t���������{R���{_?P�A���/0@7a������>�k�	)>���B��B8��@��8����E�@1����1�#�c�@�LA �m��c	��!!����]B�y���gl^c��A/$�_uy�B��@T���.B?�=�@>vh�	C-��2�� �@;s�?ש�����	��W8��\�m�̮�����pB6#��B*�=B(z<�B/��?�q������@Y�@;��@U	)�@��@{m��@���  � A��A;��VARH�A �WB�H���I@/P��8�rn>�е0�������s� ��_�_k�۱0'B�����0@��0 ��F �B��02D-ADH � AE�0�0 �W@BpG��?��?�^����E?��a@n�_�B6�W@ �1�@���@	�@]�?ԥz�A\�T����>O��(�J8��