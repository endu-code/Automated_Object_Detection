��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CESS0s!_81s!J3�> �! � �$SOFT�T_�IDk2TOTAL7_EQs $�0�0�NO�2U SPI_OINDE]�5Xk2SCREEN_(4�_2SIGE0�_?q;�0PK_FI�� 	$THK�YGPANE�4 �� DUMMY1"dDDd!OE4LA!�R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Dc@�D5�F6�F7*�F8�F9�G0�G�G@JA�E�GbA�E�G1�G!1�G �F�G2�B!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HO30IO�0� }%�SMACRO�ROREPR�X� D+��0��R{�T UT�OBACKU��0 �)DE7VIC�CTI*0�A� �0�#�`B�S�$INTERVA�LO#ISP_UN9I�O`_DO>f7�uiFR_F�0AI�N�1���1c�C�_WAkda�jOF�F_O0N�DEL��hL� ?aA�a1bc?9a�`C?��P��1E��#sATB��d��MO� �cE' D [M�c���^qREV�BI�Lrw!XI� QrR�  � OD��P�q$NO�^PM�Wp�t�r/ "�w� �u�q�r�0�D`S p �E RD_E�pCq�$FSSBn&$CHKBD_SE^e�AG G�"$SLOT_��2=�� 	V�d�%��3 a�_EDIm  O � �"��PyS�`(4%$EP�1��1$OP�0�2��a�p_OK�UST1P_C� ��d���U �PLACI4!��Q�4�( raCOM9M� ,0$D�����0�`��EOWBn�IG�ALLOW� �(K�"(2�0VAARa��@�2ao�L�0;OUy� ,Kva�y��PS�`�0M_O�]����CCFOS_UT~p0 "@�1�3�#�ؗ`X"��}R0  4F IMCM�`O#S�`��Hupi �_�p�BA�!���M/ �h�pIMPEE_F�N��N���@O���r�D_�~�n�Dry�F� dCC_��r0  T� '��'�DI�n0"��pu�P�$I�������F�t XF� GRP0��M=q�NFLI�7��0U�IRE��$g"� S�WITCH5�AX�_N�PSs"CF_�LIM� �; �0EED��!���qP�t�`PJ_dVЦMODEh�.Z`��PӺ�ELBOF � ������p� ���3���� FB/���0�>�G� �>� WARNM�`/���qP��n�NST�� COR-0bF�LTRh�TRAT�PT1�� $AC�C1a��N ��r$�ORI�o"V�RT��P_S� CHG*�0I��rT2��1
�I��T�I1��>� x i#�Q\��HDRBJ; TCQ�2L�3L�4L�5L�6L�7L� N��9s!��O`S <F +�=�O��#92^��LLECy�"MULTI�b�"N���1�!���0T�� �STY�"�R`�=l�)2`����*�`T  |� �&$��۱m��P�̱�UT�O���E��EXT�����ÁB���"2Q� (䈴![0�������<�b+�� "D"���ŽQ��<煰kc1(�9�#���1���ÂM�ԽP��" q'�3�$ L� �E���P<��`A�$�JOBn�T���l�TwRIG3�% dK� ������<���\��+��Y���_M��7& t�pFLܐBsNG AgTBA�  ���M��
�!��p� �q��0�P[`��O�'[���0tnah*���"J��_R��CDJ��IdJ
k�D�%C�`�Z����0��P_�P��@ ( @F RO.��&��t�IT�c�NOM �
����S���`TE)w@���Z�P�d���RA�0��2b"�����
$T����MKD3�T��`U31����p(5!HGb�T%1�*E�7�c�KA�b�WAb�cA4#YNT|���PDBGD��2 *(��PUt@0X��W���AX��a���eTAI^cBUF���0!+ � �7n�PIW�**5 P�7M�8M�9
0��6F�7SIMQS�@>KEE�3PATn�^�a" 2`#�"��L64FIX!,C ���!d��D�2B�us=CCI�:FPCH�P:BAD�aHCE hAOGhA]HW�_�0>�0_h@�f�Ak���F��q\'M`#�"�DE3�- l�p3G��@FSOES]FgHBSU��IBS9WC��. `{ ��MARG쀜���FACLp�SLEWxQe�ӿl��MC�/�>\pSM_JBM��Ԁ�QYC	g�e#�w0 ā�CHN-�;MP�$G� Jg��_� #��1_FP$�!TCuf!õ#@�����d�#a��V&�0�r�a;�fJR���r�SEGFR�PIO�� STRT��N��cPV5���!41�r��
r>İ�b�B��O�2` + �[���,qE`&�,q`�y�Ԣ}t��yaSI!Z%���t�vT�s� ��z�y,qRSINF }Oбc���k��`���`�`L�ĸ T`7�C3RCf�ԣCC/�9���`a�uah�ub'�MI�N��uaDs�#�G�D
�YC��C�����e�0q0��� �EV�q�UF�_�eF��N3��s�ah��Xa+p,�5!�#1�!VSCIA?� A��s1�"!3 ��`F/k��_ �U��g��]��C�� a��s�.bR�4� �����N����5a�R��HANC��$L�G��P�f1$+@NYDP�t�AR5@N^�`�a�q���c��ME�108���}0��RAө�CAZ 𨵰�%O��FCTK��s`"��S�PFADIJ�O J�ʠ�ʠ���<����Ր��GI�p�B�MP�d�p�Dba��AcES�@	�K�W_���BAS�� �G�5 � M�I�T�C�SX[@@�!62�	-$X���T9�{s�C��N�`�a~P_H�EIGHs1;�WI�D�0�aVT ACϰ�1A�Pl�<����EXPg���|��C}U�0MMENU���7�TIT,AE�%)�a2��a��g8 P� a�ED�E.`��PDT��R�EM.��AUTH?_KEY  ����R�� �b�O	���}1ERRLH� �9c \� �q-�OR�D�B�_ID�@l �PU�N_O��Y�$SCYS0��4g�-�I��E�EV�#q'�P�XWO�� �: �$SK7!f2&�T�d�TRL��; ��'AC�`��ĠINMD9DJ.D��_��bf1��f���PL�A��RWAj���SD��A��!+r|��U�MMY9d�F�10�d�&���J�<��}1P�R� 
3�PO9S��J�= ��$V$�q�PLB~�>���SܠK�?�����CJ�@����EN5E�@T��A���S�_�RECOR��B�H 5 O�@7=$LA�>$~�r2��R��`�q�b`�_DLu��0RO�@�aT[� Q��b������! }О��PAUS���dE�TURN��MR�U�  CRp�E�WM�b�AGNAL:s2$LA�!�?$PX�@$P�y A �Ax�1C0 #ܠDO�`X��k�W�v�q�GO_A7WAY��MO�ae����]�CSS_C�CSCB C �8'N��CERI����J`u�QA0�}���@�GAG� R �0�`��{`��{`OF�q�5��#kMA��X��&���LL�D� �$���sU�D)E%!�`���OVR10�W�,�OR|�'�$�ESC_$`�eDSGBIOQ��l �\�B�VIB&� �c�,�����f�=pSS�W���f!VL��P�L���ARMLO�
��`����d7%SC �bALspH�MPCh �Ch �#h �#h 5�UU���C �'�C�'�#�$'�d�#AC\4�$�pH��Ou�0�!Y��!�SB�� �`k$4�C�P3Wұ~46$VOLT37#$$`�*�^1�0�$`O1*�$o��0�RQY��2b4�0DH_THE����0xSЯ4�7ALPH�4�`���7�@ �0�qb7�rR�5�88� �×���"��Fn�MӁVHBPFUBAFLQ"D�s�`�THR��i2dB�����G(��PVP�����(������1�J2�B�E�C�E�CPSu�Y@� �Fb3���H�(V�H:U �G�
X0��FkQw�[��Na�'B���C IN{HBcFILT�� �$��W�2�T1�[� ��$���H Y6АAF�sDO��Y �Rp� fg�Q�+�c�5h�Q�iSh�QPL��Wqi�QTMOU �#c�i�Q\��X�gmb���vi�h�bAi�fI��aHIG��ca	xO���ܰ��W�"vAN�-u!��	#AV�H!Pa8$P�ד#p��R_:�A�a��B��N0�X�MCN`���f1[1�qVE�p��Z2;&f�I�QO�uh�rx�wGldDN{G|d��aF>!�9�r�aM:�U�FWA�:�Ml���X�Lu��$ !����!l�ZO�����0%O�lF�s�13�D	I�W�@��Q����_��!CURV�A԰0rCR41ͰZ �C<�r�H�v���<�`0��<�(�f�CH�QR 3�S���t���Xp�VCS_�`�ד�F���ژ���?N�STCY_ E L����1�t�1�T�U��24�2B�NI �O7������DEV�I|� F��$�5�RBTxSPI2B�P���BYX�����T��HNDG>��G H tn���L��Q�C���t5��Lo0 H���閻�FBP�{tF�E{�5�t��T��I��DO���uPMC�S�v>�f>�t�"HOTSW�`s�CP�wELE��J T��@�e�2��25�� O� ��HA7�E��344�0�LN���A�K �� MDL� 2J~PE��	A��s��tːÈ�s�JÆG!�rD"�ó�����\�T�O��W�	��/��S�LAV�L  �0INPڐ���`%��_CFd�Mw� $��ENU��OG��b�ϑ]զP�0�`ҕ�]�IDMaA�Sa��\�WR�#���"]�VE�$a�SKI�STs��sk$��	2u���J�������p	��Q���_SVh�EXCLUMqJ2M!'ONL��D�Y��|r�PE ղI_V��APPLYZP��HcID-@Y�r�_M�2=��VRFY�0��xr�1�cIOC_f�D�� 1������O���u�LS���R$D_UMMY3�!��z�S� L_TP/B�v�"���AӞ�ّ �N ���RT_�u�� �G�&r[�O D��P_;BA�`�3x�!F ��_5���H����� �� �P $�KwARG�I��� q�2O ���SGNZ�Q� �~P/�/PIGNs�l�$�^ sQ|ANNUN�@��T<�U/�ߴ�LA@zp]	Z�d~
��EFwPI�@ Rk @�F?IT�?	$TOTA%��Pd���!�M�NIY�S+���E��A[�
DAYS\�ADx�@��	�� �EFF_AX�I?�TI��0zCO�JA �ADJ_�RTRQ��Up���<P�1D �r5̀Ll�T�0? ]P�"�p��mtpd��V �0w�G���������SK�SU� ��CTRL_CA��� W�TRAN�S�6PIDLE_�PW���!��A�V曧V_�l�V ��DIAGS���X�� /$2�_SE�#TAC���t!`�!0z*@��RR��vPA���p ; SW�!�!�  ��ol��U��oOH��P�P� ��IR�r��BcRK'#��"A_Ak� ��x 2x�9ϐZs2��%l�W�0t*�x%oRQDW�%MSx��t5AX�'�"��LI�FECAL���10��N�1{"�5Z�3�{"dp5�ZU`}�MO�TN°Y$@FL9A�cZOVC@p�5�HE	��SUPP!OQ�ݑAq� Lj (CL�1_X6�IEYRJZRJWRJ�0TH�!UC|��6�XZ_AR�p6��Y2�HCOQ��MSf6AN��w$��ICTE�Y `>��CACHE�Cp9�M�PLAN��oUFFIQ@�Р�0<�1	��6
���MSW�EZ 8>�KEYIM�p��TM~�SwQq�wQ�#���TROCVIEܻ �[ A�BG�L��/�}�?� 	��?��D\p�ذST��!�R� �T� ��T� �T	��PEMA�If�ҁ��_F�AUL�]�RцĆ1�U�� �TR�E�^< �$Rc�uS�% IT��BUFW}�W��9N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTT(����sP��M��Ot�T�LwAX � ��XX~`9#�c_G�3
ЧYN_1�_�D���1 �2M�*��T�F��H@ ~g�`� 0p���Gb-sC_R�AIAK���r�t�RoQ8�u7h�qDSPq��rP��A�IM�c6�\����s2�U�@�A�s�M*`IP���s�!D��6�TH�@n�)�OyT�!6�HSDI3��ABSC���@ V`y��� �_D�/CONVI�G��H�@3�~`F�!�pd��psqSCZ"���sgMERk��qFB��Lk��pET���aeR�FU:@DUr`����x�CD,���@p;cJHR�A!��bp�ՔՔ+PSԕCʭ��C��p;��ғSp�cH *�LX�:cd�Rqa� | ����W��U��U�@�U�	�U�OQU�7R��8R�9R��0T�^�1�k�1x�1��1��1���1��1��1ƪ2RԪ2^�k�2x�2��U2��2��2��2��U2ƪ3Ԫ3^�3k�Bx�3���o���3���3��3ƪ4Ԣ]�EsXTk!0�d <�  7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr�����.�2REM� Fj��B�OVM��A�T7ROV�DT�`-�MX<�IN��0,�NW!INDKЗ
w�<׀�p$DG~q3�6��P�5�!D�6�R�IV���2�BGEA-R�IO�%K�¾DN�p��J�82�PB@>�CZ_MCM�@�1���@U��1�f ,<②a? ���P�I�!?I�E���Q����`m���g�� _0Pfqg RI�9ej�k!UP2_ gh � �cTD�p@���! a�����wBAC�ri T�Ph�b�`�) OG���%���p��IFI��!�pm�>��	�PT��"��MR2��j ��Ɛ+"�� ��\��������$�B`�x%��_ԡ�ޭ_����� M������D�GCLF�%DGDMY%LDa��5�6P�ߺ4@��Uk���? T�FS#p�Tl P���e�qP�p$EX_����1M2��2� 3�5���G ���m ���Ѝ�SW�eOe6D�EBUG���%G�R���pU�#BKUv_�O1'� �@PO�I5�5�MS��OOfswSM��E�b�@�0�0_E n �0~�� �TERM�yo�C��ORI+���p�D  �S#M_���b�q�����TA�r�����UP�Rs�s -�1�2n$�>' o$SEG,*> �ELTO��$U�SE�pNFIA�U"4�e1���#$p$UFR���0ؐO!�0̫���OT�'�TA�ƀU�#NST�P�AT��P�"PTH	J����E�P r�PV"ART�``%B`�ab�U!REL:�aSH�FT��V!�!�(_SEH+@M$���� ���@N8r����OVR�q��rSHI%0��UzN� �aAYLO����qIl����!�@��@ERV]��1�?: �¦'�2��%��5��%�RCq��EASY1M�q�EV!WJi'���}�E���!I�2��U�@D��q�%Ba��
5P�o��0�p6OR�MLY� `GR��t2b 5n� � ��UPa�U�u Ԭ")���T�OCO!S�1PO�P ��`�pC��������Oѥ`REPR�3��aO�P�b�"e�PR�%WU.X1��eo$PWR��IMIU��2R_	S�$VIS��#(AUD���Dv"w v��$H���P_ADDR��H��G�"�Q�Q�QБR�~pDp1�w H� S Z�a��e�ex�eƅ�SE��r��HS���MNvx� ���%Ŕ��O�L���p<P��-��A�CROlP_!QND�_C��ג�1�T �R'OUPT��B_�Vp	Q�A1Q�v��c_� �i���i��hx��i����i��v�ACk�IOU��D�gfsu^d��y $|�P_D���VB`bPRM_��b�HTTP_�אHaz (��O�BJEr��P��$���LE�#�s`{� � ��u�AB%_x�T~�S�@��DBGLV��KR�L�YHITCOU��BGY LO a�TEM��e�>�+P�'�,PSS|�P�JQ�UERY_FLA��b�HW��\!a|2`u@�PU�b�PIO��"�]�ӂ/dԁ�=dԁ�� �IOLUN��}����CXa�$SLZ�$I�NPUT_g�$�IP#�P��'���SLvpa~��!�\�W�C�-�B%�IO�pF�_ASv��$AL ��w �F1G�U��B0m!���0H�Y��ڑ��i᎐UOPs� `������@[�ʔ[�і"�[PP�S�IP�<�іI�2���P�_MEMB��i`� X��IP�P�b{�C_N�`����R0�����bSP��p�$FOCUSBG�a~�UJ�Ƃ �q  � o7JOG�'n�DIS[�J7�cVx�J8�7� Im!|�)�7_LAB�!��@�A��APHI�b�Q�]�D� J�7J\���� _KE}Yt� �KՀ�LMONa����$XR��ɀ��WATCH_��3���EL��}Sy~���s� �Ю!V�g� �CTR3򲓥��LG�D� �R��I�~
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�Gȴ I�F�%SO���q �Ɩ�@��v��ƴ��K�S�����w�k�N����E��\���'�"*�U�s5��@L>�4�7DAUZ�EA�pՀX�Dp�f�GH�B��OGBOO��g� C���PIT����� ��REC��S'CRN����D_p�b�aMARGf�`��@:���T�L���S�s¡�W�Ԣ�Iԭ�JG=MO�MNCH�c���FN��R�Kx�PR�Gv�UF��p0��F�WD��HL��STP��V��+���Є�RS��H�@�몖C�r4��?B��� +�O�U �q��*�a28����Gh�0PO������b��M8�Ģ��EX���TUIv�I��(� 4�@�t�x�J0@J�~�P��J0��N�a��#ANA��O"�0V�AIA��dCLEA�R�6DCS_HIP"�/c�O�O��SI��S��I�GN_�vpq�uᛀTܓd� DEV-�LL�A �°BUW`�j�x0T<$UǃEM��Ł�����A
�R��x0�σ�a��@OS1�2�3�a�`� ��ࠜh�AN%-���-�IKDX�DP�2MRO�X�Գ!�ST��Rq��Y{b! �$E&C+��p.&A&q���`� L���ȟ%Pݘ��T\Q�UE�`�Ua��_ � �@(��`�b���# �MB_PN@ �R`r��R�w�TRIqN��P��BASS��a	6IRQ6�M�C(�� ��C�LDP�� ETRQ�LI��!D�O9=4FALʡh2�Aq3zD᱌q7��LDq5[4q5ORG�)�2�8P�R���4/c�4=b-4�t�� �rp[4*�L4q5SB�@TO0Qt�0*D2FRCLMC@D�?�?�RIAt,1ID`�D� Yd1��RQQprp�DSTB
`� �F�HAXD2���G>�LEXCES?R��R�BMhPa�͠�B�D4�E�q`�`�F_A�J�C[�O�H:� K��� \���b2Tf$� ��LI�q�SREQUIRE�#�MO�\�a�XDEB�U��,1L� M䵔 �p���P�c�AA"RN��
Q�q�/�&����-cDC��B�IN�a?�RSM�Gh� �N#B��N�iPST�9� � 4��L�OC�RI���EX�fANG��A,1�ODAQ䵗�@1$��9�ZMF���� �f��"��%u#ЖVgSUP�%d�FX�@�IGGo�� � rq�"��1��#B��$���p%#by��rx���v<bPDATAK�p!E;����R��M��*�� t�`MD�qI���)�v� �t�A�wH8�`��tDIAE��sANSW��th��
�uD��)�bԣ(@$`�� PCU_�V06�ʠ�d�PLOr�$`��R���B���B�pp�����,1RR2�E��  ��V�A�/A d$CALII�@��G~�2���!V��<$R�S�W0^D"��ABC~�hD_J2SE�Q\�@�q_J3M�
G�G1SP�,��@PG�Bn�3m�u�3p�@���JkC���2'AO)IyMk@{BCSKP^:�ܔ9�wܔJy�{BQ�ܜ�����`_A1Z.B��?�EL��YAOCMP�c|A)���RT�j���1�ﰈ��@1�������Z��SMG��pԕf� ER!��a[INҠACk�p�����b�n _���@����D�/R��3DIU��CDH�@
�:#a�q$V�Fc6�$x�$���`�@���b��̂�E��H �$BEL�P����!ACCEL����kA°IRCS_R�pG0�T!��$PS�@B2L`���W3�ط9�< ٶPATH��.�Dγ.�3���p�A_ ��_�e�-B�`C����_MG�$DDx��ٰ��$FW�@��p����γ����DE���PPABN�R?OTSPEEup��O0��DEF>Q���`$USE_���JPQPC��JYh����-A 6qYN�@�A�L�̐�L�MO�U�NG��|�OL�y�INCU��a���ĻB��ӑ�AENCS���q�B�����D�IN�I�����pzC��VE�����23�_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��PR9C����MOS� gT�MOpp�@-GPERoCH  M�OVӤ �����!3�yD!@e�]�6�<�� ʓA����LIʓdWɗ��:p83�.�I�TRKӥ�AY����?Q^���m��b��`p�CQ�� MOM�B?R�0u��D����y�0Â��DU�ҐZ�S_BCKLSH_C����o�n� ��TӀ���
c��CLALJ��A��/PKCHKO0�SNu�RTY� �q���M�1�q_
#c�_U�MCP�	C���SC�L���LMTj�_AL�0X����E� � �� ���m�0h���6��PC����!H� �P�ŞCN@�"sXT����CN_��1N^C�kCSF����V6����ϡj���nnCAT�SHs �����ָ1���֙����������PA���_	P���_P0� e���0O1u�$xJG� P�{#�OG���TORQU(�p�a�~���`�Ry������"_W�� ^�����4t�
5z�
5UI;I ;Iz�F�``�!��_8�1��VC��0�D�B�21�>	P�?�B�5JRK�<�2�6~i�DBL_SM�Q:&BMD`_DLt�&BGRV4
Dt�
Dz���1H_���31�8JCcOSEKr�EHLN�0 hK�5oDt�jI��jI<1�J�LZ1�5Zc@y��1cMYqA�HQBTHWM�YTHET09�N�K23z�/Rn�r@C�B4VCBn�CqPASfaYR<4gQt�gQ4V�SBt��R?UGTS���Cq��a��P#��<�Z�C$DUu ���R䂥э2�Vӑ��Q��r�f$NE�+pI�s@�|� �$R�#QA�'UPeYg7EBHBALP!HEE.b�.bS�E�c �E�c�E.b�F�c�j�F�R�VrhVghd��lV��jV�kV�kV�kV*�kV�kV�iHrh�f��r�m!�x�kH�kH��kH�kH�kH�iOJclOrhO��nO�jUO�kO�kO�kO�kO�kO�FF.bTQ����E��egSPBAL�ANCE��RLE6�PH_'USP衅F���F��FPFUL�C�3��3��E��1=�l�UTO_p �%�T1T2t���2N W�����ǡ��5�`(�擳�T�OU���>� INSEG��R��REV��R���DI�FH��1���F�1�;�OB��;C���2� �b�4LCHgWAR��;�ABW!~��$MECH]Q��@k�q��AXk�P���IgU�i�� 
p���!����ROB��CR��ͥ#*�C���_s"T � �x $WEIGHh�9�$cc�� �Ih�.�IF ќ�LAGK�8SK��K�7BIL?�OD��U�&�STŰ�P�; �����������
�Ы�L��  2��`�"�DEBU.�L�&�n��PMMY9���NA#δ9�$D&���$��� Qw �DO_�A��� <	���~�H�L�BX�P�N�Ӣ+�_7�L�t�OH  ��� %��T����ѼT�����TgICK/�C�T1��%������N��c����R L�S���S��ž��PROMPh�E~� $IR� �X�~ ���!�MAI��0��j���_9�����t�l�R�0CO�D��FU`�+�ID�_" =�����G_�SUFF<0 h3�O����DO�� ِ��R��Ǔن�S���P�!{������	�H)��_FI��9��O�RDX� ����3�6��X�����GqR9�S��ZDTD���v�ŧ4 =*�L_NA4���|K��DEF_I[� K���g��_���i���0��š���IS`i  �萚����e��"��4�0i�Dg����D� O��LOCKEA!uӛϭ�0����{�u�UMz�K� {ԓ�{ԡ�{����}� ��v�Ա��g����� ��^���K�Փ����!w�N�P'���^����,`�W\�[R��7�TEFĨ ��OULOMB�_u�0�VIS�PITY�A�!O>Y�A_FRId��F(�SI���R��H����3���W�!W��0��0_,�EAS%��!�& �"���4p�G;穯 h ��7ƵC?OEFF_Om��H�m�/�G!%�S.��߲CA5����u�G�R` � � �$R� �X]�TME�$R�s�Z�/,)ËER�T;�:䗰��  ]�LL��S��_SV�($�~����@���� �"SETU��MEA��Z�x0�u���>��� � � �� ȰID�"���!�*��&P���*�F�'����)3��#�A��"�5;`*�ЧREC���!7�S�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I���0�MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X17ࡐMO�R�� H	�CU �A3�z�1Q�
��3���$��FV���2ՠ�AbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų7�=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	����y�7�t�#�}1� @�@;���O&E�RI#A��
N�ЈX�s�f�{��PL�}1�,RTv�m�AT�USRBTRC_T(qR��B �����$� �Ʊ��,�~0� D��`-CSALl`�SA0���]1gqXE���%���C��J�
���cUP(4����PX���؆�q��3�w� ��PG�5� $SUB�������t�JMPWAITXO��s��LOyCFt�!D=�CVF	ь�y�⻑R`�0��CC_�CTR�Q�	�IG�NR_PLt�DB�TBm�P��z�BW�)����0U@���IG��a��Iy�TNLND��Z�R]aK� N��B�0�PE�s���r���f�SPD}1� L�	�A�`gఠ�S��U!N�{���]�R!�B�DLY�2���D�B:�PH_PK��E��2RETRI�Et��2�bsR���FI�B� ����8�� 2��0DBG�LV�LOGSIYZ$C�KTؑUy#2u�D7�_�_T1@�EM�@C\1A�����R��D�FCHEC�KK�R�P�0���2�@&�(bLEc�" �PA9�T���P�C�߰PN�����AR@h�0���Ӯ�PO�~�BORMATTna F�f1h���2�S��SUXy`	�3�LBо�4�  rEI�TCH����8PL�)�AL_ � �$��XPB�q� C�,2D�!��+2�J3�D��� T�pPD�CKyp��oC� _AgLPH���BEWQo���� ��I�wp� � �b@PA�YLOA��m�_1�t�2t���J3AR���؀դ֏�laTI�A4��5��6,2MOMCP�����������0BϐAD�����\���PUBk`R�Ԑ;���;�����z4�` I$PI\D s�oӓ1yՕ�w�2�w�UZ��I��I��I�〛�p����n���y��e`�9S)bT�SPEED� G��(�Е�� /���Е�`/�e�>���M��ЕSAMP��6V��/���ЕMO�@ 2@�A��QP�� �C��n����������� LRf`kb�ІE9h�EIN09��7S.�В9
yPy�GA�MM%S���D$GGET)bP�cD]Ԛ�2
�IB�q�IN�G$HI(0;A��$LREXPA8)LWVM8z�)��g���C5�C�HKKp]�0�I_��h`eT��n�q���eT,���� ��$�� 1��iPI� RCH_D`�313\��30LE�1��1\�o(Y�7 �t�M�SWFL �M��SCRc�7�@�&��%�n�f�SV���P�B``�'�!�B�sS_�SAV&0ct5B3NO]�C\�C2^�0� mߗ�uٍa��u���u:@e;��1���8��D�P ���������)� �b9��e�GE�3���V�e�Ml�� � �YL��QNQSRlbfqXG�P �RR#dCQp� �S:AW70�B�B[�CdgR:AMxP�KCL�H����W�r�(1n�g�M�!o�� �F�P@}t$WP�u�P r�� P5�R<�RC�R�� %�6�`��� ��qsr %X��OD�qZ�Ug��ڐ>D� ��OM#w�J?\?n?�?�?���9�b"�e�]�_��� |��X0�� bf��qf��q`�ڏgzf2��Eڐ� d�FbJ�"�0���FdPB���PM�QU�� �� 8L�QCO�U!5�QTHI�H�OQBpHYSY�ES��qUE�`�"�]O���  �P�@L\�UN���Cf�9O�� P��Vu���!����OGRA�ƁcB2�O�tVuI�Te �q:pINFOB�����{�qcB�e�OI�r� (�@SLEQS��q��p�v�gqS���� 4�L�ENABDRZ�PTIONt�����Q�\��)�GCF��G��$J�q^r�� R���U�g������_ED����� ��F��PK��E�'NU߇وAUT<$1܅COPY���(��n�00MN��^�PRUT8R ��Nx�OU��$G�[rf�2�RGADJ����*�X_:@բ�$�����P��W��P���} ��)�}�EX��YCDRz�~�NSr.��F@r�LGO��#�NYQ_FREQR�W� �#�h�TsLAe#����ӄ ��CRE� s�IFl��sNA��%a��_Ge#STATUxI`e#MAIL�� ���q t��������ELEM�� �|/0<�FEASI?� B��n�ڢ�vA�]� � I�p��Y!q�]�t#A�ABM���E�p<�VΡY�BASR�Z��S�UZ��0�$q���RMS_TR;�qb ���S�Y�	�ǡ��$���>C��Q`	� 2� _�TM������ ̲�@ �A��)ǅ�i$'DOU�s]$Nj����PR+@3���rGR�ID�qM�BARS� �TY@��OTO��p��� Hp_}�!Ⱦ���d�O�P/�� � �p�`PORp�s��}���SRV��Y)����DI&0T��@��� #�	�#�4!�U5!�6!�7!�8��e�F�2��Ep$VALUt��%��ֱ|��/��� ;��1�q�����(_�AN�#�ғ�Rɀ(���TOTAL��S���PW�Il��REGGEN�1�cX��`ks(��a���`TR��R��_S� ��1ଃAV�����⹂Z�E���p�q��Vr���V_�H��DA�S����S�_Y,1�R4�S� A�R�P2� ^�IG_SE	s����å�_Zp��C_�Ƃ�E�NHANC�a�/ T ;�������INT�.��@F�Psİ_OVRsP��`p�`��Lv��o���7�}��Z�@�SLG�AA�~�25�	���D��S�BĤDEb�U�����TE�P>���� !Y���
�J��$2�IL_�MC�x r#_��`TQ@�`��q���'�BV��C�P_� 0�M��	V1�
V1�2��2�3�3�4�4�
�!���� � �m�A�2IN~VIABP���1�2�U2�3�3�4��4�A@-�C2���{p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KE�EP_HNADD"!!`$^�j)C�Q��A�$��"	��#O�a�_$A�!�0�#i��#REM�"�$��½%��!�(U}�e�$HP�WD  `#S�BMSK|)G�q�U2:�P	�COLLAB� �!K5�B��h ��g��pITI1p{9p#>D� ,�@�FLAP��$SY�N �<M�`C6��~�UP_DLYAA=�ErDELA�0�ڐ�Y�`AD�Q���QSKIP=E�� ���XpOfPNTv�A�0P_Xp�rG �p�RU@,G��:I+�:I B1:IG�9JT�9Ja�9J�n�9J{�9J9<��R=A=s� X����4�%1�QB� NFL#IC�s�@J�U�H�LwNO_H�0�"?�֌RITg��@_P�A�pG�Q� ���^�U��W��LV�>d�NGRLT�0_q���O�  " ��OS��T�_JvA V	�APPR_WEIGH�s�J4CH?pvTOR8��vT��LOO��]�D+�tVJ�е�ғA�Q�U�S�XOB'�'��1SJ2P���7�X�T�<a43DP=`Ԡ\"p<a�q\!��RDC�ѮL� �рR��R�`� �RV��jr�b�RGE��*��cNFLG�a�Z���SsPC�s�UM_<`>^2TH2NH��P~.a 1� m`�EF11��� �lQ �!#� <�p3AT� g�S�&�Vr�p�t�Mq�Lr���HO�MEwr t2'r�-?Qcu�y�t3'r���P����4'r�'�@9�K�]�o����5'r뤏��ȏڏ����6'r�!�3�E�W�i�{��7'r힟��Pԟ����8'r��@-�?�Q�c�u��S$0
�q�p�� sF��`��1�"`P����0�`/���-�IO[M��I֠��*�POW=E�� ��0rZa*��� �5ވ�$DSB GN�AL���0Cp���laS2323�� Ɍ~`��� / ICEQP��PEp��5PsIT����OPBx0ޣ�FLOW�@TR`vP��!U���CU�M��UXT�A��w�ERFAC�� Uv��)�SCH��'� tQ  _��>�f�Q$����OM���A�`T�P#UP%D7 A�ct�T��U�EX@�ȟ�U EFqA: X"�1RSPT�N����T ��PPaA�0o񩩕`EXP��IOS���)ԭ�_`���%��C�WR�A���ѩD�ag֕`ԦF�RIENDsaC2U�F7P����TOOLΫ�MYH C2LE�NGTH_VTE��I��Ӆ$S�E����UFINV�_���RGI��{QITI5B��X�v��-�G2-�G1@7�w�SG�X��_��UQQD=#���AS�Äd~C�`��q����$$C/�S�`�����S0p������VERSI� ���p��5��I𼰲�����AAVM�_Y�2 �� 0  G�5��C�O�@�.r� r�	 ����S0����������������
?Q�Y�BS���1���� < -������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO`|O�O�O�OiCC�@�XLMT��C�n�  ��DIN�O��A�Dq�EXE�H4PV_��ATQz
���LARMRE?COV �R�gLMDG�p*��5�OLM_IF *��`d�O�_�_ �_�_j�_'o9oKo]onm, 
��od b��o�o�o�o^��$�� z, A   �2D{�PPINFoO u[ �V w��������` �������*�� &�`�J���n�����DQ����
��.�@� R�d�v���������a
PPLICAT��?�P��`�HandlingTool 
�� 
V8.30�P/40Cpɔ_L?I
883���ɕ$ME
F0�G�4�-

3�98�ɘ�%�z�
7DC3��ɜ
�NoneɘV�r���ɞ@�6d� Vq_ACGTIVU��C���MODP���C�I~��HGAPON���OUP�1*�� i�m��d��Қ_����1*�S  �@������ ��Q���Կ�@��
����� �3��5�Hʵl��K�HTTHKY _��/�M�SϹ����� ����%�7ߑ�[�m� ߝߣߵ��������� �!�3��W�i�{�� ������������� /���S�e�w������� ��������+� Oas����� ��'�K] o������� �/#/}/G/Y/k/�/ �/�/�/�/�/�/�/? ?y?C?U?g?�?�?�? �?�?�?�?�?	OOuO ?OQOcO�O�O�O�O�O �O�O�O__q_;_M_ __}_�_�_�_�_�_�_�kŭ�TOp��
�DO_CLEAN9�|�pcNM  !{衮o�o�o�o�o���DSPDRYRLwo��HI��m@�o r����������&�8�J���MA�XݐWdak�H�h�X�Wd�d���PLU�GGW�Xgd��PRUC)pB�`�ka�S�Oǂ2DtSEGF0�K� �+��o �or����������%�LAPOb�x�� � 2�D�V�h�z��������¯ԯ�+�TOTA�L����+�USENUO�\� e�A�k����RGDISPM+MC.���C6�z��@@Dr\�OMpo��:�X�_STRIN�G 1	(�
��M!�S�
~��_ITEM1Ƕ  n������ +�=�O�a�sυϗϩ� ����������'�9��I/O SI�GNAL��T�ryout Mo{deȵInpy��Simulate�ḏOut���OVERRLp �= 100˲I?n cycl�̱�Prog Ab�or��̱u�St�atusʳ	HeartbeatƷ�MH Faul<	��Aler�L� :�L�^�p��������� ScûSa տ��-�?�Q�c�u��� �������������);M_q��WOR.�û����� �+=Oas �������//'.PO����M  �6/p/�/�/�/�/�/ �/�/ ??$?6?H?Z?�l?~?�?�?�?�?H"DEVP.�0d/�?O*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_|\_n_PALT	� �Q�o_�_�_�_�_o o)o;oMo_oqo�o�o��o�o�o�o�o�_GRIm�û9q�_a s������� ��'�9�K�]�o�������'�R	�݁Q ����)�;�M�_�q� ��������˟ݟ����%�7�I�ˏPREG�^����[�����ͯ ߯���'�9�K�]� o���������ɿۿ�~O��$ARG_� �D ?	����0�� � 	$O�	[D�]D��O�e�#��SBN_CONF�IG 
0˃����}�CII_S�AVE  O������#�TCELL�SETUP �0�%  OME_�IOO�O�%MO�V_H������RE�P��J��UTOB�ACK����FRA:\o�� Q�o���'`r��o���� �� f�o������*�!�3�`�Ԉ�� f����������o� {��&�8�J�\�n��� ���������������� "4FXj|�������끁�  ��_i�_\A�TBCKCTL.�TMP 6.VD� GIF PHD�_q��N�t�#��f�INI�P��Օ�c�MESS�AG�����8��ODE_D����z���O�0�c�PAUS�M!!�0� (�73�U/g+(O d/�/x/�/�/�/�/�/ �/???P?>?t?1��0$: TSK  �@-��T�f�UPDT���d�0
&XW?ZD_ENB����6STA�0��5"��XIS��UNT �20Ž� � �	 ��z���en�g�-뷛G�S�o�U@��H�����zF�Oo�}Cw*�g�^���с.�O�O�O�O/_2FM[ET߀2CMPTA�A��@�$�A-�@����@���@����]5��5�(�d5��P5�r��5F*5�3�38]SCRDCF�G 1�6%�Ь�Ź�_�_�oo(o:oLo��o�Q ���_�o�o�o�o�o�o ]o�o>Pbt�`��o9�i�GR<@�M/�s/NA��/�	i��v_ED��1�Y� 
 ��%-5EDT�-�'�GETDgATAU�o�9��P?�j�H�o�f�\�x�A��  ����2�&�!�E���: IB���~�ŏ׏m����3��&۔��D���ߟJ�����9�ǟ�4 ���ϯ�(����]�o�����5N����� �(�w��)�;�ѿ_��6ϊ�gϮ�(�C�@����ϝ�+��7�� V�3�z�(��z�����i����8��&���~�]���F�ߟ�5���B�9~������]�����Y�k�����CR�!ߖ���W�q����#�5���Y��p$�NO�_DEL��rGE?_UNUSE��t�IGALLOW �1��(�*SYSTEM*�S	$SERV�_GR�V� : REG�$�\� �NUM�
��P�MUB ULA�YNP\PM�PAL�CYC10#6 $\ULSU�8:!�Lr�BOX�ORI�CUR_���PMCNV6�10L�T4DLI�0��	����BN/`/r/�/��/�/�/�/���pLA�L_OUT ��;���qWD_AB�OR=f�q;0IT_R_RTN�7�o	�;0NONS�0�6� 
HCCFS_U?TIL #<�5�CC_@6A 2#; h ?�?�?O�#O6]CE_OPT;IOc8qF@�RIA_Ic f5�Y@�2�0F�Q�=2q&}�A_LI�M�2.� ���P�]B��KXʊP
�P�2O�Q�R�B�r�qF�PQ 5T1)TR�H�_:J�F_PARAMGoP 1�<g^�&S�_�_�_�_�VC��  C�d�`��o!o`�`�`�
`�Cd��Tii:ah:e>eBa�GgC�`~� D� D	�`m�w?��2HE �ONFI� E?�aG�_P�1#; ���o1C�Ugy�aKPAU�S�1�yC ,�������� �	�C�-�g�Q�w���@������я���rO�A��O�H�LLECT_�B�IPV6��EN. QF�3�ND�E>� �G�7�1234567890��sB�TR�����%
 H�/%) �������W���0� B���f�x���㯮��� ү+�����s�>�P� b����������ο� �K��(�:ϓ�^�|�:�B!F� �I|�IO #��<U%�e6�'�9�K���T-R�P2$��(9X�t�Y޼`%�̓ڥH���_MOR�3&��=��@XB� �a��A�$��H�6� l�~���~S��'�=�r�_A?�a�a`��@K(��R�dP��)F�ha�-�_�'�9�%
�k��G� ��%yZ�%��`�@]c.�PDB��+����cpmidbag��	�`:������p��N  #��@��.���]ܭ@s<�V^��@sg�$�fl�q>��ud1:���:J��DEF *�ۈ��)�c�b?uf.txt�����_L64FIX ,������l/ [Y/�/}/�/�/�/�/ 
?�/.?@??d?v?U? �?�?�?�?�?�?,/>#__E -���<�2ODOVOhOzO�O6&I�M��.o�YU>�c��d�
�IMC��2/����dU�C�Ӌ20�M�QT:Uw�C�z  B�i�A����A���Au��gB3�*C?G�B<�=w�i��B.��B����B��5B�$�D�%B���e�zVC�q�C�v��D���D-l�E\D��n�j��B9"��22�o�D|����� ����C�C�����
�xObi�DY4cdv`D��`/�`�v`s]E�D D��` E4�F*�� Ec��FC���u[F���E���fE��fF���3FY�F��P3�Z��@�33� ;��>L��T�Aw�n,a@��@e�5Y���a���`At��w�=�`<#�*�
��?�ozJRSMOFST (��,bIT1��D @3���
д�'�a��;��bw?��ߚ<�M�NTEKST�1O�CR@��4��>VC5`A��w�Ia+a�aORI`C6TPB�U�C�`4�s��r��:d�*��qI?�5��qT�_�PROG ���
�%$/ˏ�t��N�USER  �U�������KEY_T�BL  �����#a��	
�� �!"#$%&'()*+,-./���:;<=>?@A�BC�GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~�������������������������������������������������������������������������������͓���������������������������������耇�������������������������LCK�
�����STAT/��s_�AUTO_DO ��	�c�INDTO_ENBP���Rpq�n�`�T2����ST�Or`���XC�� �26�) 8
S�ONY XC-5�6�"b����@���F( А�HR50w���>��P�7b�t�Aff����ֿ� Ŀ�� ��C�U�0�yϋ�fϯ� �Ϝ��������-ߜ��TRL��LETE�ͦ ��T_SCREEN �ڟkcs���U��MMENU 1=7�� <ܹ� ��w��������� K�"�4��X�j��� ����������5��� k�B�T�z��������� ������.g> P�t����� �Q(:�^ p����/�� ;//$/J/�/Z/l/�/ �/�/�/�/�/�/7??  ?m?D?V?�?z?�?�? �?�?�?!O�?
OWO.O @OfO�OvO�O�O(y��?REG 8�y�����`�M�ߎ�_M�ANUAL�k�DwBCO��RIGY��9�DBG_ERRML��9�ۉq�ر_�_�_ ^QNU�MLI�pϡ�pd�
�
^QPXWOR/K 1:���_5o�GoYoko}oӍDBT;B_N� ;������ADB__AWAYfS�q/GCP 
�=�p�f�_AL�pR��bbRY��[�
�WX_�P 1<{y�n�,�%oc��P��h_M��I�SO��k@L��sON�TIMX��
�ɼ�vy
��2sMO�TNEND�1tR�ECORD 1B΋� ���sG�O�]�K��{�b���� ����V�Ǐ�]���� 6�H�Z��������� #�؟������2��� V�şz��������ԯ C���g��.�@�R��� v�寚�	���п��� c�χ�#ϫ�`�rτ� ��Ϻ�)ϳ�M��� &�8ߧ�\�G�Uߒ�� ������I������4��� �p7�n���ߤ� ���������"��� F�1���|�������� [�����i���BT�f���bTOLEoRENC�dB�'r��`L��^PCSS�_CCSCB 3IC>y�`IP�t} �~�<�_`r �K�����/�{��5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O��O�O�O_�~�LL� D��&qET�c��a C[C��PZP^r_ A�J� p� �sp��Q<GPt[	 A�p�Q�_�[? �_�[oU��p�P�pSB�V�c�(a�PWoio({h+�o�X�o�o�Y��[	r�hL�W��N:p����}6ګ�c��a�D@VB��|��G���+?��K� �otGhXGr�So�����eB   =���Ͷa>�tYB�D� �pC�p�q�aA"�H�S�Q-��q���u�d�v�����AfP `; 0���D^P�֨p@�a
�QX THQ����a aW>� �a9P��b�e:��L�^�h�Hc�́PQ �RFQ�PU�z�֟�o \^��-�?��c�u�X���zCz�ů�b2�Щ�RD�����l)*����S ̡0��]�0�.��@���EQ�p��F�X�ѿ�Uҁп�VSȺNSTCY 1E�
�]�ڿ��K�]� oρϓϥϷ������� ���#�5�G�Y�k�}���ߒ��DEVIC�E 1F5�  MZ�۶a��	� ��?�6�c���	{䰟����_HNDGD �G5�VP���R�LS 2H�ݠ��/�A��S�e�w����� ZPA?RAM I�Fg�He�RBT 2-K��8р<��WPVpC�C��,`¢PQ�Z�z��%{�C��2�jMTLU,`"nPB, s� �M� }�gT�g��
#B��!�bcy� [2Dchz�����/��/gT#�I%D��C�` �b!�R��A��A�,��Bd��A5��P��_C4kP�!�2�C��$Ɓ�]�f�fA�À��B�� �| ���/�/�T (��54a5�} %/7/d?/M?_?q? �?�?�?�?�?O�?O O%O7OIO�OmOO�O �O�O�O�O�O�OJ_!_ 3_�_�_3�_�_�_�_ �_o�_(ooLo^oЁ =?k_IoS_�o�o�o�o �o�o�o#5G �k}����� ��H��1�~�U�g� y�ƏAo�Տ���2� D�/�h�S���go���� ԟ����ϟ���R� )�;���_�q������� ���ݯ�<��%�7� I�[�m��������� }�&��J�5�n�Yϒ� �Ϗ��ϣ�ѿ���� ��F��/�Aߎ�e�w� �ߛ߭���������B� �+�x�O�a���� ��������,���%�b� M���q����������� ����L#5� Yk}��� � �61CUg �������� 	//h/���/w/�/�/ �/�/�/
?�/.?@? I/[/1/_?q?�?�?�? �?�?�?�?OO%OrO IO[O�OO�O�O�O�O �O&_�O_\_3_E_W_ �_?�_�_�_�_�_"o oFo1ojoE?s_�_�o m_�o�o�o�o�o0 f=Oa��� �������b� 9�K���o���Ώ��[o ��(��L�7�I����m������$DCS�S_SLAVE �L���ё���_4D�  љ��CFoG Mѕ��������FR�A:\ĐL-�%0�4d.CSV�� � }�� ���A Vi�CHq�z����p��|�����  ������Ρޯ̩ˡҐ-矩*����_CR�C_OUT N�������_FS�I ?њ ����k�}����� ��ſ׿ �����H� C�U�gϐϋϝϯ��� ������ ��-�?�h� c�u߇߽߰߫����� ����@�;�M�_�� ������������� �%�7�`�[�m���� ������������8 3EW�{��� ���/X Sew����� ��/0/+/=/O/x/ s/�/�/�/�/�/�/? ??'?P?K?]?o?�? �?�?�?�?�?�?�?(O #O5OGOpOkO}O�O�O �O�O�O _�O__H_ C_U_g_�_�_�_�_�_ �_�_�_ oo-o?oho couo�o�o�o�o�o�o �o@;M_� �������� �%�7�`�[�m���� ����Ǐ������8� 3�E�W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿� ��'�P�K�]�oϘ� �ϥϷ���������(� #�5�G�p�k�}ߏ߸� ������ �����H� C�U�g������� ������ ��-�?�h� c�u������������� ��@;M_� ������� %7`[m� ������/8/ 3/E/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO�sO�O�O�O�O�C�$�DCS_C_FS�O ?�����A P �O�O_?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo ~o�o�o�o�o�o�o�o 72DVz� ������
�� .�W�R�d�v������� ������/�*�<� N�w�r���������̟ ޟ���&�O�J�\� n���������߯گ� ��'�"�4�F�o�j�|� ������Ŀֿ�������G�B�T��OC_RPI�N_jϳ��� �ς��O����1�Z�U��NSL��@&�h߱� ��������"��/�A� j�e�w������� ������B�=�O�a� ���������������� '9b]o� ������� :5GY�}�� ����///1/ Z/U/g/y/�/�/�/�/ �/�/�/	?2?-???Q? z?u?��ߤ߆?�?�? �?OO@O;OMO_O�O �O�O�O�O�O�O�O_ _%_7_`_[_m__�_ �_�_�_�_�_�_o8o 3oEoWo�o{o�o�o�o �o�o�o/X Sew����� ���0�+�=�O�x� s���������͏ߏ� ��'�P�K�]�o������ �PRE_CH�K P۪�A ~��,8�2x��� 	 8�9�K���+�q���a� ������ݯ�ͯ�%� �I�[�9����o��� ǿ��׿���)�3�E� �i�{�YϟϱϏ��� ��������-�S�1� c߉�g�y߿��߯��� �!�+�=���a�s�Q� ����������� ���K�]�;�����q� ������������#5 �Ak{�� ����CU 3y�i���� ��/-/G/c/u/ S/�/�/�/�/�/�/? ?�/;?M?+?q?�?a? �?�?�?�?�?�?�?%O ?/Q/[OmOO�O�O�O �O�O�O�O_�O3_E_ #_U_{_Y_�_�_�_�_ �_�_�_o/ooSoeo GO�o�o=o�o�o�o�o �o=-s� c������� '��K�]�woi���5� ��ɏ��������5� G�%�k�}�[������� ן�ǟ����C�U� o�A�����{���ӯ�� ��	��-�?��c�u� S�������Ͽ῿�� ���'�M�+�=σϕ� w�����m������%� 7��[�m�K�}ߣ߁� ���߷����!���E� W�5�{��ϱ���e� ������	�/��?�e� C�U������������� ��=O-s� ���]���� '9]oM�� �����/�5/ G/%/k/}/[/�/�/� �/�/�/�/?1??U? g?E?�?�?{?�?�?�? �?	O�?O?OOOOuO SOeO�O�O�/�O�O�O _)__M___=_�_�_ s_�_�_�_�_o�_�_ 7oIo'omoo]o�o�o �O�o�o�o!�o1 W5g�k}�� ����/�A��e� w�U�������я��o ����	�O�a�?��� ��u���͟����� '�9��]�o�M����� ����ۯ��ǯ�#�ů G�Y�7�}���m���ſ �����ٿ�1��A� g�E�wϝ�{ύ����� ��	�߽�?�Q�/�u� ��e߽߫ߛ������� �)���_�q�O�� ������������ 7�I���Y��]����� ����������!3 WiG��}�� ��%�A�1 w�g����� �/+/	/O/a/?/�/ �/u/�/�/�/�/? �/9?K?�/o?�?_?�? �?�?�?�?�?O#OO GOYO7OiO�OmO�O�O �O�O�O_�O1_C_%? g_y__�_�_�_�_�_ �_�_o�_+oQo/oAo �o�owo�o�o�o�o �o);U__q� �������%� �I�[�9����o��� Ǐ�����ۏ!�3�M ?�i��Y�������՟ �ş����A�S�1� w���g�����������ӯ�+�=��$DC�S_SGN Q�K�c��7m� �16-MAY�-19 10:1�7   O�l�4-�JANt�08:3�8}����� N.DѤ����������h�x,rWf�*σ�^M�� � O�VERSIO�N [�V�3.5.13�E�FLOGIC 1�RK��  	���P�?��P�N�!�PROG_�ENB  ���6Ù�o�ULSE � TŇ�!�_A�CCLIM�����Ö��WRS�TJNT��c��K�EMOx̘��� ����INIT S�.�G�Z���OPT_�SL ?	,��
� 	R575���Y�74^�6_�7V_�50��1��2_��@ȭ��<�TO  �Hݷ���V�DKEX��dc����PATH A[��A\�g�y��H�CP_CLNTI�D ?��6� �@ȸ����IAG_GRP 2XK�� ,`���� �9�$�]��H�����1234567890����S�� |�����p��!�� �� H���;�dC�S���6����� .�Rv�f� �H��//�</ N/�"/p/�/t/�/�/ V/h/�/?&??J?\? �/l?B?�?�?�?�?�? v?O�?4OFO$OjO|O OE��Oy��O�O_ �O2_��_T_y_d_�_:,
�B^ 4�_�_ ~_`Oo�O&oLo^oI� �Tjo�o.o�o�o�o�o  �O'�_K6H� l������� #��G�2�k�V���B] ���Ǐُ��������(��L�B\Drx��@��PC�����4  79֐�$��>���:������ߟʟܟ���CT�_CONFIG �Y��Ӛ��egU���STB_F_TTS��
�ɠb����Û�u�O�M�AU��|��MSW�_CF6�Z��  ��OCVIEWf��[ɭ����� �-�?�Q�c�u�G�	� ����¿Կ������ .�@�R�d�v�ϚϬ� ��������ߕ�*�<� N�`�r߄�ߨߺ��� ������&�8�J�\� n���!�������� �����4�F�X�j�|�,���RC£\�e��!*�B^�������C2g{�SBL_�FAULT ]���ި�GPMSK�k��*�TDIAG' ^:�աI���UD1: 6�78901234!5�G�BSP�- ?Qcu���� ���//)/;/M/.� �
@q�|�/$�TRECP��

��/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO�i/{/xO�/UMP_?OPTIONk��F�ATR¢l��	�E�PMEj��OY_T�EMP  Èϓ3B�J�P�AP�DUNI��m�Q���YN_BRK �_ɩ�EMGDI_STA"U�aQ�SUNC_S1`ɫ C�FO�_�_�^
�^dpOoo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �E�����y�Q� �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d��z��� ����˟����%� 7�I�[�m�������� ǯٯ����!�3�E� W�i���������ÿݟ �����/�A�S�e� wωϛϭϿ������� ��+�=�O�a�{�i� �ߩ߻�տ������ '�9�K�]�o���� �����������#�5� G�Y�s߅ߏ�����i� ������1CU gy������ �	-?Qk�}� ��������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?u?�?�?�? ��?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_m? w_�_�_�_�?�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9Ke_W��� �_�_����#�5� G�Y�k�}�������ŏ ׏�����1�C�] oy��������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;���g�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� _�i�{ߍߟ߹����� ������/�A�S�e� w����������� ��+�=�W�E�s��� ���ߧ������� '9K]o��� �����#5 O�a�k}�E��� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-?GYc?u? �?�?��?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_Q?[_m__�_�?�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/I_Se w��_����� ��+�=�O�a�s��� ������͏ߏ��� '�A3�]�o����� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����9�K�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� ߑ�C�M�_�q߃ߝ� �߹���������%� 7�I�[�m����� ���������!�;�E� W�i�{��ߟ������� ����/ASe w������� 3�!Oas�� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?+= G?Y?k?!?��?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	_#?5??_Q_c_u_ �?�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o-_ 7I[m�_��� �����!�3�E� W�i�{�������ÏՏ ����%/�A�S�e� q�������џ��� ��+�=�O�a�s��� ������ͯ߯��� �9�K�]�w������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� �������'�1�C�U� g߁��ߝ߯������� ��	��-�?�Q�c�u� �����������m� �)�;�M�_�y߃��� ����������% 7I[m��� �����!3E Wq�{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ �/+?=?O?i_?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O�O�O�O�O? �$�ENETMODE� 1aj5_�  00�54_F[PRRO�R_PROG �%#Z%6�_�YdUTABLE  #[�t?�_�_�_gdRSEV_NUM 2R  �-Q�)`dQ_AUTO_?ENB  PU+S�aT_NO>a b�#[EQ(b  *U��`��`��`��`�4`+�`�o�o�oZdH�IS%c1+PSk_A�LM 1c#[ e�4�l0+�o�;M_q���o_\b``  #[a�FR�zPTCP_V_ER !#Z!�_��$EXTLOGo_REQ�f�Qi�,�SIZ5�'�ST�KR�oe�)�T�OL  1Dz��b�A '�_B�WD�p��Hf��D�_�DI�� dj5�SdDT1KRņST�EPя�P��OP�_DOt�QFAC�TORY_TUN��gd<�DR_GR�P 1e#YNad �	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ�ԟ��� 1��U�@�y�d�v������ӯ����LW
 �J�kp�,��t�ۯ�j�U���y�B��  B୰���$�  A@��s�@U�UUӾ�������Eﻀ E�`F@ F�5U/�,���L���M���Jk�Lzp��JP��Fg�f��?�  s��9��Y9}�9���8j
�6��6�;���A���O ���� � I ������[�FEATURE �fj5��JQ�Handlin�gTool � �"
PEn�glish Di�ctionary��def.4�D St�ard��  
! h�Analog �I/OI�  !�
IX�gle S/hiftI�d�X��uto Soft�ware Upd�ate  rt �sѓ�matic �Backup�3�\st��gr�ound Edi�t��fd
Camera`��Fd�e��CnrROndIm���3��Common calib UI��_ Ethe�n���"�Monitor��LOAD8�tr~�Reliaby��O�ENS�Data Acquis>���m.fdp�ia�gnos��]�i�D�ocument �VieweJ��8�70p�ual �Check Saofety*� cy�� �hanced Us��Fr�����C �xt. DI�O :�fi�� m�8���end��ErrI�L��S������s  t Pa��r[�� ���J9�44FCTN_ Menu��ve��M� J9l�TP �InT�fac{� � 744��G��p� Mask Ex�c��g�� R85��T��Proxy� Sv��  15� J�igh-S�pe��Ski
� �R738Г��m�munic��on�s�S R7��uqrr�T�d�022���aю�connecwt 2� J5���Incr��str�u,Қ�2 R�KAREL Cmod. L��ua���R860hRunw-Ti��EnvL��oa��KU�el u+��s��S/W����7�Licensye���rodu� �ogBook(S�ystem)�A�D pMAC�ROs,��/Of�fs��2�NDs�M�H�� ����M�MRC�?��ORD�E� echSto�p��t? � 84�fMi$�|� 13dx��]е�׏����Modz�witc�hI�VP��?��.� sv��2Op�tm�8�2��fi�l��I ��2g �4 !+ulti�-T�����;�PCM funY�Po|���4$�b&/Regi� r �Pri��FK+7����g Num Se-lW  F�#��� Adju���6�0.��%|� fe<���&tatu�!$�6���%��  9 �J6RDM �Robot)�sc�ove2� 561N��RemU�n@�� 8 (S�F3Se�rvo�ҩ�)�SNPX b<�I�\dcs�0}��Libr1��H� �5� f�0��[58��So� tr��ssag4%G 91��p ��&0����p/I��  (�ig TMILIBx(MӋ�Firm�����gd7���s�Ac�c����0�XATX��Heln��*LR�"1��Spac��Arquz�imu�laH��� Q���Tou�Pa��I���T��c��&��ev�. f.sv?USB po��"��iP�a��  r�"1Unexcep�t��`0i$/����H[59� VC&�r��[6���P{��RcJ�PRIN�V�; d� T@�TSP C�SUI�� r�[X�C��#Web P9l6�%d -c�1R�@4d�����I�R66?0FV�L�!FV�GridK1play C�lh@���і5RiR�R.@���R-35iA���Ascii���"�η� 51f�cUp9l� � (T�����S��@rityA?voidM �`���CE��rk�C�ol%�@�GuF� 5P��j}P����
 B�zL�t� 120C C� o�І!J��P�Бy��� o=q�b �@DCS b ./��c��O��q��`�;� ���qckpaboE4�DH@�OT�~��main N��r�1.�H��an.�t�A> aB!FRLM����!i ���MI 7Dev�  (�1�G h8j��spiJP@��� �@��Ae1/�r����!hP� M-A2� i��߂^0i��p6�PC��  �iA/'�Pass�wo�qT�ROS� 4����qeda�SN��Cli�����G6x Ar�� 47��!���5s�DER\��Tsup>RtОI�7 (M�a�T2�DV�
�3D Tri-���&��_�8;�
�A�@Def�?����Ba: d7eRe p 4t0���e�+�V�st6�4MB DRAM��h86΢FR�O֫0�Arc� v#isI�ԙ�n��7|� ), �b�He�al�wJ�\h��C'ell`��p� �sh[��� Kqw�c�� - �v���pX	VCv�tyy�s�"^Ѐ6�ut� �v�m���xs ���TD_0��J�m�` �2��a[�>R ts=i�MAILYk��/F2�h��ࠛ 9�0 H��F02]�q2�P5'���T1C��5�����FC��U�F�9�GigEH�S�t8�0/A� if�!2v��boF�dri=c� �OLF�S�����" H5k�OgPT ��49f88���cro6���@��l�ApA�Sy�n.(RSS) �1L�\1y�rH�L� �(2x5�5�d�pCV�x9����est�$S�Р��> \pϐSS�F�e$�tex�D �o���A�	� BP����a�(R00�Qi#rt��:���2)�D���1�e�VKb@l �Bui, n��WACPLf��0��Va��kT�XCGM��D��L8����[CRG&a&�YBU��YKfL�p�pf��k�\sm�ZCTAf�@�О�Bf2�и��V#�s���� r���CB���
Pf���WE��!��
���T�p��DT�&4 Y�V�`���EH����
�61�Z��
�R=2�
�E 	(Np��F�V�PK�B����#��Gf1`?GD���H�р?I�e ����LD�L��N��7\s@���`����M��dela�<,��2�M�� "L[P��`?��_P�%�����S��-F��TSO�W�J5�7��VGF�|�V;P2֥ 5\b�`0�&�cV:���T;T�� �<�ce,?V{PD��$
T;YF��DI)�<I�'a\so<��a-�6J�c6s6�4L�M�V9R�h���Tri�� ���5�` �f�@��������P
� ����`��IOmg PH�[l�6�I/A  VP�S��U�Ow��!%S|�Skastdpn)���t�� SWIMEkST�BFe�00��-Q� �_�PB�_�RGued�_�T�!�_��S ��_bH573�o2c2��-oNbJ5�N�Iojb)�Cdo�cx E��o�_�lp��o�TdP �o�c�B�or�2.r�ٱ(Jsp�EfrSE�o�f1�}�r3 R�GoeELS��sL ����s�����B	�0�S\ $�F�ryz�ftl�o~�g�o����������?�����P   �n�&�"�l ��T �@<�^��Y��e�uy8Z���alib���Γ��ɟ3���埿�\v ��e\c�6�Z�qf�T�v�R VW�r��8S��UJ91��0��i�ů[c91+o�wy8���847� :��A4�j��Q��t6�<m���vrc.����0HR���ot�0ݿN��  ��8ޯf�460�>eS0L�97���U�ЄϦ�60.� g�н�+���'�ܠ�Ϻ�8co��D	M߱U"�����ߕp�i�߲T! ��n	a;�� ���u%��ⅰI��loR�d��1a59gϱŭ�&��95�ϔ�R����1��?��o�#��1A��/���vt{�UWe0ǟ���ￇ73[���97�ρ�C W���62K�=fR���8���������d����2 �ڔ����@�@y" "http������t7 �� v 3R7��78�����4�� ��TTPT��#	��ePCV�4/v߀�j�Q�Fa�7��$N�0�/2�rI�O�)/;/M/6.sv�3�64i�oS�l? torah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4c.K?�g'�)�s24g?�� (B�O�d�\iOA5sb�?U_�?vi�/i��/��/Wn��`�o%�F o�4l�$of��oXF� I)xo�cmp\�7��mp���duC`��lh����o(A�_Bt� �o]6P��m�I?0�w�@���naO��	4*O0wi�%P�?"�bsg?�]7�YE$M���8woVJ�/ե311?o��DMs�BC��7J�\���r(�52�XFa AP��ڟ<�v�`/şaqqs����/Of���1�9�VR`K���ph�քH5+��=�IN/¤SkiW�/�IF��_�%��fs�I�O�l����"<𜿚$�`�����\jԿz5bO�vr�ouς�3(�ΤH (DϮ��?sG��|� �F�Ou�������D)O��*�3P$�FӅ�@k��ϻ���럴� �P�L��ʿ��pbox��ߦebo���Sh$ �>�R.�0wT{����fx6��P��D`��3��#_I\m;YEe�OԆM�hxW��=Ete,���dct\���O$kR���d���Xm*���ro30��D�l�j9��Vx'�  FC����|@�ք f?6K�ARE0�_�~ (1Kh��.cf����WpoO�_K�up���a���H/j#- 3Eqd/�84���$qu�o��/ o2o?DVo<�7C�)�s�NJ�Ԇ�|?�3l\sy`�?�40�?Τwio��u]?�w58�?,F�a$OJ�
?Ԇ"io��!�V��u&A��P�R�ߩ5, s��v1�\  Hg552B�Q21p�0R78P5�10.R0  n�el J61�4Ҡ/WA�TUP��d8P54�5*�H8R6��9_VCAM�q97P�CRImP\1tPUI�F�C8Q28  i�ngsQy0��4P P6�3P @P PSCH~��DOCVڀD �PCSU���08Q�0=PqpVEIcOCr��� P54Pwupd�PR69aP܄��PSET�pt\!hPQ`Qt�8P7`Q�!?MASK��(P?PRXY���R�7B#POCO  /\pppb36���@PR�Q��b1Pd60Q^$cJ539.eHsb~��vLCH-`~(�OPLGqK\bPQ0]`��P(`GHCR��4`S�awund�PMCSIPR`e0aPle5=Ps�p(`DSW� �  qPb`0`�aPa��(`PRQ``Tq�RE`(Poa601P�<cPCM�PHcR0@q\j23b�V�`pE`�S`UPvisP�`E` c�`UPcPR9S	a�bJ69E`s�FRDmPsRMC�N:eH931PHcS�NBARa�rHLB��USM�qc�Pg5�2�fHTCIP0cT�MIL�e"P�`eJ� �PA�PdSTPT�X6p967PTEL��p��P�`�`
Q8P8$Q48>a"PPX�8Pc95�P`[�95qq�bUEC-`F
�PUFRmPfahQCvmP90ZQVCO�`�@PVIP%�53�7sQSUIzVSX��P�SWEBIP�SH�TTIPthrQ6�2aP�!tPG���cI�G؁�`c�PGSξeIRC%��cH7�6�P�e Q�Q|�Ror��R51P s:PL�P,t53=P8u8=P
y�C�Q6]`�b�P�I��q52]`sJ5�6E`s���PDsCLt�qPt5�\rd�q375UP cR8���u95P sR55]`,s � P8s��P�`CP�P�P�SJ77P0\o�6��cRPP�cR6�ap�`�QtaT�379P`�64�Pd387]`�d90P0c ��=P,���5�9ta�T91P� ��1P(Sܒ��Qpai�P06�=P- C�PF�T`	���!aLP PTS�p.L�CAB%�I Б�IQ` ;�H�UPPa[intPMS�Pa�иD�IP|�STY%�t7\patPTO�b8�P�PLSR76�`�5�Q��WaNN�Pa�ic�qNNE`�OsRS�`�cR681Pwint'�FCB�P"(�6x�-W`M�r���!(`OBQ`pluug�`L�aot �`GOPI-���PSP�Z�PPG�Q7�`7�3ΒPRQadv�RL��(Sp�P�S��n�@�E`��� �PTS-��q W��P�`apw�`8��P`cFVR�Plc�V3D%�l�PBV�I�SAPL�Pcy�c+PAPV1�pa�_�CCGIP - uU��L�Prog+PGCCR�`�ԁB�Pi �PԁK=�"L�PH��p��(h�<�P���h�̱�@g�Bـ
�TX�%���CTC��ptp��2��P927"0ҝPs2�Qb��;TC-�rmt;�	`�#1ΒTC9`HcC[TE�Perj�EIPp.p/�E�P�c�ЮI�use��Fـverv�F%���TG�Pp� CP��%�d -h��H-�Tra�PCT�I�p��TL� TRS���p�@נ��IP�PTh�M%�lex�sQTMQ`ver, �p�SC:���F��P�v\e�PF�IPSV�"+�H�$cj�ـtr��aCTW-���CPVsGF-��SVP2mPOv\fx���pc�bؚ�e��bVP4�fx�_m��-��SVPD�-��SVPF�P_m�o�`V� cV��t�\��LmPove4���-�sVPR�\t|�tPV�Qe5.W`V6�*u"��P}�o`�М�`��CVK��N�I�IP��CV����IP=N9�Gene���D���D�R�D����  ��f谔�pos.^��inal��n�D�DeR���`��d�P��omB���on,����R�D�R��\��T�Xf��D$b��omp��� "N��P��m����! ��=C-qf����=FXU�����g F��(��Dt II��r�D���u�� "����Cx_ui X�������f2��h	Crl02��D,r9ui�Ԣ>� it2c�0�co��e"���Խا(.)� ����� ���� IQnQ �{I[ ��_= �wo��,bD�� ��|GG�� �����{4 �e� �vʷ� ��&�� 2��Z u{z������ ��TW&q~q� 5�׷&�o�? ;0��  ��2� �y�� ���W&��� ?�3� {A��e�/> ��\�3&T���� 77߸ ��{�� ���� �ֵ��&��8� �l1��S��) ���d *�J� F's� ~��� 6:0ݙ ��,��s�{�- Q�v� ���� �,սT �ZBLx6�ۯ�6 ��6����Par ��s�>�E��j�6dsq��F  ���������Dhel�����ti-S�� �Ob��Dbcf�O���V��t OFT��P< A�_�V�ZI��D���V\�qWS��= d7tle�Ean�(b{zd��titv�JZ�z�Ez XWO� H6�6���5 �H�6H691�E4܀TofkstF� Y�682�4�`�f8�04�E91�g�`3<0oBkmon_�E��xeݱ�� qlm��W0 J�fh��B�__  ZDTfL0��f(P7�Eckl`KV� �6|��D85��ّ�m\b����xo܊k�ktq��g2`.g���yLbkLV�ts��IF�bk������Id I/�f��GR� �han�L��Vy��%���%ere�����io��� ac�- A��n�h���cuA2Cl�_�^ir��)�dg��	.�@�& G��R630���p v��p�&H�f��un���R57v�OJa�vG�`Y��owc��-ASF��O��7���SM������
af��rafLa�vl�\F c�w a���?VXpoV� �30��NT "L�FFM��=����yPh	a�G-�w�� �m2.�,�t��̹π6ԯ��sdF_�MC'V����D����fslm�is�c.  �H5522��21�&dc.pR7�8����0�708J614V�ip ATUtu�@�OL�545Ҵ�INTL�6�t8 ?(VCA����sseCRI���ȑ��UI���rt�\rL�28g��N�RE��.f,�63�!��,�SCH�d =Ek�DOCV���p���C,�<�L�0Q�i;sp��EIO��xEF,�54����9���2\sl,�SETp���lр�lt2��J7�ՌMA�SK��̀PR�XY҇��7���O[CO��J6l�3�<l�� (SVl�A��H�L�@Օ��539fRsv���#1���LCH���OPL]Gf�outl�0���D��HCR
sv�g��S@�h��CSa�!�{�50��D�l�q5!�lQ��DSW��aS����̀��OP����7��PR���L<�ұ�(Sgd���gPCM���R0 �\s��5P՝���0����n�q� AJ�1��N�q�2��PRS�a���69�� (A?uFRD�Խ���RMCN���9�3A�ɐCSN�BA�F9� HLB��� M��4���h��2A�95z�HTC�aԈ�TMIL6�j�95,��857.v,PA1�ito��oTPTXҴ JK�'TEL��piL��i XpL�80�I)��p.�!��P;�J95�ԏs "N���H�U{EC��7\cs��FR��<Q��C��5;7\{VCOa�,����IP1jH��S;UI�	CSX1�A�WEBa��HsTTa�8�R62���m`��GP%�IG� %tutKIPG�Sj�| RC1_m�e�H76��7�P�ws_+�?x�R;51�\iw�N�L��H�53!��wL�98!�h�R66��H����Ԡ���@;J56��1���N0��9�ej��L���R5`%��A|�5q�r�`,�8 5��{165!��@�"�5��H84!�29���0��PJ���n; B[�J77!ԨӃR6�5h3n���y36P��3R6��-`;о pԨ@��exeK�J87��#J90�!�stu+�~@!�۵�k90�koAp�B����@!�p�@|BA�g*�n@!��Q��#06!�@[�F�FaPb�6��́,�TS�w NC[�CAB$iiͰl1I��R7��p@q�y�CMS1�rog+QM�� �� sTY$x�CTOa�nv\+��1�(�,�6�con�~0�Ի15��JNN�%ep:��P��9ORS%tx���8A�815[�FCBaUnZQ�P!�p�p{��CMOB���"G��OL��x�O�PI�$\lr[�S�Š�T	D7�U��CP�RQR9RL���S��V�~`���K�ETS�$1��0���3\�Ԩ�FVR1�LZQ�V3D$ ���BV�a�SAPL1�CL�N[�PV��	rCC1Gaԙ��CL�3�CCRA�n "Wr!B�H�CSKQ�n\0�p��)�0CTPn�ЌQe��p.!$bCt�aT0U��pCTC�yЋRC�1�1 (�s��trsl,�r��
TX��;TCaerrm�r��MC"�s��#CT]E��nrr�REa��XPj�^��rmcH�^�a"�P�QF!$����$p "�rG,1�tTG$c8��Q�H�$SCTI�!� s��CTLqdACCK�Rp)��rLa�R82��M��YPk�.���OF��.���e��{�CN���^�1�"M�^�a�С�Q`US���!$��M�QW�$m�VGF�$R M�H��P2�� H5�� ΐq��ΐ�$(M-H[�VP�uoY���h�$)��D��hg���VPF��"MHG�̑`e!�+�V/vpcm�N��ՙ�N��$��VPRqd)��CV�x�V� "�X�,�1��($TIa�t\mh:��K��etpK��A%Y�VP%ɠ�!PN����GeneB�rip����8��extt���Y�m�"�(��HB� ��)��x��������Ȣ�res.�yA�ɠn����*���p�@M�_�N��6L���Ș�yAvL�Xr�Ȉ2��"R;�Ƚ\rax��	P�� h86���Gu+ʸ�Ͽ�Se0Lɨm�9�69�P����r�Ȩ2�ɹ1��n2��h� �0L�XR}�R�I{�e� L�x���c �Ș���N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1��/�k�@���A���ruk�ʘ L�scop��H�}�ts{������s��9��j7965��Sc��h���5 J9�{�
t�PL�J	een���t I[
x�comr��Fh�L�4 J���fo��DIF�+�6�Q����rat�i|��p��1�0�
R	8l߾�M�����PB��8� �j�mK�@X�HZ����N��oڠ��3�q��v�i���80�~�l� Sl�yQ��tpk�xb�j�.�@�R� d������,/n(�8�A8�0���
:�O8��<�Q}�CO���PT.��O (��.�Xp�|�~H���?�v� �wv��8�228�pm���722�j7�^�@ƙ���c�f�=Yvr���vcu���O�O�O�O�_#_5_7�3Y_��w3v4{_�_w�ʈ��ust_�_�cus�_�Z��oo,o>opPo�io��nge���(pLy747�jWe�lʨHM47ZKE�q {���[m�MFH�?�(wsK�8J��n���o��fh9l;��wmf���?� :�}(4	<g 9J{��II)̏މ9w��X�774kﭏ&/7ntˏ݊e+���3se�/�aw��8ͤɐ��EX \�!+: X�p��~�00��nh��,:Mo+�xO��1 �"K�O��\a��# 0��.8���{h�L?��j+�mon�:��tL�/�st�?-�w�: ���)�;��(=h��;
d Pۻ�{: 7 ��� �J0֛�re�����STD�!treLANG���81�\tqd����<���rch.��x����htwv��WWָ� R79��"Lo�51 (�I�W�h�Ո�4֧aww� �v�y �623c�h a?�cti�֘!�$X�iؠ�t �Ձn,�։����j<��"AJP@�3�p�vr{�H�6��!���- SeT� Ex3�) G�J934��{LoW�4 (S������� <���91 ��8!4�j9�所+�d��y�
��	�btN�ite{�R ��I@ Ո�����P��������	 ����Z�vol ��X ��9�<�I�p����ld*���F�86!4{��?��K�	��k扐�֘1�wmsk��M�q�Xa�Ae����p���0RBT�1ks.?OPTN�qf��U$ RTCam T��y��U��y�� U��UlU6L�T@�1Tx����SFq��Ue�6T��USP; W�b DT�qT2h�T�!/&+��8TX�U\j6&��U U�Usfd�O&�&ȁT���662DPN�abi��%�Q�%62V� �$���%�� �#(�(6{To6e St�%���#5y�$�)5(To�%tT0�%5�W6�T���%�#�#orc���#I���#���%c�ct�6ؑ?�4\W6965"p6}"�#\j536���4�"��?kruO O,Im ?Np�C �?t�0<O�;�e �%���?�
;gcJ7 "AV<�?�;avsf�O__&_8WtpD_V_0GT�F|_:UcK6�_�_9r�O�3e\s�O2^�y`O:�migxGvNgW! m�%��!�%T�$E A{6�po6̀�#37N�)5R5�_2E���$0���$Ada�Vd���V�?;Tpz7�_�e7DDTF9���#8�`�%��4~y�ted Z@0�A}�@�}�04N�}�0}���}�dc& }����u 6�v��v1�u1\b�u$2}�<��}� R83�u�"x}��"}�valg���Nrh�&�8�J��Y�o�ue��� j7q0�v=1��MIG�uerfa��{q����E�N�ء��EYE�ce A���� �pV�e�A!���2Յ�Q �%��u1�e�i�@��@H�e����J0� '��b��T��E In��B�  W�|��5�37g����(MI�t�Ԇr��ݟ�Cam���nеv!g�U -�v J߆8⹖0F���P�y�ac���28���Rɏ jo��2�� djd�8r}�� og\k�0��gܕ�wmf�Fro/� Eq'�4"}��3 J8��oni[��ᅩ}Ĵ��C o� ��ʛ��m@�R�e��{n�Д�V��o������  �����裆"P�OS\����ͯ mcenϖ�⑥OMo��43��� �(Coc� An[�t���"Fe�a\�vp��.��ocflx$�le��`8�hr�tr�NT�w CF+�x E/�at	qi�M�ӓxc�֌p�f�lx����Z�c�x��
0 h��h8f��mo��=� H����)� (�vSER�,���g�0߆0\�r�vX�= ��I � - �ti��H���VC�828�5ص�L"�RC��n �G/���w�P�y�\v�vm "o�lϚ��x`��=e�ߠ-�R-3?������vM [��AX/2�)�S�r�xl�v#�0��h8�߷=� RAX�AТ����9�H�E/�Rצ����h߶"R�Xk��F�˦85ή�2L/�xB88�5_�q�Ro�0iA��5\rO�9�K��v����8���.�gn "�v��88��8s�i ?�9 �����/�$�y O�MS"����&�9R H784&�`�745�	pp��p��ycr0C�Rc�hP0� j�-�a�%?o��6D950R7tsrl��ctlO��APC���j�ui�"�L���  ����K^棆!�A��qH���&-^7����� ��616C�q�794h����� M�ƔI��99���(��$F�EAT_ADD �?	���Q~%P  	�H ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n���������TDEMO �fY   WM_��� �����//%/ R/I/[/�//�/�/�/ �/�/�/�/?!?N?E? W?�?{?�?�?�?�?�? �?�?OOJOAOSO�O wO�O�O�O�O�O�O�O __F_=_O_|_s_�_ �_�_�_�_�_�_oo Bo9oKoxooo�o�o�o �o�o�o�o>5 Gtk}���� ����:�1�C�p� g�y�������܏ӏ� ��	�6�-�?�l�c�u� ������؟ϟ���� 2�)�;�h�_�q����� ��ԯ˯ݯ���.�%� 7�d�[�m�������п ǿٿ���*�!�3�`� W�iϖύϟ������� ����&��/�\�S�e� �߉ߛ��߿������� "��+�X�O�a��� ������������� '�T�K�]��������� ��������#P GY�}���� ��LCU �y������ /	//H/?/Q/~/u/ �/�/�/�/�/�/?? ?D?;?M?z?q?�?�? �?�?�?�?
OOO@O 7OIOvOmOO�O�O�O �O�O_�O_<_3_E_ r_i_{_�_�_�_�_�_ o�_o8o/oAonoeo wo�o�o�o�o�o�o�o 4+=jas� �������0� '�9�f�]�o������� ��ɏ�����,�#�5� b�Y�k���������ş ����(��1�^�U� g������������� ��$��-�Z�Q�c��� ����������� � �)�V�M�_όσϕ� �Ϲ���������%� R�I�[߈�ߑ߫ߵ� ��������!�N�E� W��{�������� �����J�A�S��� w������������� F=O|s� ����� B9Kxo��� ���/�/>/5/ G/t/k/}/�/�/�/�/ �/?�/?:?1?C?p? g?y?�?�?�?�?�? O �?	O6O-O?OlOcOuO �O�O�O�O�O�O�O_ 2_)_;_h___q_�_�_ �_�_�_�_�_o.o%o 7odo[omo�o�o�o�o �o�o�o�o*!3` Wi������ ��&��/�\�S�e� ������������� "��+�X�O�a�{��� �������ߟ��� '�T�K�]�w������� ���ۯ���#�P� G�Y�s�}�������� ׿����L�C�U� o�yϦϝϯ������� �	��H�?�Q�k�u� �ߙ߫��������� �D�;�M�g�q��� ��������
���@� 7�I�c�m��������� ������<3E _i������ �8/A[e �������� /4/+/=/W/a/�/�/ �/�/�/�/�/�/?0? '?9?S?]?�?�?�?�? �?�?�?�?�?,O#O5O OOYO�O}O�O�O�O�O �O�O�O(__1_K_U_ �_y_�_�_�_�_�_�_ �_$oo-oGoQo~ouo �o�o�o�o�o�o�o  )CMzq�� �������%� ?�I�v�m����������ُ���;�  2�Q�c�u��� ������ϟ���� )�;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����� ��1CUg y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����'>9  :> Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{��������/=C6Yk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A���$FEAT_D�EMOIN  VE��q��>�Y�_INDEXf�u���Y�ILECOM�P g������t�T���S�ETUP2 h������  �N ܑ��_AP2�BCK 1i��  �)B���%�C�>���1�n� E����)���M�˯�� �����<�N�ݯr�� ����7�̿[��ϑ� &ϵ�J�ٿWπ�Ϥ� 3�����i��ύ�"�4� ��X���|ߎ�߲�A� ��e�����0��T� f��ߊ�����O��� s�����>���b��� o���'���K������� ��:L��p��� �5�Y�}�$ �H�l~�1 ��g�� /2/� V/�z/	/�/�/?/�/ c/�/
?�/.?�/R?d? �/�??�?�?M?�?q?@O�?O<O���P�� 2�*.V1RCO�O�0*�O�O`�3�O�O�5w@PC�O|_�0FR6:�O"=^�Oa_�KT���_ �_&U�_�\h�R_�_�6�*.FzOo�1	�(SoEl�_io�[STM �b�o�^+P�o��m�0iPen�dant Panel�o�[H�o �g��oYor�ZGIF |��e�Oa��ZJPG �*��e���z��JJS�����0�@���X�%
Ja�vaScriptُ�CSʏ1��f��ۏ %Casc�ading St�yle Shee�ts]��0
ARGNAME.DT��
�<�`\��^���Д�៍�АDISP*ן���`$�d��V��e��CLLB.cZI��=�/`:\���\�����Col�labo鯕�	P�ANEL1[�C�%��`,�l��o�o�2 a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V���zό��!ߘ�TPEINS�.XML(�@�:\�<����Custo�m Toolba�r}��PASSW�ORD���>FR�S:\��� %�Password Config� �?J���C��"O��3� ����i����"�4��� X���|�����A��� e�����0��Tf �����O�s ��>�b�[ �'�K���/ �:/L/�p/��/#/ 5/�/Y/�/}/�/$?�/ H?�/l?~??�?1?�? �?g?�?�? O�?�?VO �?zO	OsO�O?O�OcO �O
_�O._�OR_d_�O �__�_;_M_�_q_o �_�_<o�_`o�_�o�o %o�oIo�o�oo�o 8�o�on�o�!� �W�{�"��F� �j�|����/�ďS� e���������T�� x������=�ҟa��� ���,���P�ߟ񟆯 ���9����o���� (�:�ɯ^�����#� ��G�ܿk�}�ϡ�6� ſ/�l�����ϴ��� U���y�� ߯�D��� h���	ߞ�-���Q߻���߇��,��$FI�LE_DGBCK� 1i������ (� �)
SUMM?ARY.DG,���OMD:`�����Diag Su�mmary���
CONSLOG���y����$���Co�nsole lo�g%���	TPACCN��%g������TP Acco�untinF����FR6:IPKD?MP.ZIP�����
��)����Exc?eption-�����MEMCHEC�K�����8�M�emory Da�ta��LN�=)�RIPE����0�%� �Packet L�E���$Sn�S�TAT*#�� %LSta�tus�i	FTAP�/�/�:��mment TB�D=/� >)ETHERNE��/o�/�/��Et�hernU<�fi�guraL��'!DCSVRF1//)/�B?�0 verify allE?��M(5DIFF:? ?2?�?F\8diff�?}7o0CHGD1�?�?�?�LO �?sO~3&��
I2BO)O;O�O� bO�O�OGD3p�O�O�OT_ �O�{_
VUPDAT�ES.�P�_��FORS:\�_�]���Updates �List�_��PS�RBWLD.CM�o���Ro�_9�P�S_ROBOWEyL^/�/:GIG��o>_�o�Gig�E ��nosti�cW�N�>�)}�aHADOW�o�o�ob�Sha�dow Chan�ge��8+"rNOTI?=O���Notif�ic�"��O�A=�PMIO�o���h��f/��o�^U�*�UI3�E�W��&{�UI������B� ��f��_�������O� ��������>�P�ߟ t������9�ί]�� ���(���L�ۯp��� ���5�ʿܿk� Ϗ� $�6�ſZ��~��w� ��C���g���ߝ�2� ��V�h��ό�߰��� Q���u�
���@��� d��߈��)��M��� ������<�N���r� ���%�����[���� &��J��n� �3��i��" �X�|�� A�e�/�0/� T/f/��//�/=/�/��/�$�$FILE�_�PPR�P���� �����(MDONLY� 1i5�  
 �z/Q?�/u?�/ �?�?t/�?^?�?O�? )O�?MO_O�?�OO�O �OHO�OlO_�O_7_ �O[_�O_�_ _�_D_ �_�_z_o�_3oEo�_ io�_�oo�o�oRo�o vo�oA�oew �*��`�����&�O��*VIS�BCK,81;3*�.VDV����F�R:\o�ION\�DATA\��/���Vision� VD file ̏��&�<�J�4�n� �����3�ȟW���� ��"���F�՟�|�� ����m�֯e������ 0���T��x������ =�ҿa�s�ϗ�,�>� ��b���ϗϼ�K� ��o��ߥ�:���^�����ϔ��*MR2_�GRP 1j;��C4  B�}�	 71�������E�� E�  �F@ F�5U�������L����M��Jk��Lzp�JP���Fg�f�?� � S����9�Y�9}�9���8j
�6���6�;��A� � ���BH��B���B���$�������������@UUU#�����Y�D�}� h����������������
C��_CFG� k;T �M���]�NO {:
F0�� � \�RM_CHKTYP  0��}�000��O=M_MIN	x�g��50X� �SSBdl5:0��bx�Y����%TP_DEF'_OW0x�9��IRCOM���$GENOVRD�_DO*62�T[HR* d%d�o_ENB� �/RAVC��mK�� ��՚�/3�/���/�/�� ��M!OUW s���}��ؾ��8��g�;?�/7?Y?[? 7 C��0����(7l�?�<B�?B�����2��*9�N SMT�T#t[)��X�4�$�HOSTCd1u�x���?�� kMCx��;zO�x�  27.0z�@1�O  e�O �O	__-_;Z�O^_p_��_�_�LN_HS	anonymous�_ �_�_oo1o yO��FhFk�O�_�o�O�o �o�o�oJ_'9K ]�o�_���� �4o�XojoG�~�o ^�������ŏ��� ��1�T���y��� ��������,�>�@� -�t�Q�c�u������� ��ϯ���(�^�� M�_�q�����ܟ� � ݿ��H�%�7�I�[� ��ϑϣϵ����l� 2��!�3�E�Wߞ��� ¿Կ����
������ �/�v�S�e�w��� �����������+� r߄ߖ�s�����߻� ���������'9K ]�������� �4�F�X�j�l>�� }������ //1/T��y/�/��/�/�/.D\AENT� 1v
; P!\J/?  ��/ 3?"?W??{?>?�?b? �?�?�?�?�?O�?AO OeO(O�OLO^O�O�O �O�O_�O+_�O _a_ $_�_H_�_l_�_�_�_ o�_'o�_Koooo2o {oVo�o�o�o�o�o �o5�oY.�R�v��zQUICC0���3��tA14��"����t2���`�r�ӏ!ROU�TERԏ��#�!?PCJOG$����!192.168.0.10�~�sCAMPRTt�P�!d�1m������RT폟�����$N�AME !�*!�ROBO���S_CFG 1u�)� �A�uto-star�tedFTP&��=?/֯s�� ��0�B��f�x��� ������S������ ,���������ϼ�ޯ ���������ʿ'�9� K�]�oߒ�ߥ߷����������SM %y�{�U�ό��� �������
��.�@� c���v������������z�%�7�I�K�8 �\n���k�� ���3�FX j|����a��7/M*/</ N/`/r/9�/�/�/�/ ��/�/?&?8?J?\? �m?���?�//�? �?O"O4O�/XOjO|O �O�O�?EO�O�O�O_ _0_w?�?�?�?�O�_ �?�_�_�_�_o�O,o >oPoboto�_o�o�o �o�o�oK_]_o_L �o�_�o�����o � ��$�6�Y�Y��~�������ƏZ�_ERR w3�я��PDUSIZ  �g�^�p���>~�WRD ?r��Cq�  guestb�Q�c��u�������`�SCD�MNGRP 2x�r�����H�g�\�b�K� 	�P01.00 �8`�   �� �   B�  ��� ���H���L���L��L������O8�����l�����Ua4�  �Ȥ� ��8���\���)j�`�;�������d�.�@�R�ɛ__GROUېy�����	ӑ���QUPD  ?u�����İTYg�����TTP_A�UTH 1z��� <!iPen'dan��-�l����!KAREL�:*-�6�H�KC�]�m��U�VISION SET���ϴ�!�����R� 0��H�Bߏ�f�x�����߮���CTRL C{����g�
���FFF9E3���AtFRS:D�EFAULT;��FANUC W�eb Server;�)����9�K��܀����������߄W�R_CONFIGw |ߛ ;���IDL_CPU�_PCZ�g�B��I�y� BH_�MI�Nj�)�}�GNR_�IO��g���a�N�PT_SIM_D�_�����STAL�_SCRN�� ����TPMODNT�OL������RTY`��y���� �ENO����Ѳ]�OLNK 1}��M���������eMA�STE��ɾeSL?AVE ~��c>�O_CFGٱ�BUO�O@CY�CLEn>T�_A�SG 1ߗ+�
 ����// +/=/O/a/s/�/�/�/��/��NUM�z�
@IPCH��^RTRY_CN Z���@��������� @kI��+E�z?E�a�P_M�EMBERS 2Y�ߙ� $���2����ݰ7�?�9a�S�DT_ISOLC�  ����$J_23_DSM+��3JOBPROC�N��JOG��1��+�d8G�?��+�O�/?
�LQ�O__/_�O S_e_w_�_`�O H�m@��E#?&BPOS�REQO��KANJ�I_���a[�MON ����b�yN_goyo�o�o�o�$Y�`3�<� ��e�_ִ��_L���"?`�EYLOGGIN�LE��������$LANGUAGgE ��<T�Y {q�LGa2�	��b���g�xP�� � ��g�'Զ�b���>�M�C:\RSCH\�00\<�XpN_D?ISP �+G�pH��O�O߃LOC�p�Dz���AsO�GBOOK �������󑧱����X�����Ϗ���`�a�*��	p� ����!�m��!���=p�_BUFF 1�p��2F幟����՟D� Col�laborativǖ���F�=�O�a� s�������֯ͯ߯����B�9�K���DC�S �z� =���'�f��?ɿۿ����H@{�IO 1��� ~?9Ø�� 9�I�[�mρϑϣϵ� ���������!�3�E� Y�i�{ߍߡ߱����ߴ���E��TMNd �_B�T�f�x���� ����������,�>� P�b�t�������L��SEVD0��TYPN1�$6���QRS"0&��<2�FL 1�"�J0���������GTP:pO>F�NGNAM1D��mr�tUPS�GI�"5�aO5�_LO{ADN@G %��%TI�pZUZ�AUN#�(MAXUALRM�'���(���_PR"4F0�d��1�B_PNP�� V 2�C	�MDR0771�ߕ�BL"806=3%�@ �_#?�hߒ|/�C��z��6��/���/Po@P �2��+ �ɖ	�T 	t  ��/�%W?B?{?� k?�?g?�?�?�?O�? *OONO`OCO�OoO�O �O�O�O�O_�O&_8_ _\_G_�_�_u_�_�_ �_�_�_o�_4ooXo joMo�oyo�o�o�o�o �o�o0B%fQ �u������ ��>�)�b�M����� {��������Տ�� :�%�^�p�S��������D_LDXDI�SApB�MEM�O_APjE ?=C
 �,� (�:�L�^�p�������� 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%A �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A�z�4��~�K��������K:z�j]�Q_D��^��PL_NAME �!3%,�!�Default �Personal�ity (fro�m FD) �R�R2� 1�L?6(L?�,0	l d���� ����//(/:/ L/^/p/�/�/�/�/�/�/�/ZX2u?0?B? T?f?x?�?�?�?�?\R<?�?�?O O2ODO�VOhOzO�O�O�OZZK`\R�?�N
�O_\TP�O:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHo_)_~o�o �o�o�o�o�o�o  2DVhz�[omo ����
��.�@� R�d�v���������Џ�� Ef  Fb� F7���   ��!��d��@�R�6�t��� ���l���ʝ����� ݘ���� "�@�F�d���� "�|��ݐA�  ϩ�U[�$n�B��E ��� � @D�  &�?�� �?�@��A@�;f��FH�� ;�	l,�	 '|��j�s�d�/>��� ��� �K(��Kd$2�K ��J7w��KYJ˷�ϜJ�	�ܿ�� @�I���_f�@w�z��f򿿾γ�N�������	Xl�����_��S�ĽÔ�}�I ����5�?��  ����A�?oi#�;����� ���l� �Ϫ�-���ܛ�G�G�Ѳ��@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=�����в@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj��a�Be�Ci��#��Bи�ee^��^^ȹBР ��P����̠�����ADz՟�n�3��C��i�@�R�R�Y���� { �@� ����  ���?�ff0������n� ɠ #ѱy9G
(���I�	(�@uP~����t��t���>����;�C�d;��.<���<�g�<F+<L�������,��d�,�̠?fff�?��?&&��@���@x��@��N�@���@T�H�ِ�!-�ȹ �|��
`���� ���//</'/`/`r/]/�/��eF�� �/�/�/�/m?��/tJ?�(E��G�#�� FY�T?�?P? �?�?�?�?�?O�?/O O?OeOk��O�IQO G�?�O1?�OmO_0_�B_T_������A _�_	_�_�_�_ o���A��An0 bФ/o �C�_Uo�_�Op���؃o�o�o�o���W������oC�E�� q�H�d�����a@q��e�F�Bµ�WB]�NB2��(A��@�u�\?�D��������b�0�|�u�R����
x~��ؽ��B�u*C��$�)�`�$ ����GC#����rAU�����1�eG�D�I��mH�� I:��I�6[F�﫹C�I���J�:\IT��H
~QF�y���p�*J��/ I8Y�I��KFjʻCe �o��s�����Џ��� ߏ�*��N�9�r�]� �����������۟� ��8�#�\�G�����}� ����گů���"�� �X�C�|�g�����Ŀ �������	�B�-� f�Qϊ�uχ��ϫ��� �����,��P�b�M� ��qߪߕ��߹����� ��(��L�7�p�[��@�������s($�ϳ�3:����$���3���d�,��4��@�R�wa�ǲ��l�~�wa����e����wa4 �{������(L�:ueP�P~�A �O������	����G2 W}h����� �/���O�O7/m/[(d=�s/U/�/�/�/ �/�/?�/1??U?C?�y?�=  2 E�f9gFb��77�b9fB)aa)`C9A`	�&`w`@-o�?w`e�@O)O�?MO�Ow`�?@�?�O�O�O�O9c?�0T�A7ht4w`w`�!w`xn
  �O9_K_]_o_�_�_�_ �_�_�_�_�_o#ozz�Q ��h��G����$MR_CA�BLE 2�hO �a�T� @@�0�Ae��a�a��a��`��0�`C��`�aO8�tB�^n�d��`�aE�4�E�#��o�f�#��0�|�0�DO��By`���Š��bED4E�c,��o�g8  ���Cu�07�d4
v�ے�0 �b���XE�Z&�lȠ`y`
qC�p�bHE݈
v#g�5DͣҮ�qz�lҠ`�p�0�q�p�b0�
v׸%c���b=%	E;h��u/o�c -��4tH�\�?�9�K� ]�o�ԏϏ��
�ɏۏ�@���?��eo �a���������b����� �����`�	 ����@������% �*�}0�6 ��ݐ�����`���	����@������*,� ,�-�\c�OM �ii���3� � ���%% 23�45678901�i�{� f��������ԋ��1����
���`�not �sent3������;�TEST�FECSALGRG  e�qiG�1d.�Zš
:�� �D�CbS�Q�c�u��� 9�UD1:\ma�intenanc?es.xml��ֿ�q� =���DEFAULT�-�i4\bGRP 2�M�  =��a��{p  �%�Force�s�or checkS  ���b�z��p����h5-[ �ϻ�������ϖ�D�%!1s�t cleani�ng of co�nt. v�ilation��}�R��+��[�ߔߦ߸�z��mech�gcal`�����!�0��h5k�@��R�d�v�����(�rolle_Ƶ����/���(�:�����Basic q�uarterly�������,������0����M��M��:C@"GpP�a�b`i4�������#AC���M"��{�Pbt���S�uppq�greaCse���?@/&/8/J/\/��C+ �ge��. batBn�y`/��/h5	/ �/�/�/? ?_�ѷen'�v��/�/��/��?�?�?�?�?ѣG=?O�qp"CrB1O��0�/`OrO�O��O�O�t$��Lf�B�C-m��A�O:�OO@$_6_H_Z_l_�t*�cabl�Om���B�S<m��Q�_:�
_ �_�_oo0oo)(Ӂ/�_�_���_�o�o�o��o�o�O@ha�u1�l�2r xm�<qC:��op������ReplaW�fUȼ2�:�._4�F�X�j�|�m�$%���o�������#� ��
��.�@���d��� ŏ׏����П���� U�*�y�����r����� ����	�q��?�߯c� 8�J�\�n���ϯ���� �ڿ)����"�4�F� ��jϹ�˿������� �����[�0�ϑ�f� �ϊߜ߮�����!��� E�W�,�{�P�b�t�� ���߼�����A�� (�:�L�^�������� ������� $s� H������q��� ��9]o�V hz���U�# �G/./@/R/d/� �/�/��//�/�/? ?*?y/N?�/�/�?�/ �?�?�?�?�???Oc? u?JO�?nO�O�O�O�O+J�r	 H�O�O_ _6M2_@OBE:_p_>_ P_�_�_�_�_�_ o�_ �_oHoo(oZo�o^o po�o�o�o�o�o �o� :z �bA?�w  @�q _ ���Fw�� ��H* �**  @q>v�p2T�f�x�:�p������ҏ��eO ^C7�Տ#�5�G�	�k� }���ُ���c���� �W��C�U�g���ß )�����ӯ���	�� -�w�����9��������m�Ͽ��=�O�E�	A�$MR_HI_ST 2�>uN��� 
 \�$Force� sensor �check  1�23456789�0q�3����ß��N}SB�� -319.8 �hours RU�N 9.�Y�!1�st clean�ing of c�ont. ven�tilation�0ÄϖϨ�-�Y�޹�mech��ca�li�%Ό4��o��DN�t��95���1����rol�leh�+�=�O���Y�Basic �quarterlyߒߤ߶�
O4�F� �(�����b�t� ����������M�_� ���:�����p���:��SKCFMAP � >uQ���r5�������ONREL  .��3���EXC'FEN��:
���QFNCXJJO�GOVLIM8d�Ná ��KEY8z��_PAN7�����������SFSPDTYqPxC��SIG�|:��T1MOT��G��_CE_G�RP 1�>u\�D����� /Ⱥ��/�/U/ /y/0/n/�/f/�/�/ �/	?�/???�/c?? \?�?P?�?�?�?�?�?�O)OOMO,���QZ_EDIT5 )�TCOM_CFG 1���[�O�O��O 
�ASI 	�y3�
__+[!_O_��>O�_~bHT_ARC_U�քT_MN_oMODE5�	UAP_CPL�_�gNOCHECK� ?�� �� o.o@oRodovo �o�o�o�o�o�o�o�*!NO_WA�IT_L4~GiN�T�A���EUwTo_ERRs2���3��ƱJ������>_)��|MO�s��}x:Ov���8�?����� l���rPARAM�r�����j���x5�5�G� =  r� b�t�s�X�������������֟�0�����b�t�����SUM_RSPACE������Aѯۤ�$OD�RDSP�S7cO�FFSET_CAqRt@�_�DIS���PEN_FIL�E:�7�AF�PT?ION_IO���q�M_PRG %��%$*����M�WORK �y=f ��춍�D��������	 ������gT���RG_DSBOL  ��C�{�u��RIENTT5O7 ��C� �A �UT_SIM_Dy����V�LCT ���}{B �٭��_PEqX�P=��RAT�W� dc��UP� ���`���`e�w�]ߛߩ��$��2r�L6(L�?���	l d������&�8�J� \�n��������� �����"�4�F�X���2�߈����������� ��*�<w�T fx������p�J`��ˣG���Tz�P g������/ "/4/F/X/j/|/�/�/ �/���/�/??0? B?T?f?x?�?�?�?�? �?�?�?�/�/,O>OPO bOtO�O�O�O�O�O�O �O__(_:_��O�C�y_�]2ӆ��_ �^�_�_�W^]^]��/ooSog�Hgroho zo�o�o�o�o�oF`��#|`�A�  �9y����OK�1�k�����}<�EA��nq @D� � �q����nq?��Cᾄs�q1� ;��	l��	 |��Q�s�r�q>��u �sF`H<z�H~�H3k�7GL�zHpG�99l7�k_�B�T�F`C4��k�HJ���t��-�Ae��}�k�����s�?��  �ሏ�����EeBVT����dZ�������ڏ ���q-�PFk�y�{FbU����n@6�  ���z�Fo��Be	'� � ���I� �  ��:p܋=���8ڟ웆�@�� �B�,���B���g�rAgN����  '|�X��g��B��p��BӀC׏����@ � #�Bu�&��ee�^^މB:p2���>�m�6p�Z���Dz?o}�܏ ������׿������Ǒ���� f�  � ��M���*�?��ff�_8�J�ܿ 3pϑ�ñ8�Чϵ�H�q.·�(����P�� �'��s�tL�>��/��;�Cd;��.�<߈<�g�?<F+<L ���^oiΚrd@��r6p?offf?�?&�����@��@x���@�N�@���@T싶�Z�� �ћtމ�u�߈w	�x� �ti�>�)�b�M��q� ������������� :�%�^�������W����S�E�  G�>aF�� Fk��� ������1U@y d������q� �	��{�A��h� ����a��ird��A{/w/J/5/n/vA��A���":t�/ C^/�/Z/ ލ?���/�/1??����W����g��pE� ~1�?04q�0
1�1@IӀ���BµWB]��NB2�(A����@�u\?����������b�0��|�uR�����
�>�ؽ���Bu*C���$�)`�? ����GC#����rAU�����1�eG����I�mH��� I:�I��6[F���C�4OI��J�:�\IT�H
~�QF�y�Ol@���*J�/ I8�Y�I��KFjʻC��-?�O�O_ _>_)_b_M_�_�_�_ �_�_�_�_o�_(oo %o^oIo�omo�o�o�o �o�o �o$H3 lW�{���� ���2��V�h�S� ��w�����ԏ����� ��.��R�=�v�a��� ����П����ߟ�� <�'�`�K�]������� ��ޯɯ��&�8�#��\��3(J���3:�a������J�3��c4�������x�����1����ڿ<��1���e���14 �{2�2�r�@`ϖτϺϨ��%PR�	P���!�h�!��K�6�o�Z����� u�|ߵߠ�������� ��3��W�B�{�f�4� ��������d�A�� ��!��1�3�E�{�i��������������  �2 Ef�7Fb-�7��6B�!�!�� C9� �� �0@ �/`r������#x��+=��3?, V�8v�R�0�0��0�.
 D���� �//%/7/I/[/m/p/�/�:� ��ֻ��G���$PA�RAM_MENU� ?2���  DEFPULSE�+�	WAITTM�OUT�+RCV�? SHEL�L_WRK.$CUR_STYL� ;4<OPTJJ?�PTB_?Y2C/?R?_DECSN 0�� �<�?�?�?�?�?OO ?O:OLO^O�O�O�O�O��O�!SSREL_�ID  .������EUSE_PRO/G %�*%�O0_�CCCR0�B���#�CW_HOST �!�*!HT�_=ZT ��O_�Sh_zQ�S�_><[_TIME
2�F�XU� GDEBU�G�@�+�CGINP?_FLMSKo5isTRDo5gPGAb`e %l�tkCHCo^4hTYPE�,� �O�O�o#0B kfx����� ����C�>�P�b� ��������ӏΏ��� ��(�:�c�^�p������7eWORD ?�	�+
 	RySc`��PNS�ՙC4�JOv1���TE�P�COLЀէ�2��gLP �3�����OjTRA�CECTL 1�v2��! ��/� �Қ��q�DT Q�2��Ǡ��D � �:����Ԡ�Ԡ��}��ׯ���;� 4��4��4���;�u�:�q:���;�8�	�8�
8�8�8��8�8�8��@:�
8�8���� �T��ٱ޴��� ؿ�$�6���
�l�~� @�R�dϞϰ������� ��
��V�h�zߌߞ� ����������
�,�>�@P�*�<�v��*�����˶; +8�+ (��)��*���� ��%�7�I�[�m�� �������������� !��5�G�Y�k�}��� ����ſ��С� *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6@u bt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� ��V�߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�?��?�?�1�$PGT�RACELEN � �1  ����0��6_�UP ���e�A@�1@��1_CFG ��E�3�1
@�
<D�0<DZO<C�0�uO$BDEFSPD� �/L�1�0���0H_CONF�IG �E�3� �0�0d�D�&�2 �1�APpDsAl�A�0��0IN'@?TRL �/MOA�8pEQPE�E��G�A<D�AIWLID(C�/M	bT�GRP 1ýI� l�1B � �����1A��33FC� F8� E�� @eN	�A�AsA�Y�Y�A�@?� 	 vO�Fg�_ ´8cokB;`baBo,o>oxobo��o�1>о�?B�/�o�o~�o =%<��
 C@yd��"�������  Dz@�I�@A0�q� � ������ˏ���ڏ� ��7�"�4�m�X���|����Ú)ґ
V7�.10beta1�HF @�����Aq��Q�  �?� �B���P�p �C��~&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@p���f������ҡr�R�ܣ�Rљ����1�i�������t<B!CeQKNO?W_M  lE7F�bTSV ĽJ�BoC_�b�t��������������1�]aSM��SŽK ���	�NB�0����ĿK���-�bb��A�RP���`�0�Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1=�K
 4MU�iǨj� K�]�oߠ� �ߥ߷�������2�� #�h�G�Y��}������
������,�2r7�I��1�<t�H��P3^�p�����,�A4��������,�5(:,�6Wi{�,�7����,��8�!3,�MA�D�6 F,�OV_LD  KD��xO.�PARNUM�  �MC/%�S+CH� E
9'!8G)�3Y%UPD/���E�/P�_CMP_0��0@�0'7E�$�ER_CHK�%05H�&�/�+RS����bQ_MO�+?=5_�'?O�_RES_G6��:�I�o�?�?�? �?O�?O7O*O[ONO OrO�O�O�{4]��<�?�Oz5���O__ |3 #_B_G_|3V b_ �_�_|3� �_�_�_|3 � �_�_o|3Oo>o<Co|2V 1�:�k1�!�@c?�=2T?HR_INRc0i!�}�o5d�fMASS6�o Z�gMN�o�c�MON_QUEUE �:�"�j0��UO�N� U1Nv�+DpENDFqd?`y�EXEo`u� BE�npPAsOPTIO�Mwm;DpPROGR�AM %$z%�Cp}o(/BrTASK�_I��~OCFG� �$��K�D�ATA��T���j12/ď֏��� ���+�=�O�a�����������͟��INFO�͘��3t��!� 3�E�W�i�{������� ïկ�����/�A�@S�e�w�����Θ�a '��FJ�a K_N���T��˶ENB�g ڽw1��2��G�N�2�ڻ P(O�=���]�ϸ�@���v� ��u�uɡdƷ_E?DIT �T���|��G�WERFL�x��c)�RGADJ {Ҷ�A�  $Ձ?j00��a�Dqձ���5�?�$�ʨ�<u�)%e��0����FӨ�2�R��+	H;pl�G�b_�u>�pAod�t$��*�/� **:�j0�$�@�5AY�T���^��q�� �b~�L��\�n��� ������������� 4�F�t�j�|������� ������bLB T�x����: ��$,�Pb ���/���� /~/(/:/h/^/p/�/ �/�/�/�/�/V? ?? @?6?H?�?l?~?�?�? �?.O�?�?OO O�O DOVO�OzO�O_�O�O �O�O�Or__._\_R_ d_�_�_�_�_�_�_�f	g�io�pWo�o{d� �o�~o�ozoB�PREF �R��p�p
�IOR�ITY�w[���M�PDSP�q��pwU�T6����ODUC-T3�����;OG��_TG��8���ʯrTOENT �1׶� (!?AF_INE�p,�~7�!tcp7�>_�!udN���?!icmv���֯rXYK�ض���q)� ,�����p��&�	��R�9� v�]�o�����П����@��*��N�`�*�s�K��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE �R��:�w!d��连�2s�9Ks���PORT_N�UM�s�p����_CARTRE�P{p�Ω�SKST�A�w d�LGS6)�ݶ��tӁp�Unothin�g�������{��T?EMP ޾y���'e��_a_seiban�o\��ol� ��}߶ߡ��������� "���X�C�|�g�� ������������	� B�-�f�Q���u����� ��������,< bM�q��������(L�VOERSIyp�w}� disab�ledWSAVE� ߾z	26�00H768S?�!ؿ����/C 	5(�r)og+^/y�e{/�/�/�/�/�*�,/? �p���]_�p 1�Ћ� �����W�h?z?�W*pURGE«�B�p}vgu,�WFF�0DO�vƲ�vW%���4(�C�WRUP_�DELAY ��\κ5R_HOT �%Nf�q׿GO�5R_NORMAL&H��r6O�OZGSEMI�jO�O�O(qQSKI%PF3��W3x=_ 98_J_\_]�_�_{_ �_�_�_�_�_�_	o/o AoSoowoeo�o�o�o �o�o�o�o+= aOq����� ���'��7�]�K��������)E�$RAF{���K/�zĀÁ�_PARAM�A3���K @.�@�`�61�2C<��y��C�6$�B�ÀBTIF�4`�R�CVTMOUu�vc��ÀDCRF3}��I �+UC�AqD��2�=\�(?���]�
�ޅ����4��+_���;��Cd;��.<�߈<�g�<?F+<L���Ѱ��d�u�L������� ϯ����)�;�M��_���RDIO_T?YPE  M=U��k�EFPOS1 ;1�\�
 x4/�����+�$/<�� $υ�pϩ�D���h��� ���'������o�
� ��.ߤ�Rߌ������ ��5���Y���i��*� <�v���r������� ��U�@�y����8��� \�����������?��xc����2 1�KԿX�T�x��3 1�����nY�S4 1�'9K�/�|'/�S5 1����/�/�/�/:/S6 1�Q/c/u/�/�-??Q?�/S7 1��/�/
?D?�?�?�?>d?S8 1�{?�?��?�?WOBO{O�?SM?ASK 1L�8�O�D�GXNO���Fx&�^��MOTEZ�hŻ��Q_ǁ�%]�pA݂��PL_RA�NG!Q]�_QOWE/R �ŵ�P1V�SM_DRYPR/G %ź%"O�_��UTART ���^�ZUME_PR�O�_�_4o��_EX�EC_ENB  x��#�e�GSPD`pO`WhՅjbTDBro�jRM�o�hING�VERSION �Ź#o�)I_AIRPURhP� �O(�MMT_ҡ@T�P#_ÀOB�OT_ISOLC��NTV@A'qhuN�AME�l��o�JO�B_ORD_NU�M ?�X#q�H768  �j1Zc@�r
��rV�s���r�?�r?��r�pÀPC_TI�MEu�a�xÀS2�32>R1�� �LTEACH PENDANw��:GX�!O �Maintena�nce Cons�j2����"��?No UseB�׏ ������1�C�y�V��NPO�P@�YQ��cS�CH_Lf`�%^ �	ő~��!UD1:�z��R�@VAIL�q�@�Ӏ�J�QSPA�CE1 2�ż ��YRs�i�@Ct��YRԀ'{��8�?��˯���� "���7�2�c�u����� G���߯ѿ򿵿�(� �u�AC�c�u����� Ͻ�߿���ϵ��(� �=�_�qσϕ�C߹� �����߱��$��9� [�m�ߑߣ�Q����� �߭��� ���	�W�i� {���M�������5� ��.S�e�w��� ��I������� *?as��E �����/&// ;/]o����� �/2/�/?"?�/7?Y/ k/}/�/�/O?�/�/�?��?�?O0OOKA�o�*SYPpM*��8.30261 �yB5/21/2018 A �WP�fG|�H�_TX`�� !$COMM�E�$US�Ap $EN�ABLEDԀ$sINN`QpIOR�B��@RY�E_SIG�N_�`�AP�AIT\�C�BWRK�BD<��_TYP�CRIN�DXS�@W�@%VF{RI{�_GRPԀ$UFRAM�r�SRTOOL\VMY�HOL�A$LE�NGTH_VTE�BTIRST�T ? $SECLP�X�UFINV_PO�S�@$MAR�GI�A$WAI�T�`�ZX2�\�VG-2�GG1�AI�@�S��Q	g�`_WR�BNO_USE_DI�B^uQ_REQ�BC�C�]S$CUR_T�CQP�R"a^f �G�P_STATUS>�A @ �A3`X�BLk�H$zc1�h��P@���@_�F�X �@E_MLoT_CT�CH_�J6�`CO�@OL�E�C�GQQ$W�@w��b#tDEADLO�CKuDELAY_CNT�a3qGt�a�$wf 2 �R1[1$X<�2*[2�{3[3$Zwy �q%Y�y�q%V�@�c�@��b$V�`�RV�UV�3oh>b�@ � q�d�0arMSKJ��LgWaZ�C`NRK�P�S_RATE�0�$���S
`�Q�TAC���PRD���e�SD*��a4�A�0�DG�A� 0�P�flp bquS2ppI�#`\
`�P 
�S\`�  �A�R_�ENBQ ��$RUNNER_SAXI�<`ALPL�Q��RU�THICQ�$FLIP7��DT�FEREN��R�IOF_CHSU�IW��%V)�G1����$P�řA�Q�Pݖ_J�F�PR_P�	�RV_DATA�A�  $�E�TIM���$VA�LU$�	�OP_ �  �A�  2 �S�C*�	� �$ITP_!�SQ]P�NPOU}�o�TOT�L�o�DSP��JO�GLIb��PE_P�Kpc�Of�i��PX�]PTAS�$KE?PT_MIR��¤2"`M�b�APq�aE�@�y�q�g@١c�vq�PG�BRK6��x���L�I��  �?�SJ�q�P�ADE�z�ܠBSOCz�M�OTNv�DUMM�Y16Ӂ$SV��`DE_OP��S�FSPD_OVR4
���@LD�����OR��TP8�LEb��F������OV��CSF��F����bF��d�ƣ&c)�fQc�LC�HDLY��REC�OV���`��W�PM��gŢ�RO�������_F�?� @v�S� �NVER�@�`O�FS�PC,�CSWD�ٱc�ձ���B����T�RG�š�`E_F�DO��MB_CM4}���B��BLQ�¢�	�Q�̄Vza�BUP��g��G
��AM����@`KՊ�e�_M�!�d�AMf�Q��T�$CA����DF����HBKd�v���I�OU��I'R��PA����������p���~��DVC_DB�S�!�x�Q�!�s�d�9�1�A��9�3A��AT�IO�0��͠��U0S����WaAB��R�+c�`tá`DؾA��_�AUXw�SUBCPUP���S�`�����3Եжc���3�FLyA�B�HW_Cwp�"�Ns&�]sAa��_$UNITS�M�>F�ATTRIz�Z�ެ�CYCL�CNE�CA���FLTR�_2_FI��TARTUPJp����Aƴ�LP������_S�CT*cF_F�F_P���b�FS��+�K�CHA/Q��*�d�RSD��Q�����Q���_TH�PRO8r���հEMPJ���rG�T� ��Q�DI�@y�RAOILAC/�bMX�CLOf�xS��ځ����拁���PR#�S�`app�C� {	��FUNC���RIN`QQP� �ԱRA)]R ���AƠ��AWAR�֓��BLZaWrA0kg�ngDAQ�B�rkLD�र&q��M�K���TI����j��$�@R�IA_SW��AF
��Pñ#��%%�p89r1��MOIQ���gDF_~P(�PD"�LM-�FA�PHR�DY�DORG�H�; _QP�s%MULCSE~Pz���*�� �J��Jײ��FAN_ALMLVG���!WRN�%HARDP��UcO�� K�2$SHADOW�]�kp�a02��� ST�Of�+�_^�w�AU�{`R��eP_SBR�z5���:F�� ��3MPINF?�p\�4��3REGV&/1DG�+cVm �C��CFL(��?�D�AiP���Z`�� �8����Z�	 �P(Q�$�A$Z�Q �V�@�[�
� ���EG��o���kAAR���㌵2�axG���AXE��ROB.��RED��W�QD�_�Mh�SYA��AF�:�FS�GWRI�P~F&�STR����E�˰EEH�)��D�a\2BkPB6P��=V��DvЗOTO�1)���ARYL�tR�v�3����FI&�ͣ$LI�NKb!\��Q�_�3S���E��QXY�Z2�Z5�VOFF����R�R�XxPB��ds�G�cFI�03g�������_J��'�ɲ�S�&qR0LTV[6���aT�Bja�"�bC���D�U�F7�TURB� X��e�Q�2XP�ЊgFL�E���x@��`�U9Z8���� +1	)�K��Mw��F�9��劂����OR!Qj��G;W3��� #�Ґd ���uz����1N�tOVE�q_�M�� ё?C�uEC�uKB�v'0 �x-�wH��t��� & `��qڠ�B�ё�u��q�wh�ECh����E)R��K	�EP�$���AT�K�6e9`e�W���AXs� '��v�/�R ��� �!�� ��P��`�@�`�3p�Yp�1�p �� �� �� (��  8�� H�� X�� h�� �x�� ������DEBU�$%3�I��·RAB���ٱ�s9V��� 
d�J� ����@񘧕������ �Q���a���a��3q���Yq+$�`%"<�cLA�B0b�u�'�GR�O���b<��B_ s��"Tҳ*`�0A�u�p�uq�p1}�ANDGp��������U��p1��  �ѷ0�Qθuݸ��P�NT0���SERsVE �Z@ $`�EAV�!�PO ����nP!�P@�$!�Y@  $.>�TRQ�b
=��B2G�K�%"2\��~� _  l���5�D6ERRVb(�I��V0`;���TOQ:�7�L�@
�R��e %G�%�Q�� <�50�F� ,�`�z��>�RA� 2� d!�����S�  M��pxU �����OCuG�  }��COUNT6Q���FZN_CFG�F� 4#��6��T G4�_�=�����Î�^VC ���M ��"��$6��q ��F!A E� &��X�@� ������A����A9P��P@HEL�0�ҿ 5b`B�_BAS��RSR�6�CSH����1�Ǌ�2��3��4���5��6��7��8��}�ROO����Pf�PNLEA�cAB)�ܫ ��ACKu�IN2O�T��(B$UR0� =�_PU��!0��OU+�Pd�8j���� V��TPFWD�_KAR��� ��R�E(ĉ P�P�>QUE�:RO�p�`r0P1I� x�j�P�8f��6�QSEM��0t��� A��STYL�3SO j�DIX�&p�����S!_TMC�MANRQ��PE�NDIt$KEY?SWITCH����kHE�`BEA�TM83PE{@LEP��>]��U��F���SpDO_HOeM# O�@�EF�p�PRaB�A#PY�C�� O�!���OV_�M|b<0 IOCM��dFQ��k�HKYA D�Q�7��	UF2��M���p�c�FORC�3WARڅ"J�OM|@ G @S�#o0U)SUP�@1�2&3&�4E���T�O��L����8UNLO�v�D4K$EDU1 � �SY�HDD�NF� M�BL�OB  p�S�NPX_AS��� 0@�0��81$�SIZ�1$VA�{���MULTIP�-��# A� � $��� /$4`�BS��0�C���&OFRIFBO�S����3� NF�ODBUP߰�%@3;9(�q����Z@ x��SI��TEs�r�c�SGL�1T�Rp&�Н3B��@�0STM�Tq�3Pg@VBW<�p�4SHOW�5@��SV��_G�� 3p$PCJ�PИ����FB�PHSPb AW�EP@VD�0�WC� ���A00��PB XG XGP XG$ XG5VI6VIU7VI8VI9VIAVIBVI�XG�YF�0XG�FVH��XbI1oI1�|I1�I1�I1�I1��I1�I1�I1�I1��I1�I1�I1Y1�Y2UI2bI2oI2
|I2�I2�I�`�X�I�2p�X�I2�I2�I2*�I2�I2Y2Y�pT�hbI3oI3|I3�IU3�I3�I3�I3�IU3�I3�I3�I3�IU3�I3Y3Y4�iU4bI4oI4|I4�IU4�I4�I4�I4�IU4�I4�I4�I4�IU4�I4Y4Y5�iU5bI5oI5|I5�IU5�I5�I5�I5�IU5�I5�I5�I5�IU5�I5Y5Y6�iU6bI6oI6|I6�IU6�I6�I6�I6�IU6�I6�I6�I6�IU6�I6Y6Y7�iU7bI7oI7|I7�IU7�I7�I7�I7�IU7�I7�I7�I7�IU7�I7Y7T��kVP� UD�y"Dՠ��
<A62��ut�R��CMD� ���M5�Rv�]��Q_h�R���e�����<�YSL���  � �%\2��+4�'���W�BVALAU��b��'���FH��ID_L���HIr��I���LE_���㴦�$0C�SA~C�! h �VE_BLCK���1%�D_CPU 5ɧ 5ɛ �����C��� ��R " � PWj��#0��LA�1SBћì����RUN_FLG �Ś����ĳ ����������H���Х����TBC2��# � @ B��e �S�p8=�FTDC�����V���3d�Q�T!HF�����R�L�?ESERVE9��F��3�2�E��Н��X -$��LE�N9��F��f�RA���W"G�W_5�b�14��д2�MO-�T%	S60U�Ik�0�ܱF����[�DEk�21LgACEi0�CCS#0�� _MA� j��z��TCV����z�T�������.Bi�'AH�z�'AJh�#EM5�"��J��@@i�V�z���2Q �0&@o�h�6��JK��VK9��0{���щ�J0�����JJ��JJ��AAAL���������4��5�ӕ N1�������.�LD�_�1�v�CF�"% `�GROU���1�A�N4�C�#m REQ�UIR��EBU��#��6�$Tk�2�$���zя #�&{ \�APPR� �C� 0�
$OPE=N�CLOS��St��	i�
��&' �MfЩ���W"N-_MG�7CB@��A���BBRK�@NOLD@�0RTMO_5ӆp1	J��P�����@���������6��1�@ m1�#�(� ������'��+#PATH ''@!6#@!�<#� � 9'��1SCA��l�6IN��UCJ�[1� C0@UM�(Y  ��#�"�����*���*���� PAYLOA�~J2LؠR_A	N^�3L��91�)�1AR_F2LSHg2B4LO4�!F7��#T7�#ACRL_@�%�0�'�$��H���.�$HA�2FL�EX��J!�) P�2�D߽߫��|�0��* :�� ��z�FG]D����z���%�F1]A�E�G4�@F�X�j�|���BE�� �����������(� �X�T*�A���@�XI��[�m�\At�T$g�QX <�=��2TX���emX �������������������+	�J>+ �-�K]o|�٠cAT�F�4�ELFP�Ѫs�J� *� J�EmCTR�!�AT�N�vzHAND_VB.��1��$7, $8`F2Avԍ��SWKs�-?� $$M*0. �]W�lg��PZ����A��� 1����:QAK��]AkAzP��LN�]DkDzePZ G��C�ST_hK�lK�N}DY�� � A����0��<7]A <7W1�'��d�@g`�P�������8"Os"�. M�2D�%"p�H��~�ASYIMj%0�� j&-��-W1�/_�{8� �$ �����/�/�/�/ 3J<�:9�/�89�D_VI�v����V_UNI�ӛ��cD1J����╴�W<�� n5Ŵ�w=4��9��?�?<�uc�4�37%�H���/�j��0��DIzuO��8�k�>0 �`��I��A��#���@ģ����@��HQl� �1 � /�MEB.Qp��9�ơT}�PT�;pG �+ /A� ���'��T��0 $DUM�MY1��$PS�_�@RF�@;�$�b�'FLA@ Y�P(c|��$GLB_TP�ŗ���p9 P�q��2 X� �z!ST9�� S�BRM M21_V��T$SV_ERb*0O�p����CL�����AGPO��f�GLv~�EW>�3 4H ��$YrZrW@�x�A1+�A���";��"�U&�4 8`N�Z�"�$GI�p}$&� -� �Y��>�5 LH {��}�$F�E��NEA�R(PN�CF��%PT�ANC�B;�JOG܌@� 6Mp$JOINTwa' d��MSET>�7  "x�E��HQtpS{r��|up>�8� �p�U.Q?�� LOC�K_FOV06���B�GLV�sGLt�T?EST_XM� 3�'EMP����Ҏ_�$U&@%�w`24� Y��5��2�d���3��CE- ����_ $KAR�QM��TPDRA)������VECn@��IUھ�6��HEf�TO�OL�C2V�DREN IS3ER6�N�@ACH� 7?1Ox �Q�29Z�H �I�  @$R�AIL_BOXEzwa�ROBO���?��HOWWA�R�1�_�zROLMj��:qw�jq� ��@ O_Fkp!� d�l>�9�� +�R O8B: �@��c�OU�;��Һ�3ơ�r�q_�/$PIP��N&`H��l�@��#@CORDEDd�p >f��fpO�� < D ��OB⁴sd����Kӕ���qS;YS�ADR�qf���TCHt� =� ,8`ENo��1A�k�_{�-$CqKuP�VWVA��> Ǥ  &��PR�EV_RT�$�EDITr&VSHWRkq�֑ &R:�%v�D��JA�$�a?$HEAD�6�4� �z#KE:�E��CPSPD�&JM%P�L~��0R*P�ģ?��1%&I��S�rC�pNE; �q�wOTICK�C��MJq�3�3HN��@ �@� 1Gu�!_GP8p6��0STY'"x�LO�љ�2l2?�A� t 
m G3%%�$R!{�=��S�`!$��w`���ճ���9Pˠp6SQU��E<��u�TERC�0���TSUtB  ����hw&`gw�Q)�p1O����@IZ��{���^�PR�kюB�1XPU���E_DYO��, XS�K~ƧAXI�@���UR�pGS�r� ^0�&���p_) �ET�BP(m��o��0Fo��0A|���Rԍ���a�p1@R�Cl>@P��b_�yUr� �Y��yU��yS��yS�� �UЇ�U���U���U�] ��Ul[��Y�bXk�]�Cm�����d�S�SC�� D h��DS~0��Q�SPL���eATހ���A�]0,2N�ADDRE�S<B} SHIF�{s��_2CH�pr�I��=q�TVsrI��E"���a�Ce�
��
;�VW�A��'F \��q��0l|\A@�rC�_B"R{z�p�ҩq�TXSCWREE�Gv��1TINA���t{�����A�b?�H T 1�ЂB�����I��Ap��BE�y RRO������� B���d�UE�4I �g�!p�S���RSM]0�GU�NEX(@~Ƴ�j�S_S�ӆ��Á։񇣣��ACY�0� 2-H�pUE;�J���\��@GMT��Lֱ��A��O	�BBL�_| W8���K �Լ0s�OM��LE�/r��� TO!�s�RwIGH��BRD
�%qCKGR8л�T�EX�@����WIDTH�� �B�|�<���I_��Hi� OL 8K���_�!=r���R:�_��HYґ��O6q�Mg0I紐U��h�Rm��LUMh��FpE#RVw��P���`��N��&�GEU�R��FP)�)� LIP��(RE%@�a)ק@�a�!��f �5�6�7�8Ǣ#B�à�@���tP�fW�Sv@M�USR&�OO <����U�Qs�FOC)��P�RI;Qm� :���T�RIP�m�U)N����Pv��0���f%��'���@�0 qQ����AG �0aT� �a>q�OSт%�RPo���8�R�/�A�H�L�q4����U¡�SU�g��¢p5N��OFF���T��}�O�� 1R������S�GUN���6�B_SUqB?���,�SRTN��`TUg2��mCOR�| D�RAUrPE�T<Z�#'�VCC��	3�V AC36MgFB1�%K"PG ��W (#��AST�EM�����0P�E��T3G�X �<\ ��MOVEz�A��AN�� ���M�>��LIM_X��2� ��2��7�,�����ı�
�BVF�`E�+��~��04Y��IB(�7���5S��_Rp� x2��� WİGp+@��}СP��3�Zx ���3A���A�ݠCZ��DRID����V�y08�90� De�MY_UBYd���6�ш@��!��X��P�_S��3��L�KB�M,�$+0DEY�(#EX`�����UM_MU� X����ȀCUS�� ���G0`PACI���а@�Հ:��:,�:����R!E/�3qL�+��:z[��TARG�БP�r��R<�\C d`��A��$�	���AR��SW2 ��-I��@Oz�%qA7p�yREU�U�01�,��HK�2]g0��qP� N� �EAM0GWOR����MRCV3�^ ����O�0M�C�s	p���|�REF_� ��x(�+T� ����������3_RCH4(a�P�І��hrj�NA�5��0�_ ���2����L@��n�@@OU~7wp6����Z��a2[��RE�p�@;0\�c�a'2]K�@SUL��]���C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��Q5(I�]7q�}�Tg`4D�`�0.`0�AP_�HUC�5SA��CMPz�F�6�5�5�0_�aR��a�1I\!yX�9��VGFS��_ad ��M��0p�UF_x��B� �ʼ,RO��Q��'��6��UR�3GR�`.��3IDp���)�D`�;��A��~�IN��H{D���V��J���S͓UWmi=�0����TYLO*�5�����bt m+�cPA� �cCACH�vR�UvQ���Y��p�#CF�I0sFR�XT���Vn+'$HO����P!A 3�XBf�(1 ���$��`VPy� ^b_S�Z313he6K3he1�2J�eh chG�chW�A�UMP�j��IM5G9uPAD�ii�IMRE�$�b_SIZ�$P����0 ��ASYNBUF��VRTD)u5tqΓ?OLE_2DJ�Qu�5R��C��U��vPQ�uECCUlV�EMV �U�r�WVIsRC�aIuVTPG����rv1s��5qMPL�Aqa��v���0�c�m� CKLAS��	�Q�"��d  ��ѧ%ӑӠ@}¾�$8�Q���Ue |�0!�rSr�T�#0! 񕠄r�iI��m�vK�B�G��VE�Z�PK�= �v�Q�&�_HO|�0��f � >��3�@Sp�SLOW�>�RO��ACCaE���!� 9�VR�#0���p:���AD���F��PAV�j�� D����M_B"���^�'JMPG ��g:�#E$SSC��x&�HvPq��hݲvQS�`rqVN��LEXc�Gi T`�sӂ��Qn�FLD �DEsFI�3�02���:��P2�Vj'� �A��V�4[`MV_PIs��t`���A�@��FI��|�Z��Ȥ�����A����A��~�GAߥ1 LsOO��1 JCB�इXc��^`TcPLA!NE��R��1F�c�����pr�M� [`������S����f����A@f��R�Aw�״tU�΁pRKE��d�VA�NC������ �k���ϲ�|"R_AA� l��2� �p�p�#B�m h�@���O K�$������kLЍ0OU&A�"A�Y
p�pSK�TM@F�VIEM 2l p��P=���n <<�x�dK�UMMYK1�P��`DT`M�|!CU��#AU���o $��TIT>�$PR�����OP���VSH�IF�r�p`�J�Q���fOxE$� _R�`UTc���� s��q������G�"�G�޵'�T�$�SC9O{D7�CNTQ i� l�>a�-�a�;�a�H�@a�V���1�+�2u1���D����  ]� SMO�Uq�d�a�JQ�����aI_�R[�r�n�*@�LIQ�AA/`�XV%R��s�n�TL���oZABC�t��t�c�
|!ZIP���u���LVbcL�n"���MPCF�x�v:�$�� �~��DMY_LN��p�����@y�w Ђ�(a�u� MCM�@C>bcCART_�D�PN� $J71D��=NGg08Sg0�BUXW� ��UXEUL|ByX���	��zZ��x 	����m�YH�Db  �y 80���0EgIGH�3n�?(� �H����$z ����|�����$B� K�d'��_��L3�RV�S�F`���OVC �2'�$|�>P&���
q���5D�TR�@ �V�1�SPHX��!{ ,� *�<�$R�B2 2� ���C!��  �@V+| b*c%g!� �b)g"�`V*�,8�?�V+�/V.��/�/?�/�/V(7%3 @/R/d/v/�/6?�/�/ �?�?�?O4OOION;4]?o?�?�?�?SO�? �?�O_�O0_Q_8_f_N;5zO�O�O�O�Op_ �O_o8o�_MonoUo�oN;6�_�_�_�_�_ �oo%o4Uj�r�N;7�o�o�o�o �o� BQ�r�5���������N;8��� ��Ǐ=�_�n���R�टş��ڟN;G �� џ�
����?���W�i�{� ������ï�.��� ����A��dW�<� N�|�������Ŀֿ� ޯ���0�B�_�R� d�꿤϶��������� ����*�L�^��r� ��
�������������&�8�J�l�~� `ҟ @����� ��ߩ��-���� &�,���9�{����� a��������������� A'Y��� �������a#1�
��N;_MODE  �^�S ��[�Y�B���
/\/*�	|/�/R4CWOR�K_AD�	�"��T1R  ����� �/� _INT�VAL�+$��R_OPTION6� �q@V_D�ATA_GRP �27���D��P �/~?�/�?�9��?�? �?�?OO;O)OKOMO _O�O�O�O�O�O�O_ �O_7_%_[_I__m_ �_�_�_�_�_�_�_!o oEo3oioWoyo�o�o �o�o�o�o�o /eS�w��� ����+��O�=� s�a�������͏��� ߏ��9�'�I�o�]������$SAF_DO_PULS� ��~������CAN�_TIM�����ΑR ��Ƙ�5�5�;#U!P"�1!��� �?E�W�i�{��� ��.�ïկ�����V'(~�T"2F�D��dR�I�Y��2�o+@a얿����)��u��� k0ϴ��w_ ��  T� �� �2�D�)�T D��Q�zόϞϰ� ��������
��.�@� R�d�v߈ߚ�/V凷�����߽�|�R�;�o ��W�p��
�t��Diz$� �0 � �T"1!� ���������� ������*�<�N�`� r��������������� &8J\n� ������� "4FX ��࿁ �������/ `4�=/O/a/s/�/�/��/�/�/�/�!!/ �0 ޲k�ݵu�0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ ok$o6o HoZolo~o�o�o�o�o 1/�o�o 2DV hz�/5?���� ����&�8�J�\� n���������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u��� ���`Ò�ϯ�� ��)�;�M�_�q����������˿ݿ� �p���3� ���&2�,��	123�45678v�h!B!��*�Ch���0�ϵ� ���������!�3�9� ��\�n߀ߒߤ߶��� �������"�4�F�X� j�|�h�K߰������� ��
��.�@�R�d�v� ������������� *<N`r�� �����& ��J\n���� ����/"/4/F/ X/j/|/;�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�/�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_�?L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o=_�o�o�o �o�o�o 2DV hz�����h������u�o.�@��R���Cz  B}��   ���}2&� � _��
���  	�_�2�Տ����_�Kp������ď i�{�������ß՟� ����/�A�S�e�w� ��������N����� �+�=�O�a�s����� ����Ϳ߿���'ψ9�K�_������<�v�_��$SCR_�GRP 1
�� �� t� ��� ���	 ������������ ����_������)�a�����&�DE� DW8���l�&�G��CR-35i�A 901234�567890���M-20��8���CR35 ��:�
��������������:֦�Ӧ�G���"&������	��]��o����:��G�H���>���� �������&���ݯ:��j����g������B�t��������r��A����  @�����@� ( ?	�=��Ht�P
��F@ F�`z �y������  �$H��Gs0^p��B��7 ��/�0//-/f/ Q/�/u/�/�/�/8��� P�� 7%?����"?�W?-2?<���@]? H�1�?t�ȭ7�������?-4AA, �&E@�<�@G�B-1 3OZOlO�-:HA�H�O�O|O P�B(�B�O�O_���EL_DEFA�ULT  ��_���S?HOTSTR#]A�7RMIPOWER�FL  i�/U�YTWFDO$V �/URRVENT �1����NU� L!DUM_�EIP_-8�j!AF_INE#P<�_-4!FT�_->��_;o!��`o ��*o�o!RPC�_MAIN�ojh�8vo�o�cVIS�oiiy��o!TPp�PU�Ydk!�
PMON_PR'OXYl�VeZ��2r��]f��!RDM_SRV�r�Yg�O�!R��dk��Xh>���!
�`�M��\i���!?RLSYNC�-9�8֏3�!RO�S�_-<�4"��!�
CE4pMTCO�M���Vkn�˟!	���CONS̟�Wl캟�!��WAS�RC��Vm�c�!���USBd��Xn R���Noӯ������� !��E��i�0���W�RVICE_KL� ?%�[ (%�SVCPRG1���-:Ƶ2ܿ�˰3��	�˰4,�1�˰5�T�Y�˰6|ρ�˰7@�ϩ�˰�����9����ȴf�!�˱οI� ˱��q�˱ϙ�˱F� ��˱n���˱���˱ ��9�˱��a�˱߉� �7߱��_����� ���)����Q�� ��y��'���O��� �w�������� ����˰��İd�c� �����= (as^���� ��/�/9/$/]/ H/�/l/�/�/�/�/�/ �/�/#??G?2?k?V? }?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O�O�O�O	_�O-_���_DEV ~�Y�MC:5X�d�GTGRP� 2SVCP��bx� 	� 
 ,
�PCP5_�_�T�_ �_�_o�_'o9o o]o Do�ohozo�o�o�o�o �o�o5{�_g �������� ��?�&�c�u�\��� ����Ϗ���J\)� ��M�4�q���j����� ˟ݟğ��%��� [�B��f������ٯ �������3��W�i� P���t���ÿ���ο ���A�(�e�L�ί ��RϿ��ϸ������  ��O�6�s�Zߗߩ� ���ߴ������'�~� ��]���h���� ���������5��Y� @�R���v��������� @�	��?&cu \������� �;M4qX� ������/�%/ /I/[/B//f/�/�/ �/�/�/�/�/�/3?? W?�L?�?D?�?�?�? �?�?O�?/OAO(OeO LO�O�O�O�O�O�O�O��O_iV �NLy�6 * 		S=>��+c"_�VU@Tn_Y_B����B�2�J�j�0Q´~_g_�_0Q%�JOGGING��_�^7T(?VjZ��Rf��Y��A�/e�_%o7e�Tt�] /o�o{m�_�o�m?Qi �o�o;)Kq%��o�}os�� ����9�{`�� )���%���ɏ���ۏ �S�8�w��k�Y��� }���ş���+��O� ٟC�1�g�U���y��� ����'����	�?� -�c�Q���ɯ����w� ��s����;�)�_� ����ſOϹϧ����� ����7�y�^ߝ�'� ��ߵߣ�������� Q�6�u���i�W��{� ������=��M��� A�/�e�S���w����� �������=+ aO������u� ��9']� ��M����� �/5/w\/�%/�/ }/�/�/�/�/�/=/"? 4?�/?�/U?�?y?�? �?�??�?9?�?-OO =O?OQO�OuO�O�?�O O�O_�O)__9_;_ M_�_�O�_�Os_�_�_ o�_%oo5o�_�_�o �_[o�o�o�o�o�o�o !coH�o{� �����; �_ �S�A�w�e������� я���7���+��O� =�s�a������П� ����'��K�9�o� ������_���[�ɯ�� �#��G���n���7� ��������ſ���� a�Fυ��y�gϝϋ� �ϯ�����9��]��� Q�?�u�cߙ߇ߩ��� %���5���)��M�;� q�_���߼��߅��� ����%��I�7�m��� ����]����������� !E��l��5� ������_ D�we��� ��%
//��� =/s/a/�/�/�/��/ !/�/??%?'?9?o? ]?�?�/�?�/�?�?�? O�?!O#O5OkO�?�O �?[O�O�O�O�O_�O _sO�Oj_�OC_�_�_ �_�_�_�_	oK_0oo_ �_co�_so�o�o�o�o �o#oGo�o;)_ Mo����o� ���7�%�[�I�k� ���������ُ� ��3�!�W���~���G� i�C����՟���/� q�V������w����� ���ѯ�I�.�m��� a�O���s�������߿ !��E�Ͽ9�'�]�K� ��oϑ�����Ϸ� ���5�#�Y�G�}߿� ����m���i������ 1��U��|��E�� ��������	���-�o� T������u������� ����G�,k���_ M�q���� ���%[I m���	��� //!/W/E/{/��/ �k/�/�/�/�/	?? ?S?�/z?�/C?�?�? �?�?�?�?O[?�?RO �?+O�OsO�O�O�O�O �O3O_WO�OK_�O[_ �_o_�_�_�__�_/_ �_#ooGo5oWo}oko �o�_�oo�o�o�o C1Sy�o��o i�����	�?� �f�x�/�Q�+���Ϗ �����Y�>�}�� q�_�������˟��� 1��U�ߟI�7�m�[� }����ǯ	��-��� !��E�3�i�W�y�ϯ ��ƿ�������� A�/�eϧ���˿UϿ� Q���������=�� dߣ�-ߗ߅߻ߩ��� �����W�<�{��o� ]���������/� �S���G�5�k�Y��� }��������������� C1gU���� ��{����	? -c���S�� ����/;/}b/ �+/�/�/�/�/�/�/ �/C/i/:?y/?m?[? �??�?�?�?? O?? �?3O�?COiOWO�O{O �O�?�OO�O_�O/_ _?_e_S_�_�O�_�O y_�_�_o�_+oo;o ao�_�o�_Qo�o�o�o �o�o'ioN` 9������ A&�e�Y�G�i�k� }�����׏���=�Ǐ 1��U�C�e�g�y��� �֟���	���-�� Q�?�a���ݟ��퟇� �ϯ��)��M��� t���=���9���ݿ˿ ��%�g�Lϋ��� mϣϑϳ�������?� $�c���W�E�{�iߟ� �߯������;���/� �S�A�w�e������ �������+��O� =�s������c����� ������'K��r ��;������ �#eJ�}k �����+Q"/ a�U/C/y/g/�/�/ �//�/'/�/?�/+? Q???u?c?�?�/�?�/ �?�?�?OO'OMO;O qO�?�O�?aO�O�O�O �O__#_I_�Op_�O 9_�_�_�_�_�_�_o Q_6oHo�_!o�_io�o �o�o�o�o)oMo�o A/QSe�����%{,p�$S�ERV_MAILW  +u!��*q~�OUTPUT��$�@�RV� 2�v  $�� (�q�}��SA�VE7�(�TOP1�0 2W� d? 6 *_�π(_������#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u����������Ͽݷ��Y�P��'�FZN_C�FG �u�$�~����GR�P 2�D� ?,B   A[�*q�D;� B\���  B4~�R�B21��HELL���u��j�k��2�����%RSR �������
�C�.�g� Rߋ�v߈��߬������	���-�?�Q��  �_�%Q���(_���,p��⦼�ޖ�g�2,pd�����HK 1�� ��E�@�R� d��������������� ��*<e`r����OMM ������FTOV_�ENB�_���HO�W_REG_UI��(�IMIOFW�DL� �^�)WAIT���$V�1�^�NTIMn���VA�|_)_UNIT����LCTRY�B�
�MB_H�DDN 2W� 2�:%0 �pQ/ �qL/^/�/�/�/�/�/��/�/�"!ON_ALIAS ?e�	f�he�A?S?e? w?�:/?�?�?�?�?�? OO&O8OJO�?nO�O �O�O�OaO�O�O�O_ "_�OF_X_j_|_'_�_ �_�_�_�_�_oo0o BoTo�_xo�o�o�o�o ko�o�o,�oP bt�1���� ���(�:�L�^�	� ��������ʏu�� � �$�Ϗ5�Z�l�~��� ;���Ɵ؟����� � 2�D�V�h�������� ¯ԯ���
��.�ٯ R�d�v�����E���п ���ϱ�*�<�N�`� r�ϖϨϺ���w��� ��&�8���\�n߀� �ߤ�O���������� ��4�F�X�j�|�'�� �����������0� B���f�x�������Y� ��������>P bt����� �(:L�p ����c�� / /$/�H/Z/l/~/)/ �/�/�/�/�/�/? ?�2?D?V?]3�$SM�ON_DEFPR�O ����1 �*SYSTEM*�0m6RECAL�L ?}9 (� �}xyzr�ate 61=>�147.87.1�49.40:93�08  �=102�96 �1�9517�2]?O+M}8co�py virt:�\output\�tcpserv3�.pc md: �over =>3�70278�0357235 �?�O�O�.O@Afrs:or�derfil.d�atCDtmpback\�?�1yO
__��L/?Bmdb:*.*�O�O�O_�_�_67D3x�D:\H_�P�Z_�0s_�_o(o;@4�Ua�_�_�5�_o�o �o<ONO`OrO�o' �O�OU_p_��8_ J_en_��#��_Io [o�_�����4oFoW� jo|���2D�h ��������]��x� 	��.�@�ӏd���� ��,���O�a�t���� )�<�N�ן������ ��U�ޟp����%�8� ˯ݯn� ϑϣ϶�G�@Y��~��!ߴg
�7 ������ ߑߣ߶ey�?�67516�>�o߁��$�dtp?disc 0������������dt�pconn 0 �H�Z�l�~��!��g9 ?�Q�G��������/�0��Z���p���% ����Z������� }5��Pbu��*}<�otes�t_�aer�l16�2791424:263469 � ��2�D�����z/ /���������/�/ .@�dv/�/?�/ ��/�/��/�?�?� ��a?w?�?O-/?/ �?c/�?O�O�O�/P? ]O�/�O_(_;?�O�O q?_�_�_9�K_]_o_��_o$o����27168���_o�o�o�? �?ROSiyo
/OAO��oTh�o��7��$SNPX_AS�G 2�����q� P� 0 '%�R[1]@1.1,��y?�7%�!� �E�(�:�{�^����� ��Տ��ʏ���A� $�e�H�Z���~���џ ����؟�+��5�a� D���h�z�����ů� ԯ���
�K�.�U��� d�������ۿ���� ��5��*�k�N�uϡ� ���ϨϺ������1� �U�8�Jߋ�nߕ��� �����������%�Q� 4�u�X�j������ �������;��E�q� T���x��������� ��%[>e� t������! E(:{^�� ����/�/A/ $/e/H/Z/�/~/�/�/ �/�/�/�/+??5?a? D?�?h?z?�?�?�?�? �?O�?
OKO.OUO�O dO�O�O�O�O�O�O_ �O5__*_k_N_u_�_ �_�_�_�_�_�_o1o oUo8oJo�ono�o�o��d�tPARAM ��u�q W�	��jP�d9p��ht��pOF�T_KB_CFG�  s�u�sOP�IN_SIM  �{vn��p��pRVQSTP_DSBW~r"t��HtSR Zy� � &!pOB1�95_SERV �M���vTOP�_ON_ERR � uCy8�PTN� Zuk��A4�RING_�PR�D��`VC�NT_GP 2tZuq�!px 	r���ɍ���׏��wV}D��RP 1�i p�y��K�]�o� ��������ɟ۟��� �#�5�G�Y���}��� ����ůׯ����� F�C�U�g�y������� ��ӿ��	��-�?� Q�c�uχϙϫ����� ������)�;�M�_� qߘߕߧ߹������� ��%�7�^�[�m�� ������������$� !�3�E�W�i�{����� ����������/ ASew���� ���+=O vs������ �//</9/K/]/o/ �/�/�/�/�/�/?�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?OO�)�PRG_COUNT8v�k�GuKB'ENB��FEMpC:t�}O_UPD 1>�{T  
4Or �O�O�O__!_3_\_ W_i_{_�_�_�_�_�_ �_�_o4o/oAoSo|o wo�o�o�o�o�o�o +TOas� �������,� '�9�K�t�o������� ��ɏۏ����#�L� G�Y�k���������ܟ ן���$��1�C�l� g�y���������ӯ�� ��	��D�?�Q�c��� ������ԿϿ��π�)�;�d�_�q�=L_INFO 1�Eo�@ �2@���������� ����`y*�d��h'��¬���=`y;MYSDOEBUGU@�@����d�If�SP_PA�SSUEB?x�L_OG  ���C���*ؑ�  ���A��UD1:�\�ԘΥ�_MPC �ݵE&�8�A��V�� �A�SAV �!�������X����SVZ�TEM_TIME 1"����@ 0  �f����������$T1SVGUNYS�@VE'�E���ASK_OPTICONU@�E�A�A+��_DI��qOG�BC�2_GRP 2#�I�����@�  �C���<Ko�CFGg %z��� �����`��	�. >dO�s�� �����*N 9r]����� ��/�8/#/\/n/v$Y,�/Z/�/�/H/ �/?�/'??K?]�k? =�@0s?�?�?�?�?�? �?O�?OO)O_OMO �OqO�O�O�O�O�O_ �O%__I_7_m_[_}_ _�_�_�X� �_�_o o/o�_SoAoco�owo �o�o�o�o�o�o =+MOa��� ������9�'� ]�K���o��������� ɏ���#��_;�M�k� }��������ß�ן ��1���U�C�y�g� �������������� 	�?�-�c�Q�s����� �����Ͽ���� )�_�Mσ�9��ϭ��� ����m���#�I�7� m�ߑ�_ߵߣ����� ������!�W�E�{� i������������ ��A�/�e�S�u�w� ������������+ =O��sa��� ����9' ]Kmo���� ���#//3/Y/G/ }/k/�/�/�/�/�/�/ �/??C?��[?m?�? �?�?-?�?�?�?	O�? -O?OQOOuOcO�O�O �O�O�O�O�O__;_ )___M_�_q_�_�_�_ �_�_o�_%oo5o7o Ioomo�oY?�o�o�o �o�o3!CiW ������� ��-�/�A�w�e��� �������я��� =�+�a�O���s����� ��ߟ͟��o�-�K� ]�o�ퟓ�����ɯ����צ��$TBC�SG_GRP 2�&ץ� � �� 
 ?�  6�H�2�l� V���z���ƿ��������(�d��E+�?�	 H�C���>����G����C�  Aq�.�e�q�C��>�'�33��S�/]϶��Y��=Ȑ� C\ g Bȹ��B����>����P���B%�Y�z��L�H�0�$����J�\�n�����@�Ҿ������� ��=�Z�%�7�����?3�����	�V3.00.�	�cr35��	* ����
��������� 3��4�   {�CT�v�}��J2�)����~��CFG +ץ�'� *�������I����.<
�<bM �q������ �(L7p[� �����/� 6/!/Z/E/W/�/{/�/ �/�/�/.�H��/?? �/L?7?\?�?m?�?�? �?�?�? OO$O�?HO 3OlOWO|O�O����O ӯ�O�O�O!__E_3_ i_W_�_{_�_�_�_�_ �_o�_/oo?oAoSo �owo�o�o�o�o�o�o +O=s�E� ��Y����� 9�'�]�K�m������� u�Ǐɏۏ���5�G� Y�k�%���}�����ß şן���1��U�C� y�g�������ӯ���� ��	�+�-�?�u�c� ���������Ͽ�� �/�A�S�����qϓ� �ϧ��������%�7� I�[���mߣߑ߳� �����߷��3�!�W� E�{�i������� ������A�/�e�S� u������������� ��+aO�s ��e�����' K9o]�� �����#//G/ 5/k/}/�/�/[/�/�/ �/�/�/??C?1?g? U?�?y?�?�?�?�?�? 	O�?-OOQO?OaO�O uO�O�O�O�O�O�O_ __M_�e_w_�_3_ �_�_�_�_�_oo7o %o[omoo�oOo�o�o �o�o�o!3�o�o iW�{���� ���/��S�A�w� e�������я����� ��=�+�M�s�a��� ������ߟ�_	�� �_ן]�K���o����� ��ۯɯ���#��� Y�G�}�k�����ſ׿ ��������U�C� y�gϝϋ��ϯ����� ���	�?�-�c�Q�s� u߇߽߫�������� )��9�_�M����/� ���i������%�� I�7�m�[��������� ����������EW i{5����� ���A/eS �w�����/ �+//O/=/_/a/s/ �/�/�/�/�/�/?'? ��??Q?c??�?�?�? �?�?�?�?O�?5OGO YOkO)O�O}O�O�O�O��N  �@S �V_R�$TB�JOP_GRP �2,�E��  ?�V	�-R4S.;\��@�|u0{SPU �>��UT �@�@LR	 �C�� �Vf  C����ULQLQ>�s33�U�R����U��Y?�@=�ZC]��P��ͥR��P  B��W$o/g�C��@g�dDwb�^���ee�ao�P&ff�e=��7LC/kaB �o�o�P��P�efb_-C�p��^g`��d�o�PL�Pt<߿eVC\  �Q@��'p�`�  A��oL`�_wC�?BrD�S�^�]��_�S�`<PB���P�anaa`C�;�`L�w�aQox�p�x�p:��X�B$'tMP@�PCH S��n���=�P��x��trd<M�gE� 2pb����X�	�� 1��)�W���c���� ��������󟭟7�@Q�;�I�w���;d�V�ɡ�U	V3.�00RScr35QT*�QT�A��� E�'E��i�FV#F�"wqF>��F�Z� Fv�RF��~MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
�D���E'
EMK�E���E�ɑ�E�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F��v�F�u�<#�
/<t���ٵ=��_��V ��R�p�V9� ]ES/TPARtp�HFP�*SHR\�ABLE� 1/;[%�SDG�� �W�G�GȡG� WQG�	G�
�G�GȖ�QG��G�G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ�H����w�S]�CS !� ������������ �&�8�J�\�n����� �������� ]\�`�� 	��(�:�����
���.�@�w�NUM�  �EEQ��P	P ۰ܰw�_?CFG 0���)r-PIMEBF_�TTb��CSo�,V�ERڳ-B,R� 11;[ 8$��R�@� �@&  ������ �//)/;/M/_/q/ �/�/�/�/�/?�/? J?%?7?M?[?m?>�@ �?�?�?�?�?�?�?O #O5OGOYOkO}O�O�O �O�O�O�O�O__1_�C_U_g_y_�_�_l_��Y@cY�MI__CHAN8 c} cDBGLV���:cX�	`ETHERAD ?f�\`��?�_uox�oQ�	`ROUTV!	
!�d�o�l?SNMASKQhc>ba255.uߣ�'9ߣY�OOL�OFS_DIb���U;iORQCTROL 2		���~T�����#� 5�G�Y�k�}������� ŏ׏�����.���R�V�PE_DET�AI/h|zPGL_�CONFIG �8�	���/c�ell/$CID?$/grp1V�̟ ޟ����Ӏ�o?� Q�c�u�����(���ϯ ������;�M�_� q�����$�6�˿ݿ� ��%ϴ�I�[�m�� �ϣ�2���������� !߰���W�i�{ߍߟ���%}F�������@/�A�C�i�H�E� �����������?�� .�@�R�d�v������ ����������*< N`r���� ���&8J\ n��!���� �/�4/F/X/j/|/ �//�/�/�/�/�/? ?�/B?T?f?x?�?�? +?�?�?�?�?OO�? >OPObOtO�O�O�O����User �View ��}}�1234567890�O�O�O_#_5_�=T�P��]_���I2 �I:O�_�_�_�_�_�_X_j_�B3�_GoYoko@}o�o�o o�op^46o �o1CU�ovp^5�o�����	�h*�p^6�c�u�����������ޏp^7 R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3��O�M�_�q��������y  e��Yz���	��-� ?�Q���uχϙ�俽�@��������>��e� 5i��c�u߇ߙ߽߫� d������P�)�;�M� _�q��*�<��i��� ������)���M�_� q�������������� ��<�û��=Oas ��>����* '9K]f�Q� ������/� %/7/I/�m//�/�/ �/�/n<��^/?%? 7?I?[?m?/�?�?�?  ?�?�?�?O!O3O�/ <׹��?O�O�O�O�O �O�?�O_!_lOE_W_@i_{_�_�_FOXG9+_ �_�_oo(o:o�OKo po�o)_�o�o�o�o�o( ��	g�0�oM _q���No�� ��o�%�7�I�[�m� &l�n��Ə؏� ��� ��D�V�h��� ������ԟ柍�g� ڻ}�2�D�V�h�z��� 3���¯ԯ���
�� .�@�R���3uF�鯞� ��¿Կ������.� @ϋ�d�vψϚϬϾ� e�w���U�
��.�@� R�d�ψߚ߬����� ������*���w� ��v�������w� ����c�<�N�`�r� ����=�w��-����� *<��`r� ���������  ��1CU gy�������   -/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O�_!_3_E_W_i_� � 
��(  �>%( 	 y_�_ �_�_�_�_�_o	o+o -o?ouoco�o�o�o�Z* �Q &�J\n��� ���o���9�(� :�L�^�p�������� �܏� ��$�6�}� Z�l�~�ŏ����Ɵ؟ ���C�U�2�D�V��� z�������¯ԯ��� 
��c�@�R�d�v��� ��᯾�п�)��� *�<�N�`ϧ����Ϩ� ���������&�8� �\�n߀��Ϥ߶��� ������E�"�4�F�� j�|�������� ����e�B�T�f�x� ������������+� ,>Pb���� ������( o�^p���� ��� /G$/6/H/ �l/~/�/�/�/�// �/�/?U/2?D?V?h?pz?�?�/�`@ �2��?�?�?�3�7�P���!frh:\t�pgl\robo�ts\m20ia�\cr35ia.xml�?;OMO_OqO��O�O�O�O�O�O�O ���O_(_:_L_^_ p_�_�_�_�_�_�_�O �_o$o6oHoZolo~o �o�o�o�o�o�_�o  2DVhz�� ����o�
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟� ݟ��&�8�J�\�n� ��������ȯߟٯ�� �"�4�F�X�j�|��������Ŀ־�8.1� �?@88�?�ֻ�ֿ�3� 5�G�iϓ�}ϟ��ϳ� �������5��A�k��U�wߡ߿��$TP�GL_OUTPU�T ;�!�! ������� �,�>�P�b�t��� �����������(� :�L�^�p�������������2345678901�������� �"��BTf x��4�����
}$L^p ��,>��� / /$/�2/Z/l/~/�/ �/:/�/�/�/�/? ? �/�/V?h?z?�?�?�? H?�?�?�?
OO.O�? <OdOvO�O�O�ODOVO �O�O__*_<_�OJ_ r_�_�_�_�_R_�_�_ oo&o8o�_�_no�o �o�o�o�o`o�o�o "4F�oT|����\��}���� �0�B�T�e�@�������� ( 	 ��Џ������ <�*�L�N�`������� ��ޟ̟���8�&� \�J���n��������� ȯ���"������� *�X�j�F�����|�¿ Կ��C���ϱ�3�E� #�i�{�忇ϱ�S��� �������/ߙ�S�e� ߉ߛ�y߿���;��� ����=�O�-�s�� �ߩ��]�������� '����]�o������ ������E�����5 G%W}������ g���1�U g	w�{��= O	//�?/Q///u/ �/��/�/_/�/�/�/ �/)?;?�/_?q??�? �?�?�?�?G?�?O�? OIO[O9OO�O�?�O �OiO�O�O�O!_3_�O _i_{__�_�_�_�_��_�R�$TPOF?F_LIM >�op>:��mqb�N_SV`  �l�jP_MON7 <6�dop�op2l�aSTRTCHK =6��f� bVTCO�MPAT-h�afVWVAR >Mm��h1d �o ��oop`ba_D�EFPROG �%|j%ROB195_SERV	��j_DISPLA�Y`|n"rINST�_MSK  t|; ^zINUGp�o�dtLCK�|}{QU?ICKMEN�dtoSCRE�p6�~�btpscdt��q��b*�_.�S�T�jiRACE_�CFG ?Mi��d`	�d
?�~u�HNL 2@|i����k r͏ߏ ���'�9�K�]�w�ITEM 2A��� �%$1234567890����  =<��П��  !���p��=��c��^��� �������.���R�� v�"�H�ί��Я��� ���*�ֿ���r�2� ������4�޿�ϰ��� &���J�\�n���@ߤ� d�v��ς������4� ��X��*��@��� ���ߨ�������T� ��x������l��� �����,�>�P����� ��FX��d����� �:�p"� �o�����F 6HZt~��N/ t/�/��// /2/�/ V/?(?:?�/F?�/�/ �/j?�??�?�?R?�? v?�?QO�?lO�?�O�O O�O*O|O_`O _�O 0_V_h_�Ot_�O__ �_8_�_
oo�_@o�_ �_�_Lodo�_�o�o4o �oXojo3�oN�or���o��s�S��B���z�  h��z ��C�:y
 P�v�]�����UD1:\������qR_GRP �1C��� 	 @Cp���$� �H�6�l�Z��|������f���˟���ڕ?�  
���<�*� `�N���r�������ޯ ̯��&��J�8�Z����	�u�����sS�CB 2D� �����(�:�L��^�pς��|V_CONFIG E����@����ϖ�OUT?PUT F�������6�H�Z� l�~ߐߢߴ������� �����#�6�H�Z�l� ~������������ ��2�D�V�h�z��� ������������
� .@Rdv��� ����)< N`r����� ��//%8/J/\/ n/�/�/�/�/�/�/�/ �/?!/4?F?X?j?|? �?�?�?�?�?�?�?O O/?BOTOfOxO�O�O �O�O�O�O�O__+O >_P_b_t_�_�_�_�_ �_�_�_oo'_:oLo ^opo�o�o�o�o�o�o �o $����!�b t������� ��(�:�-o^�p��� ������ʏ܏� �� $�6�G�Z�l�~����� ��Ɵ؟���� �2� D�U�h�z�������¯ ԯ���
��.�@�Q� d�v���������п� ����*�<�M�`�r� �ϖϨϺ�������� �&�8�J�[�n߀ߒ� �߶����������"� 4�F�W�j�|���� ����������0�B� S�f�x����������� ����,>Pa� t��������(:L/x���k}gV� K���//&/8/ J/\/n/�/�/�/W�/ �/�/�/?"?4?F?X? j?|?�?�?�?�/�?�? �?OO0OBOTOfOxO �O�O�O�?�O�O�O_ _,_>_P_b_t_�_�_ �_�O�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����o� ��� �2�D�V�h� z��������ԏ��� 
��.�@�R�d�v��� ������Ϗ����� *�<�N�`�r������� ��˟ޯ���&�8� J�\�n���������Ż��$TX_SCR�EEN 1G�g�}�ipnl/��gen.htmſ�*��<�N�`ϽPa�nel setupd�}�dϥϷ����������ω�6�H� Z�l�~ߐ�ߴ�+��� ����� �2�߻�h� z������9�g�]� 
��.�@�R�d���� �����������}� ��<N`r�� ;1��&8 �\��������QȾUALRM_MSG ?��� �Ȫ-/?/ p/c/�/�/�/�/�/�/��/??6?)?Z?%S�EV  -��6"ECFG �I��  �ȥ@�  A�1 �  B�Ȥ
  [?ϣ��?OO%O7O IO[OmOO�O�O�G�1�GRP 2J�;; 0Ȧ	 �?�O� I_BBL_N�OTE K�:T��lϢ��ѡ�0RDEF�PRO %+ (%N?u_Ѡc_�_�_ �_�_�_�_o�_o>o�)oboMo�o\INU?SER  R]�O��oI_MENHI�ST 1L�9  �(�0 ���)/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,1133�,1�oDVhz~�s� }9361 �����r�$�6� H�Z�l�~������Ə ؏����� �2�D�V� h�z�	�����ԟ� ��
���.�@�R�d�v� �������Я���� �9Rq��B�T�f�x� ��������ҿ���� ϩ�>�P�b�tφϘ� '�9���������(� ��L�^�p߂ߔߦ�5� ������ ��$���� Z�l�~����C��� ����� �2��/�h� z��������������� 
.@��dv� ����_� *<N�r��� ��[�//&/8/ J/\/��/�/�/�/�/ �/i/�/?"?4?F?X? C�U��?�?�?�?�?�? �/OO0OBOTOfO�? �O�O�O�O�O�O�O�O _,_>_P_b_t__�_ �_�_�_�_�_�_o(o :oLo^opo�oo�o�o �o�o�o �o$6H Zl~i?{?��� ���2�D�V�h� z����-�ԏ��� 
����@�R�d�v��� ��)���П����� ����N�`�r������� 7�̯ޯ���&����J�\�n�����������$UI_PAN�EDATA 1N����ڱ  	�}������!�3�E�W� ) Y�}�7�뿨Ϻ����� ���i�&��J�\�C� ��gߤߋ������������"�4��X�7�� �q}�ϕ��� ������B����%�I� [�m������
����� ������!E,i {b������l�ܳ7�<N` r����-��� //&/8/�\/n/U/ �/y/�/�/�/�/�/? �/4?F?-?j?Q?�?�? %�?�?�?OO0O �?TO�xO�O�O�O�O �O�OKO_�O,__P_ b_I_�_m_�_�_�_�_ �_oo�_:o�?�?po �o�o�o�o�oo�o  sO$6HZl~�o ������� � 2��V�=�z���s��� ��ԏGoYo�.�@� R�d�v�ɏ����П ������<�N�5� r�Y�������̯��� ׯ�&��J�1�n��� ����ȿڿ���� c�4ϧ�X�j�|ώϠ� ����+��������0� B�)�f�Mߊߜ߃��� ����������P� b�t���������� S���(�:�L�^��� ��i�����������  ��6ZlS�0w�'�9�}��� "4FX)�} ��l�����/ j'//K/2/D/�/h/ �/�/�/�/�/�/�/#?�5??Y?��C�=��$�UI_POSTY�PE  C�� 	 e?��?�2QUICKM_EN  �;�?��?�0RESTOR�E 1OC�  �L?B��6OCC1O��maO �O�O�O�O�OuO�O_ _,_>_�Ob_t_�_�_ �_UO�_�_�_M_o(o :oLo^oo�o�o�o�o �o�oo $6H �_Ugy�o��� ��� �2�D�V�h� �������ԏ�� ��w�)�R�d�v��� ��=���П������ *�<�N�`�r����� ���ޯ���&�ɯ J�\�n�������G�ȿ�ڿ�����7SCR�E�0?�=�u1sc+@u2�K�3K�4K�5K�6�K�7K�8K��2UScER-�2�D�ksMê��3��4��5��6ʬ�7��8���0ND�O_CFG P�;� ��0PDAT�E ����None�2��_I�NFO 1QC�@��10%�[���I� ��m߮��ߣ������� ���>�P�3�t��i�����<-�OFFSE/T T�=�ﲳ $@������1�^�U� g�������������� ��$-ZQcu����?�
����U�FRAME  ���*�RTOL_ABRT	(�!�ENB*GRP� 1UI�1Cz  A��~��~ ���������0UJ�9MS�K  M@�;N%8�%��/�2oVCCM��V��V�#RG�#Y�9����/����D�BH��p71C����3711?�C0�$MRf2_�*S�Ҵ��	���~XC�56 *�?�6����1$�5���A�@3C��. ��8�?��OOKOx1FOsO�5�51���_O�O�� B����A2�DWO�O 7O_�O8_#_\_G_�_ k_}_�__�_�_�_�_�"o�OFoXo�%TCC��#`mI1�i������� GFS��2�aZ; �| 23�45678901 �o�b�����o�� !5a�4BwB�`56� 311:�o=L�Br5v1�1~1�2�� }/��o�a��#� GYk}�p��� ����ُ�1�C�U� 6�H���5�~���ߏ����	���4�dSEL#EC)M!v1b3��VIRTSYNC��� ���%�SI?ONTMOU�������F��#b�����(u FR:\H��\�A\�� �߀ MC��LO�G��   UD�1��EX����'� B@ �����̡m��̡  O�BCL�1�H� ��  =	 �1- n6  G-������[�,S�<A�`=��͗���ˢ��TRAIAN⯞b�a1l�
0�d�$j�T2cZ; (aE2ϖ�i��;� )�_�M�g�qσϕϧπ�������	��F�S?TAT dm~2!@�zߌ�*j$i߾߮�_GE�#eZ;��`0�
� 02���HOMIN� f������ P~�����БC�g�X����JMPERR {2gZ;
  �� *jl�V�7�������� ������
��2�@�q�hd�v�B�_ߠRE� �hWޠ$LEX��i�Z;�a1-e��VM�PHASE  �5��c&��!OFFX/�F�P2n�j�0�㜳E1@���0ϒE1!1?s33�����ak/�k�xk䜣!W�m[�� ���[����o3;� [i {����/ �O�?/M/_/q/� �/��//�/'/9/�/ =?7?I?s?�/�?�/�/ �?�??Om?O%O3O EO�?�?�O�?�O�O�? �O�O�O__gO\_�O E_�O�_�O�O/_�_�_ �_oQ_Fou_�_|o�o �_�oo�o�o�o�o;o Mo?qof-�oI� ����7�[ P���������ˏ ��!�3�(�:�i�[��ŏg�}������TD�_FILTEW�n��� �ֲ:��� @���+�=�O�a�s� ��������֯��� ��0�B�T�f�x����SHIFTMENoU 1o[�<��%��ֿ����ڿ�� ��I� �2��V�hώ� �Ϟϰ�������3�
��	LIVE/S�NAP'�vsf�liv��E��^��ION * Ub�h�menu~߃��`���ߣ���p����	����E�.�5T0�s�P�@� ���AɠB8z�z���}��x�~�P��c ���MEbЩ��<�0���M�O��q���z�W�AITDINEN�D������OK�1�OUT���S�D��TIM����o�G���#���C����b������REL�EASE������T�M�������_A�CT[�����_D?ATA r���%L����xRDI�Sb�E�$XV�R�s���$ZA�BC_GRP 1Ut�Q�,#�0�2���ZIP�u�'�&����[M�PCF_G 1v��Q�0�/� wx�ɤ� 	�>Z/  85�/0�/H/�/l$?��+�/ �/�/?�/�/???r?>�?  �D0�? �?�?�?�?�;����x�]hYLINuD֑y� ��� ,(  *VO�gM.�SO�OwO�O�M i?�O�O^PO1_�O U_<_N_�_�O�_�_�_ _�_�_x_-ooQo8o`�_�o�oY&#2z�� ���oC�e?�a?>N|�oq�����qA�$DSPHE_RE 2{6M��_ �;o���!�io| W�i��_��,��Ï�� �Ώ@��/�v���e� ؏��p���������l�ZZ�� �N