��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  !�  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d�APP�INFOEQ/ � �L A 8�!�%�! H� �&��)EQUIP w3� NAMr {�'2_OVR�$VERSI3 �� PCOUPL�ED� $!P{P_� CES0s!�_81F3K2> �!� � $SOF�T�T_IDk2TOTAL_EQs 3$�0�0NO�2U �SPI_INDE�]�5Xk2SCRE�EN_(4_2SI�GE0_?q;�0P�K_FI� 	�$THKYGPA�NE�4 � DU/MMY1dDDd!�OE4LA� R�!R��	 � $T{IT�!$I�� N �Dd�Dd �Dc@�DU5�F6�F7�F8�F9�G0�G�GJA�E�G(bA�E�G1�G1�G �F�G2�B!SBNw_CF>"
 8F CNV_J� ; �"��!_CMNT�?$FLAGS]��CHEC�8 � E�LLSETUP {� $HO30�IO�0� %�SM�ACRO�RREP	R�X� D+�0��R�{�T UTOBA�CKU�0� �)DEVIC&�CTI*0�� �0�#�`B�S$IN�TERVALO#I?SP_UNI�O`�_DO>f7uiFR3_F�0AIN�1����1c�C_WAxkda�jOFF_O0]N�DEL�hL� p?aA�a1b?9a��`C?��P�1E���#sATB�d���MO� �cE �D [M�c��^qR;EV�BILrw!�XI� QrR � � OD�P�q_$NO^PM�Wp�t�r/"�w� ��u�q�r�0D`S� p E RD�_E�pCq$FS�SBn&$CHKBoD_SE^eAG �G�"$SLOT!_��2=�� V�d�%���3 a_ED�Im   � )�"��PS�`(4�%$EP�1�1$�OP�0�2�a�p_�OK�UST1P_�C� ��d��U �PLACI4!�Q�4�<( raCOMM� ,0$D����0�`���EOWBn�IGALL;OW� (K�":(2�0VARa��@h�2ao�L�0OUy�� ,Kvay��PS�`�0M_O]�����CCFS_U	T~p0 "�1�3�#��ؗ`X"�}R0 { 4F IMCM�`O#S�`��upi �	_�p�B}�a����M/ h�pIMPEE_F�N���N���@O��r�D_(�~�n�Dy�F� d�CC_�r0  aT� '��'�DI�Pn0"��p�P줇$I������Fn�t X� GRP0���M=qNFLIx�7��0UIRE���$g"� SWITC�H5�AX_N�PS~s"CF_LIM�� � �0EED��!��qP�t�`�PJ_dVЦMOD�Eh�.Z`�PӺ�ELBOF� ���� ��p� ���3���� �FB/��0�>�G�� �� WARNM�`/��qP���n�NST� CORz-0bFLTRh�/TRAT�PT1�� $ACC1a��N |��r$ORI�lo"V�RT�P_S�� CHG�0I���rT2��1�I��T�I1��� x� i#�Q��HDERBJ; CQ�2L�U3L�4L�5L�6L��7L�8L�9{5CO`S <F +�=��O��#92��LLEC�y�"MULTI��b�"N��1�!���0T��� �STY �"�R`�=l�)2`�p���*�`T  |�  �&$��۱m��P�Ḻ�UTO���E��EXT����ÁB���"2� (䈴![0������<�b+��� "D"���ŽQ���<煰kc�q(�9�# ���1��ÂM�ԽP���" '�3�$ L� E���P<��`=A�$JOBn�T����l�TRIG3�% dK�������<���`\��+�Y�p�_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`�0Z���0��P_�P��n@ ( @F RO.���&�t�IT�c�NOM�
����S���`T)w@���Z�1P�d���RA�0��p2b"����
$T��.��MD3�T��`QU31���p(5!HGb��T1�*E�7��c�KAb�WAb�cA4#Y�NT���PDBG�D�� *(��PU�t@X��W���AX���a��eTAI^cB�UF��0!+ g� 7n�PIW��*5 P�7M�8M�9
0�6F�7SIMsQS@>KEE�3PATn�^�a" 2`#��"�L64FIX!, ���!d��D�12Bus=CCI�:FgPCH�P:BAD렀aHCEhAOGhA]HW�_�0>�0_h@�f�Ak� ��F�q\'M`#�"�:DE3�- l�p3G@��@FSOES]FgH�BSU�IBS9WC��.� ` ��MARqG쀳��FACLp�SLEWxQ�e�ӿ��MC��/�\pSM_JB M����QYC	g�e���Д0 ā�C�HN-�MP�$G� Jg�_� #���1_FP$�!TC uf!õ#�����d�#a���V&��r�a;�fJ�R���rSEGFR�PIO� STReT��N��cPV5���!41�r��
r>�İ�b�B�O�2` +�[���,qE` &�,q`y�Ԣ}t��yaSIZ%���t�v�T�s� �z�y,qRSINF}Oбc���k ��`��`�`L�ĸ �T`7�CRCf�ԣCC/�9��`a�uah�ub'�MIN��uaDs�T#�G�D�YC��C������e�q0��� �E�V�q�F�_�eF��N3�s�ah��Xa+ep,5!�#1�!OVSCA?� A��rs1�"!3 ��` F/k��_�U��g��]���C�� a�s�ﳠR>�4� �����N����5a�R�HA;NC��$LG��P�6f1$+@NDP�t�AR5@N^��a�q���c��ME�18���}0f��RAө�AZ �𨵰�%O��FCT K��s`"�S�PFADIJ�OJ�ʠ� ʠ���<���Ր��qGI�p�BMP�dp�p�Dba��AES�@�	�K�W_��BAS��� �G�5  zM�I�T�CSX[@�@�!62�	$X����T9�{sC��N��`�a~P_HEIG9Hs1;�WID�0�aVT ACϰ�1�A�Pl�<���EXP�g���|��CU�0M�MENU��7�T[IT,AE�%)��a2��a��8 P,� a�ED�E ��wPDT��REM.���AUTH_KEGY  ������ ��b�O	�!}1ERR9LH� �9 \� �q�-�OR�DB�_IDx�@l �PUN_O��>Y�$SYS0��4�g�-�I�E�EVx�#��(�PXWO��z �: $SK7!tf2%�Td�TRL��7; �'AC�`��nĠIND9DJ.D��_��f1��f���kPL�A�RWAj�D��SD�A��!+r||��UMMY9d҆F�10d�&���J�<��}1PR� 
�3�POS��J�= ��$V$�q�PL~�>���SܠRK�?����CJ�@����ENE�@T���A���S_�RECO}R��BH 5 �O�@=$LA�>$~�r2�R��`�q�bf`�_Du��0RO�@�aT[�Q��b������! }У�PAUS|���dETURN�򖒃MRU�  C�Rp�EWM�b�AG�NAL:s2$LAx�!?$PX��@$P�y A� �Ax�C0 #ܠD�O�`X�k�W�v�q�G�O_AWAY��M�O�ae���]�CSS_CCSCB �C �'N��CER�I��гJ`u�QA�0�}��@�GAG� R�0�`��{`��{`OF�q�5X��#MA��X���A��LL�D� �$���sU�D�)E%!`���OVR310W�,�OR|�'�?$ESC_$`�eDSBIOQ��l q��B�VIB&� �c,�����f�=p�SSW���f!VL���PL���ARMLO
��`����df7%SC �bALspH�MPCh �Ch P�#h �#h 5�UU� ��C�'�C�'�#�$'�d�#C\4�$�pH���Ou��!Y��!�SB ���`k$4�C�P3�Wұ46$VOL�T37$$`�*��^1��$`O1*�$,o��0RQY��2b4~�0DH_THE�����0SЯ4�7ALPAH�4�`���7�@ �0T�qb7�rR�5�8 8� ×���"��JFn�MӁVHBPFUAFLQ"D�s�`�THR��i2dBP�����G(��PVP������������1�J2`�B�E�C�E�CPSu� Y@��Fb3���H�(V �H:U�G�
X0��FkQw�[�Na�'B���C �INHBcFILT���$��W�2�T 1�[ ��$����H YАAF�sDO ��Y�Rp� fg�Q� +�c5h�Q�iSh�Q�PL���Wqi�QTMOU�#c�i�Q\��X@�gmb��vi�h�bAi�fI�aHIG��caB	xO��ܰ��W�"v�AN-u!��	#AVj�H!Pa8$P�(ד#p�R_:�A�a��T"�N0�X�M�CN���f1[1�qVAE�p��Z2;&f�I�Q�O�u�rx�wGldDEN{G|d��aF>�!�9��aM:�U�FW	A�:�Ml���X�Lu���$!����!l�ZO ����0%O�lF�s�1&3�DI�W�@���Q���_��!CUgRVA԰0rCR41ͰZ�C<�r�H�v����<�`��<�(�f�CH �QR3�S���t���Xp�VS_�`�ד��F��ژ�����&шNSTCY_� E L����1��t�1��U��24�2
B�NI O7�������DEVI|� Fv��$5�RBTx�SPIB�P���B�YX����T��H�NDG��G H !tn���L��Q��C���5��Lo0 �H��閻�FBP�{tFE{�5�t��T4��I�DO���uPMCS�v>�f>�|t�"HOTSW�`�s�%҈ELE��J T���e�2��25�2� O� ��HA7�E�8�344�0RS:����A�K �� MDL^� 2J~PE�� 	A��s��tːÈ�s�JÆG!��rD"�óɘ����\�TO��W�	x��5�?SLAV��L  \0INP�ڐ���`%ن_CF~d�M� $��7ENU��OG��b�0ϑ]զP�0`ҕ�]�IDMA�Sa��\�WR�#��"]�V�E�$a�SKI�ST�s��sk$��2u���J �������	��Q����_SVh�EXCLqUMqJ2M!ONL��"D�Y��|�PE ղ�I_V�APPL9YZP��HID-@Y��r�_M�2��VR�FY�0��r�1�cIGOC_f�� 1��d����O��u�LS����R$DUMMY�3�!���S� L_TP/Bv�"���A�|��ّ N ����RT_u�� ��G&r[�O D���P_BA�`��3x�!F ��_D5���H��\�A�P��>�� P $4 Kw�ARGI��� q�{2O[�_SGNZ��Q �~P/�/PIG!Ns�l�$�^ sQ�ANNUN��@�T<�U/�ߴ�LAzp]	Z�d~>�EFwPI�@ Rk @�F?IT�?	$TOTA%��Pd���!�M�NIY�S+���E��A[�
DAYS\�ADx�@��	�� �EFF_AX�I?�TI��0zCO�JA �ADJ_�RTRQ��Up���<P�1D �r5̀Ll�T�p? ]P�"�p��mtpd��V �0w�G���������SK�SU� ��CTRL_CA��� W�TRAN�S�6PIDLE_�PW���!��A�V曧V_�l�V ��DIAGS���X�� /$2�_SE�#TAC���t!`�!0z*@��RR��vPA���p ; SW�!�!�  ��ol��U��oOH��P�P� ��IR�r��BcRK'#��"A_Ak� ��x 2x�9ϐZs2��%l�W�pt*�x%oRQDW�%MSx��t5AX�'�"��LI�FECAL���10��N�1{"�5Z�3�{"dp5�ZU`}�MO�TN°Y$@FL9A�cZOVC@p�5�HE	��SUPP!OQ�ݑAq� Lj (CL�1_X6�IEYRJZRJWRJ�0TH�!UC|��6�XZ_AR�p6��Y2�HCOQ��MSf6AN��w$��ICTE�Y `>��CACHE�Cp9�M�PLAN��oUFFIQ@�Р�0<�1	��6
���MSW�EZ 8>w KEYIM�p��TM~�SwQq�wQ�#����OCVI�E� �[ A�B�GL��/�}�?� Q	�?��D\p�ذST��!�R� �T�� �T� �T	��PEM�AIf�ҁ��_/FAUL�]�Rц��1�U�� �T�RE�^< �$Rc�uS�% IT��BUFW}�Wr��N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTQT����sP��M��OtT�LwAX � ��X~`9#�c_G�3
?A�DYN_1�E_�D��1 �2UM���T�F���H@ g�`�� 0p��Gb-sC_R�AIK���r�t��RoQ�u7h�qDS�Pq��rP��A�IM@�c6�\����s2�U�h@�A�sM*`IP��d�s�!DҐ6�TH�@�n�)�OT�!6�HS{DI3�ABSC���@ Vy��� �{_D�CONVI�AG���@3�~`F�!pd��psqSC8Z"���sMERk��qcFB��k��pET����aeRFU:@DUdr`����x�CD,�P��@p;cHR�A!���bp�ՔՔ+PUSԕC��C��p�QғSp�cH *�LX�:cd� Rqa�| ����W��U� �U��U�	�U�OQU�7R�8R�9R��0T��^�1k�1x�1��1���1��1��1��1Jƪ2Ԫ2^�k�2x�U2��2��2��2��U2��2ƪ3Ԫ3^�	3k�x�3���o���U3��3��3ƪ4Ԣ�%�XTk!0�d <� 7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr�¸��䂴2REM� F�j��BOVM��A��TROV�DTl�`-�MX<�IN�8�0,�W!INDKЗ�
w�׀�p$DG@~q36��P�5�!D��6�RIV�����BG�EAR�IO�%K�¾DN�p��J�82���PB@�CZ_MCM��@�1��@U��1�f� ,②a? ����PI�!?I�E��Q�TQ�am��©g� _0Pfqg R�I9ej�k!UP2_� h � �cTD��p���! a�����BAC�ri T��P�b�`�) OG���%���p��IF�I�!�pm�>��	�PyT�"}�FMR2��j ��Ɛ+" ����\��������$�(B`x%��_ԡ�ޭ_���� M�������DGCLF�%DG�DY%LDa��5��6�ߺ4@��Uk�~�� T�FS#p�Tl P���e�qP>�p$EX_��B�1M2��2� 3��5��G ���m Y��Ѝ�SW�eOe6DEBUG���%�GR���pU�#BK�U_�O1'� �@PO�I5�65MS��OOfswSM��E�b���0��_E n �p�� �TERM�o�Q��ORI�+�p�@�@SM�_���b�q�/��TA�r�U}P�Rs� -�1θ�n$�' o$�SEG,*> ELT}O��$USE�pNFIAU"4�e1����#$p$UFR����0ؐO!�0����OT�'�TAƀU�#wNST�PAT��<P�"PTHJ�����E�P r�PV"ART��``%B`�abU!REyL:�aSHFT���V!�!�(_SH+@M�$���� ��@N8r�����OVRq��rSSHI%0��UN� �a�AYLO����qI�l����!�@��@ERV]��1�?:�¦'��2��%��5�%�RC<q��EASYM�q�EFV!WJi'��}�E���!I�2��U@D��q�%Ba��
5Po��0��p6OR�MY� `G	R��t2b5n� �� ��UPa�Uu �t�")���TOCO!1S�1POP ��`P�pC�������Oі�`REPR3��aOX�P�b�"ePR�%�WU.X1��e$PW�R��IMIU�2R_	S�$VIS��#(A�UD���Dv" vΥ�$H���P_AWDDR��H�G�"�Q�Q�QБR~pDp1�w H� SZ�a���e�ex�e��SE؄�r��HS��MN~vx �0��%Ŕ��OL���p�<P��-��ACROxlP_!QND_C���ג�1�T �ROUP$T��B_�VpQ�A1Q�v��c_��i���i ��hx��i���i��v�ACk�IOU��D��gfsu^d�y $|�P_D��VB^`bPRM_�b���HTTP_אH�az (��OBJ�Er��P��$��L�E�#�s`{ �s ��u�AB_x��T~�S�@�DBwGLV��KRL�Y�HITCOU�B�GY LO a�TEM��e�>�+P'�,P�SS|�P�JQUE�RY_FLA�b��HW��\!a|`�u@�PU�b�PIO ��"�]�ӂ/dԁ=dԁ~�� �IOLN���}����CXa$�SLZ�$INP7UT_g�$IP#�1P��'���SLvpa~��!�\�W�C-�B��qIO�pF_AS:v��$L ��w� �F1G�U�B0m!0���0HY��ڑv��HO��UOPs� `������[�ʔ[�і"�[PP�SIP��<�іI�2�dat�IP_MEMB��ni`� X��IP�P�b{�_N�`�����R�����bSP���p$FOCUS�BG�a~�UJ�Ƃ� �  � o7JO�G�'�DIS[�JY7�cx�J8�7� �Im!�)�7_LA�B�!�@�A��AP�HIb�Q�]�D�� J7J\���� _�KEYt� ��KՀLMONa���$XR��ɀ��?WATCH_��3L���EL��}Sy~�L��s� �Ю!V�g� �CTR3򲓥v��LG�D� �R����I�
LG_SIZ���J�q IƖ�I�FDT�IH�_�jV� GȴI�F�%SO���q  �Ɩ���v��ƴ��K�AS����w�k�N�
���E��\����'�*�U�s5��@L�>�4�DAUZ�EA`�pՀ�Dp�f�GH�Bܶq��BOO��g� C���PIT����� ��REC��S'CRN����D_p�b�aMARGf�`��@:���T�L���S�s¡�W�Ԣ�Iԭ�JG=MO�MNCH�c���FN��R�Kx�PR�Gv�UF��p0��F�WD��HL��STP��V��+���Є�RS��H�@�몖C�r4��?B��� +�O�U �q��*�a28����Gh�0PO������b��M8�Ģ��EX���TUIv�I��(� 4�@�t�x�J0@J�~�P��J0��N�a��#ANA��O"�0V�AIA��dCLEA�R�6DCS_HIP"�/c�O�O��SI��S��I�GN_�vpq�uᛀTܓd� DEV-�LL�A �°BUW`�j�x0T<$UǃEM��Ł����0�A
�R��x0�σ�a��@OS1�2�3��x�c�`� ��ࠜh�AN%-���-�IKDX�DP�2MRO�X�Գ!�ST��Rq��Y{b! �$E&C+��p.&A&8`��a� L��ȟ@%Pݘ��T\Q�UE�`�U c��_ � �@(��`�b����# �MB_PN�@ R`r��R�w�TR�IN��P��BAS8S�a	6IRQ6�q{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?(�?RIAt�� ID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCES�?R,1�AMhPa�͠�BD4+2�A�q`5�`�F_A�J��C[�O�H� K��� �\���bTf$� ��L�I�q�SREQUIRE�#MO�\�a�XODEBU��,1L� M䵔 �p���P(�c�AA,1N��
Q��q�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N��iPST9� �� 4��LOC�R�I���EX�fAN�G��A,1ODAQ䵗�@$��9�ZMF�����f��"��p�%u#ЖVSUP�%v+1FX�@IGGo�� �rq�"��1� �#B��$���p%#by���rx���vbPDATAK�pE;����Rr��M��*� t�`+MD�qI��)�v� ��t�A�wH�`��tD�IAE��sANSW���th���uD��)�AOԣ(@$`� PCU_�V6�ʠ�d&�PLOr�$`�R���B���B�p������RRR2�E��  ��V�A/A ?d$CALI�@��	G~�2��!V��w<$R�SW0^D�"��ABC�hD_�J2SE�Q�@�q_�J3M�
G�1SPH�,��@PG�n�3m�(u�3p�@��JkC��4�2'AO)IMk@{BCSKP^:ܔ9�wܔJy�{BQܜ��8���`_AZ.B���?�EL��YAOC�MP�c|A)��RT�j���1�ﰈ��@�1�������Z��S�MG��pԕ� ERl!��aINҠACk�p����b�n _�������{A��/R��DI�U�'�DH�@
�#a��q$V�Fc�$x�$���`@���b��̂�E�H? �$BELP�����!ACCEL����kA°IRC_R��pG0�T!��$PS�@B2L+0 ���W3�ط9� ٶPATH��.�γ.�3���p�A_��_��e�-B�`C���_M=G�$DD��ٰ��$FW�@�p�����γ����DE��P�PABN�ROTSPEEu��O0��DEF>Q��+0?$USE_��J%PQPC��JY����Z-A 6qYN�@A�pL�̐�L�MOU�3NG��|�OL�y�INCU��a�¢ĻBx��ӑ�AENCS����q�B�����D�IN��I�����pzC�V�E�����23_Ux ��b�LOWL�A��:�O0��0�Di�@�B�PҠ� ��PRC�����MOS� gTMO�pp�@-GPERCH[  M�OVӤ �� ���!3�yD!e�]��6�<�� ʓA����L IʓdWɗ��:p3�.��I�TRKӥ�AY ����?Q^���m�b��`pp�CQ�� MOM��B?R�0u��D���0y�0Â��DUҐZ��S_BCKLSH_C����o�n��T������
c��CLALJ��A��/PK�CHKO0�Su�RTY� �q��M�1r�q_
#c�_UMCPr�	C���SCL�n��LMTj�_L�0X����E�� � � ���m�h���L6��PC����H� ��P�ŞCN@�"XT\����CN_��N^CL�kCSF����V6Ҁ���ϡj���nCAT�SHs���� �ָ1���֙�������f��PA���_P���_P0� e���O1u��$xJG� P{#��OG���TORQU(�p�a�~����Ry������"_W��^���@��4t�
5z�
5I;I ;Iz�F�`�!��X_8�1��VC��0�D�B�21�>	P�?�B�5�JRK�<�2�6i�D�BL_SM�Q&BM�D`_DLt�&BGR�V4
Dt�
Dz��1H�_���31�8JCOSEKr�EHLN�0hK�5 oDt�jI��jI<1�J�L�Z1�5Zc@y��1MY�qA�HQBTHWMYT�HET09�NK2a3z�/Rn�r@CB4VkCBn�CqPASfa�YR<4gQt�gQ4VSB8t��R?UGTS���Cq��a��P#���Z�C$DUu ��R� �э2�Vӑ��Q�r�f'$NE�+pIs@�$|� �$R�#QA'UPepYg7EBHBALPHEE.b�.bS�E�c�E�c��E.b�F�c�j�FR�V�rhVghd��lV�jV��kV�kV�kV�kV
�kV�iHrh�f�r�m�!�x�kH�kH�kH��kH�kH�iOclORrhO��nO�jO�kUO�kO�kO�kO�kO�FF.bTQ���E���egSPBALAN�CE��RLE�PH_'USP衅F��F|��FPFULC�`3��3��E��1�l��UTO_p �%T13T2t���2NW�� ���ǡ��5�`�擊��T�OU���� I�NSEG��R�REqV��R���DIFH�f�1���F�1�;�COB��;C��2� ��b�4LCHWA�R��;�ABW!��$MECH]Q�@k�,q��AXk�P��8IgU�i�� 
���!ܭ���ROB��CR���ͥ�� �C���_s"T � �x $WEIGHh�9�$cc�� �Ih�.�IF ќ�LAGK�8SK��K�7BIL?�OD��U�&�STŰ�P�; �����������
�Ы�L��  2��`�"�DEBU.�L�&�n��PMMY9���NA#δ9�$D&���$��� Q�   �DOu_�A��� <	� ��~��L�BX�P��N��+�_7�L�t�O�H  �� %"��T���ѼT������TICK/�C�TE1��%������N��c�Ã�R L�S����S�����PROMP�h�E� $I�R� X�~ ���!�MCAI�0��j���_9�C���t�l�R�07COD��FU`�+�ID_" =����耿G_SUFF<0 �3�O����DO��ِ��R��Ǔن�@S����!{������	��H)�_FI��9n��ORDX� �����36��X���Ɩ�GR9�S��ZD�TD�SAVu�ŧ�4 *�L_N�A4���K��DEF_I[�K���g��_����i��Ɠ�š���IS`i �萚����e����4�0i��Dg����D� O|��LOCKEA!�uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ�{� ���}��v�Ա�� g������^���K‒Փ����!w�N�P@'���^���,`�W\�l[R���TEF�Ĩ �OULOOMB_u�0�wVISPITY��A�!OY�A_FR1Id��(�SI��B�R������3��
�W�W��0��09_,�EAS%��@�!�& "���4p�}G;� h ���7ƵCOEFF_AOm���m�/�G!2%�S.�߲CA5�����u�GR` � � $R� �X]�TME�$R�s�XZ�/,)�ER�T;��:䗰�  ]�LLt��S�_SV�&�($~����@�� "SETU��MEA��Z�x0��u������ � �� �� ȰID@�"���!*��&P���$*�F�'����)3��#���"�5;`:*��REC���!=��MSK_���� P	�1_USER��,��4���D�0��VEL,2�0��ȯ2�5S�I��0�M�TN�CFG}1� � ���Oy�N�ORE��3��2�0S�I���� ��\�UaX-�ܑPDE�A� $KEY_�����$JOG<EנSVIA�WC�� 1DSWy���
��CoMULT�GI�@�@C��2� 4 ��#t�+�z�XYZ���쑡���z� �@_7ERR��� ��S L�-���@��s0BB_$BUF-@X1�����MOR�� H	�CU�A3�z�1Q��
��3���I$��FV��2S�bG�� � �$SI�@ G�0VOx B`נOBJE&��!FADJU�#EEGLAY' ���SD�W�OU�мE1PY���=0QT i�0�W�DIR$ba�pےʠDYNբHe	T�@��R�^�X����OPWORK}1��,�SYSB9U@p 1SOP�aR$�!�jU�k�PR��2�ePA�0�!�cu� 1+OP��UJ��a'�zD�QIMAG�A1	��`i�IMACr�IN,�bsRGO�VRD=a�b�0�aP �`sʠ� �^uz��LP�B�@��!PMGC_E,�Q��N@�M�rǱ��1Ų��=q�SL&�~0���$OVSL\G*E��"*E2y�Ȑ�_=p�w ��>p�s���s	�����y���=q�#}1� �@�@;���O/�RI#A��
N��X�s�f�Q�{��PL}1�,RyTv�m�ATUSRBTRC_T(qR��B �����$ �Ʊ��,�~0� D��`-CSALl`�SA���]1gqXE���%���bC��J�
���UP(4����PX��؆�q��y3�w� �PG�5�� $SU�B������t�JMPWAITO��s���LOyCFt�!D=�CCVF	ь�y���R`��0��CC_CTR��Q�	�IGNR_{PLt�DBTBm�P��z�BW)����0�U@���IG�a��I�y�TNLN��Z�R]aK� N��B�0�P�E�s���r��f�SP]D}1� L	�A�`0gఠ�S��UN�{�传]�R!�BDLY��2���sRPH_P�K�E��2RETRIEt��2�b6����;FI�B� �����8� 2��0DB�GLV�LOGS�IZ$C�KTؑUdy#u�D7�_�_T1@�EM�@C\1A��ℽR��D�FCHE3CKK�R�P�0��e��@&�(bLEc�" PA9�T���P�C�߰PN�����A�Rh�0���Ӯ�PO��BORMATT naF�f1h���2�S�F�UXy`	��LBо�4�  rEIgTCH��8PL)��AL_ � $H��XPB�q� C,2�D�!��+2�J3D��� T�pPDC�Kyp��oC� _AL3PH���BEWQo����� ��I�wp �� �b@PAYgLOA��m�_1t�y2t���J3AR���؀դ֏�laTIA�4��5��6,2MOMCP�����������0BϐAD������.��PUBk`R��;����;��Ғ�z4�` I$PI\Ds�o�@�1yՕ�w�2�w�Z��I��I��I���p� ���n���y�e`��9S)bT�SPEED� G��(�Е��/��� Е�`/�e�>��M�<�ЕSAMP�6V0��/���ЕMO�@ 2@�A��QP���C�� n�����������LRf`�kb�ІE9h�EIN 09��7S.В9
�yPy�GAMM�%S���D$GE�T)bP�cD]��2
��IB�q�I�G$HI(0;A��LR�EXPA8)LWVM8z)���g���C5�CHKhKp]�0�I_�� h`eT��n�q���eT,���� ��$�� 1�iPI>� RCH_D�313\��30LE�1�1\��o(Y�7 �t�MSW�FL �M��SCRc�7�@�&��%n�f�;SV���PB``�'�!�B�sS_SAaV&0ct5B3NO]�C\�C2^�0�mߗ� uٍa��u���u:e;��1���8��D�P��� ������)��b9� �e�GE�3��V���}Ml�� � ��YL��QNQS RlbfqXG�P�RR#@dCQp� �S:AW70��B�B[�CgR:AMxP�KCL�H���W�r��(1n�g�M�!o��� �F�P@}t$W P�u�P r��P5�R <�RC�R��%�6�`���� ��qsr X��O�D�qZ�Ug�ڐ>D�[ ��OM#w� J?\?n?�?�?��9�b"��L]�_��� | ��X0��bf��qf�� q`�ڏgzf��Eڐ��>j�"�ܰ��FdPnB��PM�QU��� � 8L�QCsOU!5�QTHI�sHOQBpHYSY�3ES��qUE�`�"��O���  �P��@\�UN���Crf�O�� P���Vu��!����OGR)AƁcB2�O�tVu�ITe �q:pINF�O�����{�qcB�ve�OI�r� (�@SLEQS��q��p�vgqS���� =4L�ENABDRZ�PTIONt�����Q���)�GCF�ЎG�$J�q^r��� R���U�g����rS_ED����ѓ �F��PK���E'NU߇وA�UT$1܅COPY������n�00MNx���PRUT8R� �Nx�OU���$G[rf�5BRGAkDJ���*�X_:@�բ$�����P��W��P��} ��)�}�[EX�YCDR|��NS.��F@r�LG�O�#�NYQ_FREQR�W� �#�h�TsLAe#������ �CRE� s��IF��sNA���%a�_Ge#STA�TUI`e#MAIL�����q t��������ELEM��� �/0<�FEASI?�B��n�ڢ�1�]� � I�p��`Y!q]�t#A�ABM����E�p<�VΡY�BCASR�Z��S�UZ��0$q���RMS_TR;�qb  ���SY�	�ǡ��$����>C�Q`	� 2� _�TM�� ����̲�@ �A��)ǜ��i$DOU�s]$NLj���PR+@3���r�GRID�qM�BA�RS �TY@��O�TO�p��� Hp_"}�!����d�O�P/��� � �p�`P�OR�s��}���SReV��)����DI&0T����� #�	�#�U4!�5!�6!�7!�I8�e�F�2��Ep?$VALUt��%���ֱ��/��� !;�1�q�����(F_�AN�#�ғ�Rɀ|(���TOTAL��,S��PW�Il��REGEN�1�c�X��ks(��a���`T1R��R��_S� ��1ଃV�����⹂Z�E��p�q��Vr���7V_H��DA�S�����S_Y,1�R4�S�� AR�P2� >^�IG_SE	s��d��å_Zp��C_��~��ENHANC�a�� T ;�8������INT�.���@FPsİ_OVRsP�`p�`��Lv�҂o��7�}��Z�@�SSLG�AA�~�2 5�	��D��S�BĤ�DE�U�����T�E�P���� !�Y��
�J��$2�IL_MC�x r#_��`TQ�`��q���'�B5V�C�P_� 0ڽM�	V1�
V1��2�2�3�3
�4�4�
�!���`� � m�A�2IN~VIBP���1�U2�2�3�3�4�4�A@-�C2�p� MC_YFp+0�0L	1(1d���M50Id�%"FE� S`�R/�@�KEEP_HNA�DD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0�#i�.�#REM�"�$�P�½%�!�(U}�e�$�HPWD  �`#SBMSK|)G��qU2:�P	�COLLAB� �!K5��B�� ��g��pI�TI1{9p#>D� �,�@FLAP��$�SYN �<M�`C�6���UP_DL�YAA�ErDELAh�0ᐢY�`AD�Q�4BQSKIP=E�� ���XpOfPNTv�A�0P_Xp�rG �p�RU@,G��:I+�:I B1:IG�9JT�9Ja�9J�n�9J{�9J9<��R=A=s� X����4�%1�QB� NFL#IC�s�@J�U�H�LwNO_H�0�"?�֌RITg��@_P�A�pG�Q� ���^�U��W��LV�>d�NGRLT�0_q���O�  " ��OS��T�_JvA V	�APPR_WEIGH�s�J4CH?pvTOR8��vT��LOO��]�D+�tVJ�е�ғA�Q�U�S�XOB'�'�{�SJ2P���7�X�T�<a43DP=`Ԡ\"p<a�q\!��RDC�ѮL� �рR��R�`� �RV��jr�b�RGE��*��cNFLG�a�Z���SsPC�s�UM_<`>^2TH2NH��P~.a 1� m`�EF11��� �lQ �!#� <�p3AT� g�S�&�Vr�p�t�Mq�Lr���HO�MEwr�t2'r�-?Qcu��w3'r������
�w4'r�'�9�K�]�(o����w5'r뤏���ȏڏ����w6'r�!�3�E�W�i�{��w7'r힟��ԟ���
�w8'r��-�?�Q�Hc�u��uS$0�q�p�� sF��`)a�"`P�����`/���&-�IO[M�I֠���)�POWE��# ��0Za*���� �5��$DS=B GNAL���0�Cp��m`S232N3�� �~`��� �/ ICEQP��PE�p��5PIT����O�PBx0��FLOW�@TRvP��!U����CU�M��UXT��A��w�ERFAC��� U��ȳC�H��� tQ  _���>�Q$����O)M��A�`T�P#�UPD7 A�ct�T��UEX@�ȟ�U �EFA: X"�1RS9PT�����T ���PPA�0o񩩕`EXP�IOS���)Ԃ��_���%��C�WR�A��ѩD�ag֕`~ԦFRIENDsa�C2UF7P����TO;OL��MYH C2�LENGTH_V�TE��I��Ӆ�$SE����UFI�NV_���RsGI�{QITI5Bb��Xv��-�G2-�G17�w�SG�X��_��UQQD=#���AS��d~C�`��qᾭ� �$$C/�S�`�����S0)`|����VERSI� ���)`�5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����S0����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT��C��  ��DI�N�O�A�Dq�EXE��HPV_��AT�Qz
��LARM�RECOV ��RgLMDG �*�5�OLM?_IF *��`d�O�_�_�_�_j�_�'o9oKo]onm, 
��odb��o�o�o0�o^��$� z, �A   2D{�P�PINFO u[ �Vw��������`����� ��*��&�`�J���n�����DQ���� 
��.�@�R�d�v���𚟬���a
PPLI7CAT��?�P���`Ha�ndlingTo�ol 
� 
V�8.30P/40�Cpɔ_LI
8�83��ɕ$ME�
F0G�4�-?
398�ɘ��%�z�
7�DC3�ɜ
�No+neɘVr���ɞ_@6d� ~Vq_ACTIVU���C죴�MOD�P���C�I��HGA�PON���O�UP�1*�� Ai�m����Қ_��6��1*�  �@��������Q����Կ�@�
���=�� ���5��Hʵl�K�HTTHKY_��/�M� SϹ���������%� 7ߑ�[�m�ߝߣߵ� ���������!�3�� W�i�{�������� ������/���S�e� w��������������� +�Oas� ������ '�K]o��� �����/#/}/ G/Y/k/�/�/�/�/�/ �/�/�/??y?C?U? g?�?�?�?�?�?�?�? �?	OOuO?OQOcO�O �O�O�O�O�O�O�O_ _q_;_M___}_�_�_��_�_�_�_kŭ�TO�p��
�DO_CL�EAN9��pcNM  !{衮o�o��o�o�o��DSP�DRYRwo��HI��m@�or��� ������&�8�J���MAXݐWdak�H�h�XWd�d��>�PLUGGW�Xg\d��PRC)pB�`E�kaS�Oǂ�2DtSEGF0�K � �+��o�or�����p�����%�LAPO b�x�� �2�D�V�h� z�������¯ԯ�+�TOTAL����+�_USENUO�\�� e�A�k­�RGD�ISPMMC.�2��C6�z�@@Dr\��OMpo�:�X�_S�TRING 1	~(�
�M!��S�
��_ITwEM1Ƕ  n� �����+�=�O�a� sυϗϩϻ����������'�9�I/�O SIGNAL���Tryou�t Modeȵ�Inpy�Simu�lateḏO�ut��OVE�RRLp = 10�0˲In cy�cl�̱Pro?g Abor��̱�u�Status�ʳ	Heartb�eatƷMH �Faul	��Aler�L�:�L�^�p����������� ScûSaտ��-�?� Q�c�u����������� ����);M_q��WOR.�û� �����+ =Oas��������//'.PO����M �6/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�?8�?�?H"DEVP.�0 d/�?O*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8_J_\_n_PALT	��Q�o_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o8�o�_GRIm�û 9q�_as��� ������'�9� K�]�o�������'�R	�݁Q����)� ;�M�_�q��������� ˟ݟ���%�7�I�ˏPREG�^���� [�����ͯ߯��� '�9�K�]�o�������෿ɿۿ�O��$A�RG_� D ?	����0���  	]$O�	[D�]D���O�e�#�SBN_�CONFIG �
0˃���}�C�II_SAVE � O�����#�T�CELLSETU�P 0�%  ?OME_IOO�O�%MOV_H������REP��J��UTOBACK�����FRwA:\o� Q�,o���'`��o������ �� f�o�����*�!�3�`�Ԉ��f��� ��������o�{��&� 8�J�\�n�������� ����������"4F Xj|����p��끁  ���SYSUIF.S�V V T<pVD� MP 6.:G/IF PHD_8q��N�t#�®f�INI�Po����c�MESSA�G�����8��OD�E_D����z��Ox�0�c�PAUSM!�!�0� (q73�U/g+(Od/ �/x/�/�/�/�/�/�/ ???P?>?t?1�0$~: TSK  @-x��T�f�UPDT��d�0
&XWZD_ENB����6�STA�0��5"�X�IS��UNT 2�0Ž� � 	� ��z���eng��-뷛�#S�o�U@��H��A��tL�Oo�}Cw쀕g�^����.��O�O�O�O/_2FME�T߀2CMPTAA���@�$A�-�@���@���@���]�5��5�(d�5��P5�r��5F*5�33�8]SCRDCFG� 1�6�Ь�Ź�_�_o@o(o:oLo��o�Q�� �_�o�o�o�o�o�o]o �o>Pbt��0�o9�i�GR<@M|/�sUP_NA��/�	i��v_E�D�1�Y� 
� �%-BCK�EDT-�'�G?ETDATAU�o��9�u?�j�H�o��f�\��A��  ���2�&�!�E���:�Q���~�ŏ׏m����3��&۔�� D��ߟJ�����9�ǟ�4���ϯ�(���@�]�o�����5N� �����(�w��)�;�ѿ_��6ϊ�gϮ� (�CϮ���ϝ�+��7��V�3�z�(��z� ����i����8��&���~�)���F�ߟ�5����9~������)����Y�k�����CR�!ߖ���W� q���#�5���Y��p$�?NO_DEL��r�GE_UNUSE���tIGALLO�W 1��(�**TEM*�S	$SERV�_GR�V� : REG�$�\� �NUM�
��P�MUB ULA�YNP\PM�PAL�CYC10#6 $\ULSU�8:!�Lr�BOX�ORI�CUR_���PMCNV6�10L�T4DLI�0��	����BN/`/r/�/��/�/�/�/���pLA�L_OUT ��;���qWD_AB�OR=f�q;0IT_R_RTN�7�o	�;0NONS�0�6� 
HCCFS_U?TIL #<�5�CC_@6A 2#; h ?�?�?O�#O6]CE_OPT;IOc8qF@�RIA_Ic f5�Y@�2�0F�Q�=2q&}�A_LI�M�2.� ���P�]B��KXʊP
�P�2O�Q�R�B�r�qF�PQ 5T1)TR�H�_:J�F_PARAMGoP 1�<g^�&S�_�_�_�_�VC��  C�d�`��o!o`�`�`�
`�Cd��Tii:ah:e>eBa�GgC�`~� D� D	�`m�w?��2HE �ONFI� E?�aG�_P�1#; ���o1C�Ugy�aKPAU�S�1�yC ,�������� �	�C�-�g�Q�w���@������я���rO�A��O�H�LLECT_�B�IPV6��EN. QF�3�ND�E>� �G�7�1234567890��sB�TR�����%
 H�/%) �������W���0� B���f�x���㯮��� ү+�����s�>�P� b����������ο� �K��(�:ϓ�^�|�:�B!F� �I|�IO #��<U%�e6�'�9�K���T-R�P2$��(9X�t�Y޼`%�̓ڥH���_MOR�3&��=��@XB� �a��A�$��H�6� l�~���~S��'�=�r�_A?�a�a`��@K(��R�dP��)F�ha�-�_�'�9�%
�k��G� ��%yZ�%��`�@]c.�PDB��+����cpmidbag��	�`:��@�QF��p��N ' ���+
���]ܭ@2s<�V^��@+sg�,$� 5sfl��q��ud1:��:J��DEF �*ۈ��)�c��buf.txt�����_L64?FIX ,���� ��l/[Y/�/}/�/�/ �/�/
?�/.?@??d? v?U?�?�?�?�?�?�?|,/>#_E -���<2ODOVOhOzO�OV6&IM��.o�YU�>���d�
�IMMC��2/����dU,�C��20�M�QT:U>w�Cz  B�i��A���A����Au�gB3�*�CG�B<�=�w�i�B.��B����B��5B��$�D�%B����ezVC�q�C��v�D���D�-lE\D�n�j���29"��22o�D|������ ���C�ZC����
�xObfi�D4cdv`D��`�/�`v`s]E�D �D�` E4��F*� Ec���FC��u[F����E��fE��f�Fކ3FY��F�P3�Z��@��33 ;��>LS���Aw�n,a@��@e�5Y���a����`A��w�=�`<#����
��?�ozJR�SMOFST �(�,bIT1��D2 @3��
д����a���;��bw?���<�M�N/TEST�1O�CER@�4��>VC5`#A�w�Ia+a�aOR�I`CTPB�U�C��`4���r��:d�����qI?�5���qT_�PROG ��
�%$/ˏ�t���NUSER  �U������KEY_TBL  �����#a��	
��� !"#$%&�'()*+,-.�/��:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s������LCK�x
����STAT/���s_AUTO_D�O(	�c�IND�T_ENBP���R�pqn�`�T2����ScTOr`���XC��� 26���8
�SONY XC-�56�"b����@���F( А=�HR50w����>�P�7b�t�Af!f����ֿ� Ŀ� ���C�U�0�yϋ�f� ���Ϝ��������-���TRL��LET�E(��T_SCREEN �ڟkcs���U��MMENU 1=7�� <ܹ� ��w��������� K�"�4��X�j��� ����������5��� k�B�T�z��������� ������.g> P�t����� �Q(:�^ p����/�� ;//$/J/�/Z/l/�/ �/�/�/�/�/�/7??  ?m?D?V?�?z?�?�? �?�?�?!O�?
OWO.O @OfO�OvO�O�O(y��?REG 8�y�����`�M�ߎ�_M�ANUAL�k�DwBCO��RIGY��9�DBG_ERRML��9�ۉq�ر_�_�_ ^QNU�MLI�pϡ�pd�
�
^QPXWOR/K 1:���_5o�GoYoko}oӍDBT;B_N� ;������ADB__AWAYfS�q/GCP 
�=�p�f�_AL�pR��bbRY��[�
�WX_�P 1<{y�n�,�%oc��P��h_M��I�SO��k@L��sON�TIMX��
�ɼ�vy
��2sMO�TNEND�1tR�ECORD 1B΋� ���sG�O�]�K��{�b���� ����V�Ǐ�]���� 6�H�Z��������� #�؟������2��� V�şz��������ԯ C���g��.�@�R��� v�寚�	���п��� c�χ�#ϫ�`�rτ� ��Ϻ�)ϳ�M��� &�8ߧ�\�G�Uߒ��8�������K� �p����6��%RC7� n���ߤ������A�4���$���H�03�A�~��;��� ����9���]������|�B#Zl���zTOLEREN\��rB�'r�`L���^PCSS_CCS�CB 3C>y�` IP��}�~�< �_`r�K�����/�{��5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O_�~ֽLL� D���&qET�c�a C[C��PZP^r_W A� p� �s�p��QGPt[	 !A�p�Q�_�[? �_h�[oU�p�P�pSB�V�c�(a@�PWoio{h+�o�Xa�o�oY��[�	r�hLW��N:�p����}6ګ�c���aD@VB���|�G����+��K� A�otGhXGr�S�o����eB  _ =��Ͷa>�t&YB�� �pC�p�q
�aA"�H�S�Q-��q ���ud�v�����Af�P ` 0����D^P��p@�a
�QXTHQ����a� aW>� �a9P� �b�e:�L�^�h�Hc�́PQ�RFQ�PU�z �֟�o\^��-�?���c�u����zCz�ů�b2�Щ�R�D�����l)* ����S̡0��]�0� .��@���EQ�p�� F�X�ѿUҁп�VS�ȺNSTCY S1E��]�ڿ ��K�]�oρϓϥϷ� ���������#�5�G��Y�k�}ߏߒ��DEVICE 1F5� MZ�۶a��	�@ ��?�6�c���	{�𰟗��_HNDGD G5�VP���R>�LS 2H�ݠ� �/�A�S�e�w������ ZPARAM �I�FgHe�RBoT 2K��8р�<��WPpC�C�,`¢P�Z�z��*%{�C��2�j�MTLU,`"nPB , s��M� }�gT�g��
B��!�bcy�[2Dch z����/���/gT#I%D��CǓ` b!�R��A���A,��Bd���A�;���_C14kP�!2�C��$Ɓ��]�ffA�À���B�� �| �0��/�/�T (��5 4a5�}%/7/d?/ M?_?q?�?�?�?�?�? O�?OO%O7OIO�O mOO�O�O�O�O�O�O �OJ_!_3_�_�_3�_ �_�_�_�_o�_(oo Lo^oЁ=?k_IoS_�o �o�o�o�o�o�o #5G�k}�� �����H��1� ~�U�g�y�ƏAo�Տ ���2�D�/�h�S��� go����ԟ����ϟ� ��R�)�;���_�q� ���������ݯ�<� �%�7�I�[�m����� ����}�&��J�5� n�YϒϤϏ��ϣ�ѿ ������F��/�A� ��e�w��ߛ߭����� ����B��+�x�O�a� �����������,� ��%�b�M���q����� ����������L #5�Yk}�� � ��61 CUg����� ���	//h/���/ w/�/�/�/�/�/
?�/ .?@?I/[/1/_?q? �?�?�?�?�?�?�?O O%OrOIO[O�OO�O �O�O�O�O&_�O_\_ 3_E_W_�_?�_�_�_ �_�_"ooFo1ojoE? s_�_�om_�o�o�o�o �o0f=Oa �������� ��b�9�K���o��� Ώ��[o��(��L��7�I���m������$�DCSS_SLA�VE L��}�ё���_4D  љ�~�CFG Mѕ���������FRA:\ĐL�-�%04d.CS�V��  }�� ����A i�CHq�z������|�����"������Ρޯ̩硞Ґ-��*����_�CRC_OUT �N������_�FSI ?њ ����k�}� ������ſ׿ ���� �H�C�U�gϐϋϝ� ���������� ��-� ?�h�c�u߇߽߰߫� ��������@�;�M� _����������� ����%�7�`�[�m� ��������������� 83EW�{� ����� /XSew��� ����/0/+/=/ O/x/s/�/�/�/�/�/ �/???'?P?K?]? o?�?�?�?�?�?�?�? �?(O#O5OGOpOkO}O �O�O�O�O�O _�O_ _H_C_U_g_�_�_�_ �_�_�_�_�_ oo-o ?ohocouo�o�o�o�o �o�o�o@;M _������� ���%�7�`�[�m� �������Ǐ����� �8�3�E�W���{��� ��ȟß՟���� /�X�S�e�w������� �������0�+�=� O�x�s���������Ϳ ߿���'�P�K�]� oϘϓϥϷ������� ��(�#�5�G�p�k�}� �߸߳����� ���� �H�C�U�g���� ���������� ��-� ?�h�c�u��������� ������@;M _������� �%7`[m ������� /8/3/E/W/�/{/�/ �/�/�/�/�/??? /?X?S?e?w?�?�?�? �?�?�?�?O0O+O=O OOxOsO�O�O�O�O�C��$DCS_C_�FSO ?�����A P �O�O_?_ :_L_^_�_�_�_�_�_ �_�_�_oo$o6o_o Zolo~o�o�o�o�o�o �o�o72DV z������� 
��.�W�R�d�v��� ����������/� *�<�N�w�r������� ��̟ޟ���&�O� J�\�n���������߯ گ���'�"�4�F�o� j�|�������Ŀֿ�������G�B�T��OC/_RPI�N_j� �����ς��O����1�XZ�U��NSL��@&� h߱���������"�� /�A�j�e�w���� ����������B�=� O�a������������� ����'9b] o������� �:5GY�} ������// /1/Z/U/g/y/�/�/ �/�/�/�/�/	?2?-? ??Q?z?u?��ߤ߆? �?�?�?OO@O;OMO _O�O�O�O�O�O�O�O �O__%_7_`_[_m_ _�_�_�_�_�_�_�_ o8o3oEoWo�o{o�o �o�o�o�o�o /XSew��� �����0�+�=� O�x�s���������͏ ߏ���'�P�K�]��o����� �PRE_?CHK P۫��A ��,8��2��� 	 18�9�K���+�q� ��a�������ݯ�ͯ �%��I�[�9���� o���ǿ��׿���)� 3�E��i�{�Yϟϱ� ������������-� S�1�c߉�g�y߿��� �����!�+�=���a� s�Q�������� ������K�]�;��� ��q������������� #5�Ak{� ����� CU3y�i�� ����/-/G/ c/u/S/�/�/�/�/�/ �/??�/;?M?+?q? �?a?�?�?�?�?�?�? �?%O?/Q/[OmOO�O �O�O�O�O�O�O_�O 3_E_#_U_{_Y_�_�_ �_�_�_�_�_o/oo SoeoGO�o�o=o�o�o �o�o�o=- s�c����� ��'��K�]�woi� ��5���ɏ������� �5�G�%�k�}�[��� ����ן�ǟ���� C�U�o�A�����{��� ӯ����	��-�?�� c�u�S�������Ͽ� ������'�M�+�=� �ϕ�w�����m���� ��%�7��[�m�K�}� �߁߳��߷����!� ��E�W�5�{��ϱ� ��e�������	�/�� ?�e�C�U��������� ������=O- s����]�� ��'9]oM �������/ �5/G/%/k/}/[/�/ �/��/�/�/�/?1? ?U?g?E?�?�?{?�? �?�?�?	O�?O?OO OOuOSOeO�O�O�/�O �O�O_)__M___=_ �_�_s_�_�_�_�_o �_�_7oIo'omoo]o �o�o�O�o�o�o! �o1W5g�k} ������/�A� �e�w�U�������я ��o����	�O�a� ?�����u���͟��� ��'�9��]�o�M� ��������ۯ��ǯ� #�ůG�Y�7�}���m� ��ſ�����ٿ�1� �A�g�E�wϝ�{ύ� ������	�߽�?�Q� /�u߇�e߽߫ߛ��� �����)���_�q� O���������� ���7�I���Y��]� ��������������! 3WiG��} ����%�A �1w�g��� ���/+/	/O/a/ ?/�/�/u/�/�/�/�/ ?�/9?K?�/o?�? _?�?�?�?�?�?�?O #OOGOYO7OiO�OmO �O�O�O�O�O_�O1_ C_%?g_y__�_�_�_ �_�_�_�_o�_+oQo /oAo�o�owo�o�o�o �o�o);U__q ������� �%��I�[�9���� o���Ǐ�����ۏ!� 3�M?�i��Y����� ��՟�ş����A� S�1�w���g�����������ӯ�+�=��$�DCS_SGN �QK�c��7m�� 16-M�AY-19 10?:20   O�l��4-JANt�08�:38}�����? N.DѤ�����������M4�o���Im��P��Z�q��  O�V�ERSION �[�V3.5�.13�EFLO�GIC 1RK���  	���P�?�P�N�!��PROG_ENB  ��6Ù�o�ULSE  T����!�_ACCL{IM���������WRSTJN�T��c��K�EM�Ox̘��� ���INIT S.�G�Z����OPT_SL �?	,��
 	�R575��Y�7�4^�6_�7_�50
��1��2_�@ȭ��><�TO  Hݷ�t��V�DEX���dc����PAT�H A[�A\��g�y��HCP_�CLNTID ?<��6� @ȸ�����IAG_GR�P 2XK�? ,`��� � �9�$�]�H������123456�7890����S�� |�������!�� ��H���;� dC�S���6� ����.�R v�f��H� �//�</N/�"/ p/�/t/�/�/V/h/�/ ?&??J?\?�/l?B? �?�?�?�?�?v?O�? 4OFO$OjO|OOE� �Oy��O�O_�O2_��@_T_y_d_�_,
�B^ 4�_�_~_`Oo �O&oLo^oI��Tjo�o .o�o�o�o�o �O' �_K6H�l�� �����#��G� 2�k�V���B]���Ǐ ُ�������(��L��B\Drx�@���PC����4 � 79֐�$��>���:�����ߟʟ�ܟ���CT_CONFIG Y���Ӛ�eg�U���STBF_TTS��
��b�����t��u�O�MAU���|��MSW_CF�6�Z��  �O�CVIEW��[ɭ������-�?� Q�c�u�G�	�����¿ Կ������.�@�R� d�v�ϚϬϾ����� ��ߕ�*�<�N�`�r� ��ߨߺ�������� ��&�8�J�\�n��� !�������������4�F�X�j�|����R%C£\�e��!*�B^ ������C2g�{�SBL_FAULT ]��ި�GPMSKk��*��TDIAG ^�:�աI��U�D1: 6789?012345�G�BSP�-?Qc u��������//)/;/M/� ��
@q��/$�TORECP��

� �/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOi/{/xO��/UMP_OPT�IONk���ATR�¢l��	�EPME�j��OY_TEMP�  È�3B��J�P�AP�DU�NI��m�Q��YN_BRK _ɩ��EMGDI_S�TA"U�aQK�XPN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 J�#�%�,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;��A����O ���� � I ߵ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����⣆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7���; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  D�C����(7�?�<B�?B����2�ٸ*9�N SMTT#t�[)��X}�C�f�HoOSTCd1ux����?�� M5Cx��;zOx�  27.0�@=1�O  e�O�O 	__-_;Z�O^_p_�_�_�LN_HS	ano?nymous�_�_�_oo1o yO��FhFk�O�_�o�O�o�o �o�oJ_'9K] �o�_����� 4o�XojoG�~�o^� ������ŏ���� �1�T���y����� ������,�>�@�-� t�Q�c�u��������� ϯ���(�^��M� _�q�����ܟ� �ݿ ��H�%�7�I�[Ϣ� ϑϣϵ����l�2� �!�3�E�Wߞ���¿ Կ����
������� /�v�S�e�w���� ���������+�r� �ߖ�s�����߻��� �������'9K] ��������� 4�F�X�j�l>��} ������/ /1/T��y/�/�/�/�/.D\AENT {1v
; P!J/.?  ��/3? "?W??{?>?�?b?�? �?�?�?�?O�?AOO eO(O�OLO^O�O�O�O �O_�O+_�O _a_$_ �_H_�_l_�_�_�_o �_'o�_Koooo2o{o Vo�o�o�o�o�o�o 5�oY.�R��v��zQUIC�C0���3��t1 4��"����t2��`��r�ӏ!ROUT�ERԏ��#�!�PCJOG$����!192.16?8.0.10��s?CAMPRTt�P��!d�1m�����R�T폟�����$NA�ME !�*!�ROBO���S_�CFG 1u�)� �Au�to-start{edFTP&��=?/֯s��� �0�B��f�x����� ����S������,� ��������ϼ�ޯ�� �������ʿ'�9�K� ]�oߒ�ߥ߷�����p����SM% y�{�U�ό����� �����
��.�@�c���v������������z�%�7�I�K�8� \n���k��� ��3�FXj |����a��7/M*/</N/ `/r/9�/�/�/�/� �/�/?&?8?J?\?� m?���?�//�?�? O"O4O�/XOjO|O�O �O�?EO�O�O�O__ 0_w?�?�?�?�O�_�? �_�_�_�_o�O,o>o Poboto�_o�o�o�o �o�oK_]_o_L�o �_�o�����o�  ��$�6�Y�Y�~��������ƏZ�_ER�R w3�я�P�DUSIZ  jg�^�p���>�?WRD ?r�Cq��  guestb�Q�c�u��������`�SCDMNGRP 2xr�w���H��g�\�b�K� 	�P01.00 8~`�   � ��   B � ��� ����H���L���L��L�����O�8�����l�����a�4�  �Ȥ� �V8���\���)�5`�;��������d�.�@�R�ɛ_�GROUېy������	ӑ���Q?UPD  ?u��Y��İTYg�����TTP_AU�TH 1z�� �<!iPend�an��-�l����!KAREL:q*-�6�H�KC]��m��U�VISI?ON SET������!�����R�0� �H�Bߏ�f�x��ߜ������CTRL �{����g�
��FFF9E3���AtFRS:DE�FAULT;��FANUC We�b Server ;�)����9�K��ܭ�����������߄WR�_CONFIG ;|ߛ ;���IDL_CPU_kPCZ�g�B�I��y� BH_�MIN�j�)�}�GNR_I�O��g���a�NPT_SIM_D_������STAL_oSCRN�� ����TPMODNTOqL������RTY��0y���� �ENO����Ѳ]�OLNK 1}��M��������eMAS�TE��ɾeSLAVE ~��c�O_CFGٱB�UO�O@CYC�LEn>T�_AS�G 1ߗ+�
 ����//+/ =/O/a/s/�/�/�/�/\��NUM��=
@IPCH�^RTRY_CNZ�����@������b�� @kI�+�E�z?E�a�P_ME�MBERS 2��ߙ� $���2����ݰ7�?�9a�SD�T_ISOLC � ����$J2/3_DSM+�3JOBPROCNn��JOG��1�+��d8�#?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSR�EQO��KANJI�_���a[�MO�N ����b�y N_goyo�o�o�o�Y�`3�<� ��e�_ִ���_L���"?`EYLOGGINL�E�������$�LANGUAGE� ��<T� ,{q�LGa2�	�b�마g�xP��  U��g�'���b���>�MC�:\RSCH\0�0\<�XpN_DISP �+G�H�8�O�O߃LOCp��Dz���AsOGBOOK �������󑧱����X �����Ϗ����0a�*��	p������!�m��!���=p_BUFF 1�p��2F幟����՟D� Coll�aborativ ǖ���F�=�O�a�s� ������֯ͯ߯����B�9�K���DCS� �z� =���'�f��?ɿۿ���|H@{�IO 1��G ~?9Ø��9� I�[�mρϑϣϵ��� �������!�3�E�Y� i�{ߍߡ߱�������Z�E��TMNd�_ B�T�f�x������ ��������,�>�P��b�t�������L��S�EVD0��TYPN1�$6����QRS"0&��<2F�L 1�"�J0� �������FGTP:pOF�NGNAM1D�mrn�tUPS�GI"5��aO5�_LOA�DN@G %�%�DF_MOTN��y�� MAXUALRM�'���(��'_PR"4F0d��1��B_PNP� V� 2�C	M�DR0771ߕz�BL"8063%�@ �_#?�ߒ|/�C��z�6��/􈃟/Po@P 2���+ �ɖ	~T 	t  ��/ �%W?B?{?�k?�? g?�?�?�?O�?*OO NO`OCO�OoO�O�O�O �O�O_�O&_8__\_ G_�_�_u_�_�_�_�_ �_o�_4ooXojoMo �oyo�o�o�o�o�o �o0B%fQ�u �������� >�)�b�M�����{��� �����Տ��:�%��^�p�S�������D�_LDXDISA�pB�MEMO_{APjE ?C
 �,�(�:��L�^�p������IS�C 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%A �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A�z�4��~�K��������K:z�j]�Q_D��^��PL_NAME �!3%,�!�Default �Personal�ity (fro�m FD) �R�R2� 1�L?6(L?�,0	l d���� ����//(/:/ L/^/p/�/�/�/�/�/�/�/ZX2u?0?B? T?f?x?�?�?�?�?\R<?�?�?O O2ODO�VOhOzO�O�O�OZZK`\R�?�N
�O_\TP�O:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHo_)_~o�o �o�o�o�o�o�o  2DVhz�[omo ����
��.�@� R�d�v���������Џ�� Ef  Fb� F7���   ��!��d��@�R�6�t��� ���l���ʝ����� ݘ���� "�@�F�d���� "�|��ݐA�  ϩ�U[�$n�B��E ��� � @D�  &�?�� �?�@��A@�;f��FH�� ;�	l,�	 '|��j�s�d�/>��� ��� �K(��Kd$2�K ��J7w��KYJ˷�ϜJ�	�ܿ�� @�I���_f�@w�z��f򿿾γ�N�������	Xl�����_��S�ĽÔ�}�I ����5�?��  ����A�?oi#�;����� ���l� �Ϫ�-���ܛ�G�G�Ѳ��@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=�����в@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj��a�Be�Ci��#��Bи�ee^��^^ȹBР ��P����̠�����ADz՟�n�3��C��i�@�R�R�Y���� { �@� ���x�����?�ff������n� ɠ#�ѱy9G
(���I�(�@uP~����t�t����>����;�Cd�;��.<߈�<�g�<F+�<L�������,�d��,�̠?fff?��?&&��@���@x��@�N��@���@T��H�ِ�!-�ȹ� |��
`����� ��//</'/`/r/0]/�/��eF���/ �/�/�/m?��/J?��(E��G�#�� FY�T?�?P?�? �?�?�?�?O�?/OO ?OeOk���O�IQOG� ?�O1?�OmO_0_B_DT_������A_��_	_�_�_�_ o��A���An0 bФ/o C��_Uo�_�Op���`�o�o�o�o���W������oC�E�A q�H�d��؜a�@q��e�F�BµW�B]�NB2�(�A��@�u\�?�D��������b�0�|�uR�����
x~��ؽ��Bu�*C��$�)`��$ ���G�C#���r�AU����1��eG�D�I�m�H�� I:��I�6[F����C�I���J�:\IT��H
~QF�y���p�*J�/� I8Y�I��?KFjʻCe�o ��s�����Џ���ߏ �*��N�9�r�]��� ���������۟��� 8�#�\�G�����}��� ��گů���"��� X�C�|�g�����Ŀ�� �����	�B�-�f� Qϊ�uχ��ϫ����� ���,��P�b�M߆� qߪߕ��߹������� (��L�7�p�[��������s($��g�3:����$���3���d�,�4���@�R���㚅l�~�wa����e����wa4 �{ ������(L:JueP�P~�A�O�������	����G2W }h������ /���O�O7/m/[(d=�s/U/�/�/�/�/ �/?�/1??U?C?y?��=  2 Efn9gFb��77�9f�B)aa)`C9A`�&`w`@-o�?w`e�O )O�?MO�Ow`�?�? �O�O�O�O9c?�0�A*7ht4w`w`!uw`xn
 �O 9_K_]_o_�_�_�_�_ �_�_�_�_o#ozzQ� ��h��G����$MR_CAB�LE 2�h� �a�T� @@�0�Ae��a�a�aK��`��0�`C�`~�aO8�tB�n��d��`�aE?�4�E�#�oZ�f�#��0��0>�DO��By`���Š��bE?D4E�c,��o��g8  ���C��07�d4
v���0 �b��XOE�Z&�l�`�y`
qC�p�bHE��
v#g�5D��Q��qz�lҠ`��0��q�p�b0�
v��%c���b=%	E;h��u/o�c-� �4tH�\�?�9�K�]� o�ԏϏ��
�ɏۏ@����?��eo ��a���������b����� �����`�	 ����@�������% �*�0��6 ��ݐ�����`���	����@�������*,� ,�-�\cO�M �ii���3� � ���%% 2345678901i�B{� f����������j�1����
���`�not sGent3�����;��TESTF�ECSALGR # e�qiG�1d.�š-
:�� �DCb�S�Q�c�u��� 9�UD1:\mai�ntenances.xml��ֿq�� =��DEFAULT-���4\bGRP 2��M�  =��a��{p  �%�Force�so�r check ) ���b�z��p����h5-[ �ϻ�������ϖ�D�%!1st� cleanin�g of con�t. v�ilation��}�Rߗ+��[�ߔߦ߸�ݽ�mech�c�al`������0��h5k�@�R��d�v�����(�rol�le_Ƶ�����/���(�:�����Basic quarterly�������,����������M��M��:C@�"GpP�a�b`�4��������#C ���M"��{P�bt���Su�ppq�greas!e���?/�&/8/J/\/��C+ g}e��. batn�!y`/��/h5	/�/��/�/? ?_�ѷe�n'�v��/�/��/���?�?�?�?�?�QG=?O�qp"CrB1O��0�/`OrO�O�O`�O�t$��Lf��C!-m��A�O:�OO$_�6_H_Z_l_�t*cgabl�Om���S!<m��Q�_:�
_�_ �_oo0oo)(Ӂ/�_�_���_�o�o�o�o��o�O@haul1�l�2r xm�<qC:��op�������Repla�W�fUȼ2�:�.�_4�F�X�j�|�m�$ %���o�������#��� 
��.�@���d���ŏ ׏����П����U� *�y�����r������� ��	�q��?�߯c�8� J�\�n���ϯ����� ڿ)����"�4�Fϕ� jϹ�˿��������� ���[�0�ϑ�fߵ� �ߜ߮�����!���E� W�,�{�P�b�t��� �߼�����A��(� :�L�^��������� ����� $s�H ������q���� �9]o�Vh z���U�#� G/./@/R/d/��/ �/��//�/�/?? *?y/N?�/�/�?�/�? �?�?�?�???Oc?u? JO�?nO�O�O�O�O+J�r	 H�O�O__ 6M2_@OBE:_p_>_P_ �_�_�_�_�_ o�_�_ oHoo(oZo�o^opo �o�o�o�o�o �o �:z �bA?� ; @�q _� ��Fw�� �Hw* �** @q >v�p2T�f�x�:���8����ҏ��eO^C 7�Տ#�5�G�	�k�}� ��ُ���c����� W��C�U�g���ß)� ����ӯ���	��-� w�����9�������m�@Ͽ��=�O�E	A��$MR_HIS�T 2�>uN��� 
 \�$Force �sensor c�heck  12�34567890�q�3����ß�߉N}SB� �-319.8 h�ours RUN� 9.�Y�!1s�t cleani�ng of co�nt. ventilation0�P�ϖϨ�-�Y����mech��cal�i�%Ό4��o�oDN�t��95���1����rollAeh�+�=�O��Y��Basic q�uarterly ߒߤ߶�
O4�F�� (�����b�t��� ��������M�_�����:�����p���:�S�KCFMAP  ]>uQ��r�5�������ON�REL  .��3���EXCFEN��:
��Q�FNCXJJOG_OVLIM8dN�\� ��KEY8�=�_PAN7�P���������SFSPDTYP8xC��SIG�:>��T1MOT�G���_CE_GRoP 1�>u\�D�����/� ���/�/U// y/0/n/�/f/�/�/�/ 	?�/???�/c??\? �?P?�?�?�?�?�?O�)OOMO,���QZ_�EDIT5 )T�COM_CFG 1���[�O�O�O� 
�ASI ��y3�
__+[_O_��>O�_bH�T_ARC_U�քT_MN_M�ODE5�	U?AP_CPL�_g�NOCHECK {?�� �� o.o@oRodovo�o �o�o�o�o�o�o�*!NO_WAI�T_L4~GiNTƑA���EUwT_7ERRs2���3���ƱJ�����X>_)��|MO�s��}�x:Ov���8�?����� l��r_PARAM�r�����j���5�<5�G� =  r�b� t�s�X�������������֟�0�����b�t�����SUM_?RSPACE������Aѯۤ�$ODR�DSP�S7cOF�FSET_CAR8t@�_�DIS���PEN_FILE�:�7�AF�PTION_IO��q��M_PRG %���%$*����M�W�ORK �yf ��춍��:�� � ����9���	 ����ڍ�It��RG�_DSBL  Ľ�C�{u��RI_ENTTO7 ��C� A �UT_SIM_Dy����V�LCT ��}{B �٭��_PEX�P=�ԷRAT�W dc|��UP ���
`���e�w�]ߛ�֩��$�2r�L6(L?���	l d����� �&�8�J�\�n��� ������������"�4�F�X���2�߈��� ����������*�<w�Tfx�� �����J`�ˣG���Tz�Pg��� ���/"/4/F/X/ j/|/�/�/�/���/ �/??0?B?T?f?x? �?�?�?�?�?�?�?�/ �/,O>OPObOtO�O�O �O�O�O�O�O__(_0:_��O��y_�]2ӆ��_�^�_�_�W�^]^]��/ooSog ��Hgrohozo�o�o�o��o�oF`�#|`��A�  9y����O�K�1�k������<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	O |�Q�s�r�q>��u
��q�F`H<zH~��H3k7GL��zHpG㎁99l7�k_B�T�F`C�4��k�H���t���-�Ae���k������s���  ��ሏ����EeBV�T���dZ���π���ڏ  ���q-�Fk�y�{Fb�U���n@6��  ����z�Fo��Be	'� �� ��I� ?�  �:p܋�=���ڟ웆�@���B�,���"B���g�AgN�����  '|���g��BU��p�BӀC׏�����@  #�yBu�&�ee�/^^މB:p2����>�m�6p�Z���Dz?o}�܏������׿@������Ǒ��� f�?  � �M���=*�?�ff�_8�J�ܿ 3pϑ�ñ�8�Чϵʖq.·�(����P���'��s�t�L�>��/�;�Cd�;��.<߈�<�g�<F+�<L ��^oiΚrd�@��r6p?fff?��?&�п�@���@x��@�N��@���@T����Z���ћtމ�u �߈w	�x��ti�>�)� b�M��q������� ������:�%�^��������W���S�E� � G�aF�� Fk���������1 U@yd��� ���q��	��{� A��h�����"a��ird��A{/@w/J/5/n/vA��aA���":t�/ C^/��/Z/ ލ?��`�/�/1??���W�����g��pE� ~1�?04�0
1�1�@IӀ��Bµ�WB]�NB2��(A��@�u�\?����������b�0�|�u�R����
�>��ؽ��B�u*C��$�)�`�? ����GC#����rAU�����1�eG���I��mH�� I:��I�6[F�﫹C4OI���J�:\IT��H
~QF�y��Ol@�*J��/ I8Y�I��KFjʻC�� -?�O�O__>_)_b_ M_�_�_�_�_�_�_�_ o�_(oo%o^oIo�o mo�o�o�o�o�o �o $H3lW�{ �������2� �V�h�S���w����� ԏ�������.��R� =�v�a�������П�� ��ߟ��<�'�`�K� ]���������ޯɯ�@�&�8�#�\��3(J�ϳ�3:a������J�3��c4�������������1�ǲ��ڿ��1����e���14 �{2�2�r�`ϖτϺϔ���%PR�P���! �h�!�K�6�o�Z�����u�|ߵߠ� ���������3��W� B�{�f�4���������d�A����!��1� 3�E�{�i��������������  2 E�f�7Fb�7�b�6B�!�!� C9� 	�� �0@�/`r� �����#x�� +=�3?, V*�8v��0�0�u�0�.
 D �����//%/ 7/I/[/m//�/�:�� ��ֻ�G����$PARAM_MENU ?2���  �DEFPU�LSE�+	WAITTMOUT�+�RCV? �SHELL_WR�K.$CUR_S�TYL� 4<OsPTJJ?PTB_?�Y2C/?R_DECSN 0�Ű<�?�?�? �?�?OO?O:OLO^O��O�O�O�O�O�!SS�REL_ID  �.�����EUSE�_PROG %��*%�O0_�CCCR�0�B���#CW_HO�ST !�*!HT�_=ZT��O_�Sh_�zQ�S�_<[_TI�ME
2�FXU� GDEBUG�@�+�C�GINP_FLM3SKo5iTRDo5gWPGAb` %l��tkCHCo4hTYPE�,� �O�O�o #0Bkfx� �������� C�>�P�b��������� ӏΏ�����(�:��c�^�p�����7eWO�RD ?	�+
 �	RSc`���PNS��C4�J9Ov1��TE�P�COL�է�2��g�LP 3������OjTRACECToL 1�2��! ��Ғ����q�DT Q�2��Ǡ��D � ��ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ����Я0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~�T�� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�3��$PGTRACELEN  �1�  ����0��6_UP �����A�@�1@�1_C�FG �ET�3�1
@�<D�0�<DZO<C�0uO$BD�EFSPD ��/L�1�0��0H�_CONFIG s�E�3 �0��0d�D��2 ��1�APpDsA�A�0���0IN'@TRL' �/MOA8pEQ�PE�E��G��A<D�AILID�(C�/M	bTGRP� 1ýI �l�1B  ������1A�33F�C� F8� E/�� @eN	�A�A�sA�Y�Y�A�@� �	 vO�Fg�_ #´8cokB;`ba�Bo,o>oxobo�o�1>о�?B/�o��o~�o =%<��
C@ yd��"���x���  Dz@� I�@A0�q� ������� ˏ���ڏ���7�"��4�m�X���|���Ú)�ґ
V7.10�beta1HF �@����Asq��Q  ��?� �BܠP�p� �C��&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@���f��N����ҡ�R�ܣΪRљ���1�i{������t<B�!CeQKNOW_M�  lE7FbTSV7 ĽJ�BoC _�b�t�����������P��1�]aSM�SŽK� ���	NB�0���ĿK���>-�bb��A �RP����0�Ŗά�bQMR�S��T��iN���d���V]S�T�Q1 1�K
� 4MU�iǨj� K�]�oߠߓߥ߷� ������2��#�h�G� Y��}�������
�P�����,�27�Iߎ�1�<t�H��P3 ^�p�����,�4��������,�5(:�,�6Wi{�,�7 ����,�8��!3,�MAD�6 �F,�OVLD � KD�xO.�P�ARNUM  p�MC/%�SCH� E
9'!G)�3Y%UPD/��E�/P�_CMP_��0@��0'7E�$ER_CHK�%5H�&�/��+RS���bQ_M�O�+?=5_'?O�__RES_G6��:� I�o�?�?�?�?O�? O7O*O[ONOOrO�O �O�{4]��<�?�O z5���O__|3 #_ B_G_|3V b_�_�_|3 � �_�_�_|3� �_�_�o|3Oo>oCo|2V� 1�:�k1!�@�c?�=2THR_�INRc0i!}�o5d޲fMASS�o Z��gMN�o�cMON�_QUEUE ��:�"�j0��O�N�� U1Nv�+DpE�NDFqd?`yEXEo`u� BEnpPAsOPTIOMwm;Dp�PROGRAM %$z%Cp}o(/~BrTASK_I���~OCFG ��$��K�DATA���T���j12 /ď֏������+� =�O�a�����������͟��INFO�����3t��!�3�E�W� i�{�������ïկ� ����/�A�S�e�w�(����Θ� '��FlJ�a K_N��T��˶ENBg ڽw1���2��GN�2��ڻ P(O��=���]ϸ�@y���v� �u��uɡdƷ_EDIT� �T�����G�W�ERFL�x�c)�RGADJ Ҷ�/A�  $�?j00���a�Dqձӆ5��?��ʨ�<u�)%e������F�f��2�R��	H;p�l�G�b_�>�pA�od�t$�*z�/� **:� j0�$�@�5Y�T���^��q�߈b~�L� ��\�n������� ��������4�F�t� j�|������������� bLBT�x ����:��$ ,�Pb��� /����/~/(/ :/h/^/p/�/�/�/�/ �/�/V? ??@?6?H? �?l?~?�?�?�?.O�? �?OO O�ODOVO�O zO�O_�O�O�O�O�O r__._\_R_d_�_�_ �_�_�_�_�f	g�io �pWo�o{d�o�~o��ozoB�PREOF �Rږp�p�
�IORITY��w[���MPDS1P�q��pwUT6��Ӿ�ODUCT3�e����OG���_TG��8��ʯrTOENT 1׶�� (!AF_�INE�p,�7�!�tcp7�_�!�udN���!�icmv��ޯrXY�K�ض���q)�a ,�����p�� &�	��R�9�v�]�o� ����П������*�H�N�`�*�sK��9}p�ߢ���Ư ,�!/6쒯�����خ��At�,  � Hp��P�b�t����u�w��HANCE !�R��:�wd��迄��2s�9Ks��PORT_NUM�s��p���_C?ARTREP{p�ξ��SKSTA�w �d�LGS)�����tӁpUn?othing��������{��TEMPG ޾y��'e���_a_seiban�o\��olߒ�}߶� ����������"��� X�C�|�g������ �������	�B�-�f� Q���u����������� ��,<bM� q��������(L�VERS�Iyp�w} �disabled�WSAVE ���z	2600H�768S?�!`ؿ����/ 	5(H�r)og+^/y�e{/ �/�/�/�/�*�,/�? �p���_�p �1�Ћ� �����Wh?z?�W^*pURGE��B�p�}vgu,�WF�0DO�vƲ�vW%��4(�C��WRUP_DEL�AY �\κ5R_HOT %Nf�q׿GO�5R_NORMAL&H�r6O�OZGSEMIjO�O�O�(qQSKIPF3��W3x=_98_J_ \_]�_�_{_�_�_�_ �_�_�_	o/oAoSoo woeo�o�o�o�o�o�o �o+=aOq �������� '��7�]�K��������)E�$RA{����K/�zĀÁ_PA�RAM�A3��K; @.�@`�61�W2C<��y���C�6$�BÀBT�IF�4`�RCVT�MOUu�c���ÀDCRF3��I� �+UC�A�qD��2=\��(?��]�;
�ޅ���4���+_���;�Cd;���.<߈<��g�<F+<L���Ѱ��d�u�L�������ϯ����)�;�M�_���R�DIO_TYPE�  M=U�k�EFPOS1 1�\�'
 x4/���� �+�$/<��$υ�p� ��D���h��ό��'� �����o�
ߓ�.ߤ� Rߌ�������5��� Y���i��*�<�v��� r���������U�@� y����8���\����� ������?��c����/2 1�KԿ�X�T�x��3 1����nY|�S4 1�'�9K�/�'/�S5 1���/�/�/�/:/S6 1�Q/c/u/�/-??Q?>�/S7 1��/�/�
?D?�?�?�?d?S8 1�{?�?�?�?WO�BO{O�?SMASK 1L��O�D�GXNO���F&�^��MOTEZ�Ż��Q_ǁ�%]pA݂��PL_RANG!Q�]�_QOWER ��ŵ�P1VSM_�DRYPRG �%ź%"O�_�UTA�RT �^�ZU?ME_PRO�_�_�4o��_EXEC_ENB  ��#�e�GSPD`O`WhՅ�jbTDBro�jRM��o�hINGVERSION Ź�#o�)I_AIoRPURhP �O\(�MMT_�@T�P�#_ÀOBOT__ISOLC�NTV�@A'qhuNAME��l��o�JOB_O�RD_NUM ?��X#qH�768  j1Z�c@�r�rV��s��r�?�r?�r�pÀPC_TIMEu�za�xÀS232>R�1�� L�TEACH PE�NDANw�:GX��!O Mai�ntenance_ Consj2���"��No UseB�׏�������1�C�y�V�NPO��P@�YQ�c�S�CH_L`��%^ �	ő��!OUD1:럒�R�@�VAIL�q@�Ӏ��J�QSPACE1w 2�ż ��@YRs�i�@Ct�YRԀ�'{��8�?� �˯����"���7� 2�c�u�����G���߯ ѿ򿵿�(��u�A C�c�u�����Ͻ�߿ ���ϵ��(��=�_� qσϕ�C߹������� ���$��9�[�m�� �ߣ�Q������߭���  ���	�W�i�{��� M�������5���. S�e�w�����I�� �����*? as��E��� ��/&//;/]o ������/2/�/ ?"?�/7?Y/k/}/�/ �/O?�/�/�?�?�?O�0OOKA��*S�YPpM*�8.3�0261 yB5/�21/2018 �A �WPfG|��H�_TX`� !�$COMME��$USAp� $ENABL{EDԀ$INN`�QpIOR�B�@RY~�E_SIGN_�`��AP�AIT�C�BW�RK�BD<�_TYyP�CRINDXSp�@W�@%VFRI{��_GRPԀ$U�FRAM�rSRTO�OL\VMYHOL��A$LENGT�H_VTEBTIR�ST�T  $�SECLP�XUFI�NV_POS�@$MARGI�A?$WAIT�`�Z�X2�\�VG2�GG1�AI�@�S�Q	g�`�_WR�BNO_US�E_DI�BuQ_R�EQ�BC�C]S$?CUR_TCQP�R�"a^f �GP_S�TATUS�A @ �A3`�BLk�H�$zc1�h�P@����@_�FX ��@E_MLT_C�T�CH_�J�`CO��@OL�E�CGQQ�$W�@w�b#tDEADLOCKu�DELAY_CNaT�a3qGt�a$wf� 2 R1R[1$X<�2[2�{3[3$Zwy�q%Y�y��q%V�@�c�@�b$V4�`�RV�UV3oh>b>�@ � �d�0NarMSKJ�LgWa�Z�C`NRK�PS_R7ATE�0$���S�
`�Q�TAC��PR�D���e�S*��a4�A�0�DG�A 08�P�flp bquS�2ppI�#`
`�P� 
�S\` � �A�R_ENB�Q �$RUNNER_AXI��<`ALPL�Q�RU�T�HICQ$FL�IP7��DTFER�EN��R�IF_C	HSU�IW��%V)�CG1����$PřA�Q��Pݖ_JF�P�R_P�	�RV_�DATA�A � $�ETIM|���$VALU$��	�OP_  � �A  2� �SC*��	� �$IT�P_!�SQ]PNPOU�}�o�TOTL�o�D�SP��JOGLI�b��PE_PKpc�O�f�i��PX]PTA�S�$KEPT_GMIR��¤"`M�b&�APq�aE�@��y�q�g@١c�q�PG�BRK6�x���L�I��  ?�SJ��q�P�ADEz�ܠB�SOCz�MOTN�v�DUMMY16�Ӂ$SV�`DE�_OP��SFSP�D_OVR
��f�@LD����OR��[TP8�LE��F��l����OV��SF��F����bF�d�ƣ&c�)�fQc�LCHDL}Y��RECOV���`��W�PM��gŢ�#RO������_F�?�� @v�S �NVsER�@�`OFS�PC,�CSWDٱc�ձ����B����TRG�|š�`E_FDO���MB_CM}���B��BLQ�¢	�Q�̄Vza�BUP�g��G
��AM���@`�KՊ�e�_M!�d�A�Mf�Q��T$CAԕ���DF���HB�Kd�v���IOU2��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�y3A��ATIO�0��͠��US����WaAB��R+c�`t��`DؾA��_AUX~w�SUBCPUP���S�`����3Եжc8���3�FLA�B�HW_Cwp"�Ns&��]sAa��$UN�ITS�M�F�AT�TRIz�Z�CY{CL�CNECA����FLTR_2_�FI��TARTU�PJp����A��LPx������_SCT*cF_F�F_P���b��FS��+�K�CHA�/Q��*�d�RS�D��Q����Q���_TH�PROr���հGEMPJ���G�T�� �Q�D�I�@y�RAILAiC/�bMX�LOf�xS��ځ���拁��V��PR#�S`appz�C� 	���FUNC���RI�N`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ngDAQ�B�rkLD�र&q�M�K���TI���j���$�@RIA_[SW��AF��Pñ#��%%�p9r1���MOIQ���DF_l~P(�PD"LM-�{FA�PHRDY�DORG�H; _QP|�s%MULSE~P�z���*�� J��J�ײ��FAN_A�LMLVG��!WR=N�%HARDP���UcO�� K2$SHADOW]�kp�a802��� STOf�+�Y_^�w�AU{`R<��eP_SBR�z5����:F�� �3MPINF?�\�4�λ3REGV/1DG��+cVm �C�CFL4(��?�DAiP���Z`�� �����Z�g	 �P(Q$�A$Z�Q V�@�[��
� ��EG0��o���kAAR�����2�axG��AX�E��ROB��RE%D��W�QD�_�Mh�CSYA��AF��FS�G�WRI�P~F&�ST�R����E�˰EH�H)��D�a\2kPB6P��=V��Dv�OTOr�1)���ARYL�`tR�v�3���FI&�~ͣ$LINKb!�\��Q�_3S��8�E��QXYZ2�Z�5�VOFF���R��R�XxPB��`ds�G�cFI�0�3g�������_J��'�ɲ�S&qR0LT2V[6���aTBja�"2�bC���DU�F]7�TUR� X���e�Q�2XP�ЊgFL�E���x@�`�U9Zy8���� 1	)�%K��Mw��F9���8������ORQj��G;W3���#�Ґd ����uz����1�tOV	E�q_�M��ё?C�u EC�uKB�v'0�x-�w H��t���& `��q ڠ�B�ё�u�q�wh�0ECh����ER��K�	�EP����AT�K�6e9e�W���AXs�'��v� /�R ����!��  ��P��`��`�3p�Yp�1�p�� � � �� (�� 8�� H� � X�� h�� x�� �������DEBU��$%3�I��·RA!B���ٱ�sV��� 
d�J、��@� ����������Q���a ���a��3q��Yq+$�`�%"<�cLAB0b8�u�'�GRO���b<��B_s��"T ҳ*`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Q`θuݸ��PNT0~���SERVE �NZ@ $`EAV�!�PO�����nP!�P@�$!Y@�  $>�TREQ�b
=��BG�K��%"2\��� _ � l��5�D6ESRRVb(�I��V0`�;���TOQ:�7�L��@
�R��e G�%ĩQ�� <�50F� �,�`�z�>�RA~� 2 d!�2����S�  M�`�pxU ����OCu�G�  ��C�OUNT6Q ]�P@FZN_CFG�F� 4#��6��T G4�_�=�����Î�^VC ���M ��"��$6��q ��F!A E� &��X�@� ������A����A9P��P@HEL�0�ҿ 5b`B�_BAS��RSR�6�CSH����1�Ǌ�2��3��4���5��6��7��8��}�ROO����Pf�PNLEA�cAB)�ܫ ��ACKu�IN2O�T��(B$UR0� =�_PU��!0��OU+�Pd�8j���� V��TPFWD�_KAR��� ��R�E(ĉ P�P�>QUE�:RO�p�`r0P1I� x�j�P�8f��6�QSEM��0t��� A��STYL�3SO j�DIX�&p�����S!_TMC�MANRQ��PE�NDIt$KEY?SWITCH����kHE�`BEA�TM83PE{@LEP��>]��U��F���SpDO_HOeM# O�@�EF�p�PRaB�A#PY�C�� O�!���OV_�M|b<0 IOCM��dFQ��h�HKYA D�Q�7��	UF2��M���p�c�FORC�3WAR�"�OM|@ � @S�#o0U)SP��@1�2&3&4RE���T�O��L�y��8UNLOv��D4K$EDU1  ��SY�HDDN�F� M�BLO�B  p�SN�PX_AS�� �0@�0��81$S{IZ�1$VA{�~��MULTIP-���# A� � $��� /4`��BS��0�C���&F'RIFBO�S����3� NF�ODBUP߰�%@3;9(���܋�Z@ x��SI���TEs�r�cSG%L�1T�Rp&�Н3xB��@�0STMTq2�3Pg@VBW�p�4�SHOW�5@�SmV��_G�� 3p�$PCJ�PИ���F�B�PHSP A�W�EP@VD�0WC�� ���A00 ��PB XG XG XGT$ XG5VI6VI7VIU8VI9VIAVIBVI@�XG�YF�0XGFVH���XbI1oI1|I1��I1�I1�I1�I1��I1�I1�I1�I1��I1�I1Y1Y2�UI2bI2oI2|I2�I2�I�`�X�I2p�X��I2�I2�I2�I2
�I2Y2Y�p�hbIU3oI3|I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3�IU3Y3Y4�i4bIU4oI4|I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4�IU4Y4Y5�i5bIU5oI5|I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5�IU5Y5Y6�i6bIU6oI6|I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6�IU6Y6Y7�i7bIU7oI7|I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7�I�7Y7T��VP� UD�y"ՠ��Q
<A62��t��R��CMD� ��Mb5�Rv�]��Q_hЁR���e����<�Y�SL���  � �%\2��+4�'��xW�BVALU���b��'���FH�ID�_L���HI��I���LE_��㴦��$0C�SAC��! h �VE_BLCK��1>%�D_CPU5ɧ  5ɛ �����C�� ���R " � �PWj��#0��LA��1SBћì���R?UN_FLG�Ś� ���ĳ ���������šH���Х��T�BC2��# � @ B��e �S�88=�FTDC�����V���3d�Q�TH�F�����R�L�ESERVE9��F���3�2�E��Н��X -$��LEN`9��F��f�RA��LW"G�W_5�b�1�њд2�MO-�T%S60U�Ik�0�ܱF�����[�DEk�21LA3CEi0�CCS#0�� _MA� j��z玤�TCV����z�T �������.Bi�'A�$z�'AJh�#EM5���J��@@i�V�z���2Q �0&@o�h��JK��VK9��{����щ�J0����J�J��JJ��AAL����������4��5�ӕ N1������J.�LD�_�1* v�CF�"% `�GROU���1�A�N4�C�#m REQ�UIR��EBU��#��6�$Tk�2�$���zя #�&{ \�APPR� �C� 0�
$OPE=N�CLOS��St��	i�
��&' �MfЩ���W"N-_MG�7CB@��A���BBRK�@NOLD@�0RTMO_5ӆp1	J��P�����@���������6��1�@ )!�#�(� ������'��+#PATH ''@!6#@!�<#� � 9'��1SCA��l�6IN��UCJ�[1� C0@UM�(Y  ��#�"�����*���*���� PAYLOA�~J2LؠR_A	N^�3L��91�)�1AR_F2LSHg2B4LO4�!F7��#T7�#ACRL_@�%�0�'�$��H���.�$HA�2FL�EX��J!�) P�2�D߽߫��|�0��* :�� ��z�FG]D����z���%�F1]A�E�G4�@F�X�j�|���BE�� �����������(� �X�T*�A���@�XI��[�m�\At�T$g�QX <�=��2TX���emX �������������������+	�J>+ �-�K]o|�٠cAT�F�4�ELFP�Ѫs�J� *� J�EmCTR�!�AT�N�vzHAND_VB.��1��$7, $8`F2Avԍ��SW�
"-?� $$M*0. �]W�lg��PZ����A��� 1����:QAK��]AkAzP��LN�]DkDzePZ G��C�ST_hK�lK�N}DY�� � A����0��<7]A <7W1�'��d�@g`�P��������" 1B$. �M�2D%"��H����A'SYMj%0�� j&!-��-W1�/_�{8 � �$�����/�/�/�/ 3J<�:9�/�\89�D_VI�v�|���V_UNI�����cD1J����╴� W<��n5Ŵ�w=4��9 ��?�?<�uc�4�3���%�H���/0�j��0�DIzu�O����k�>0) �`��I��A��# ���@ģ���@��IP�l� 1 � /�ME.Qp��9�ơT}�PT�;pG �+ Gt� ���'���T�0 $�DUMMY1��o$PS_�@RF�@�;�$b�'FL�A@ YP(c|��?$GLB_TP�ŀ����9 P�q��2c X� z!ST9��� SBRM M2�1_V�T$SV_ER*0O�p����SCL����AGPO�¶f�GL~�EW>�3s 4H �$Yr�ZrW@�x�A1+�A����";�"�U&�4 �8`NZ�"�$G�I�p}$&� p-� �Y�>�5 LH \{��}$F�E��NEAR(PN�CF<��%PTANC�B;��JOG�@� 6�9�$JOINT�wa?pat �MSE]T>�7  x�E��HQtpS{r��up>�8�� �pU.Q?��� LOCK_F�OV06���BGLV��sGLt�TEST�_XM� 3�EMP������_�$1U&@%�w`24� Y�B��5��2�d��3���CE- ���� $K�AR�QM��TPD�RA)�����VECXn@��IU��6��{HEf�TOOL�C�2V�DRE IS�3ER6��@AC)H� 7?Ox ӦQ�29Z�H I� � @$RAIL__BOXEwa�oROBO��?��?HOWWAR�1�<_�zROLMj���:qw�jq� �@ O{_Fkp! d�l>�9��
 R OB8B:��@�c�KOU�;�Һ�3ơ��r�q_�$PIP��N&`H�l�@���#@CORDED�d�p >f�fpO�� �< D ��OB⁴sd���Kӕи��qSYS�A�DR�qf��TCH�t� = ,8`E�No��1Ak�_{��-$Cq=GSf�VW�VA��> � � &��PREV�_RT�$ED�ITr&VSHWRBkq�֑ &R:�v��D��JA�$�a$HEAD�6�� ��z#KE:�E�CPwSPD�&JMP��L~��0R*P��?���1%&I��S�rC��pNE; �q�wTICK�C��M�1��5{HN��@ @�8 1Gu�!_GPp6���0STY'"xLO��:�2l2?�A tk 
m G3%%$R!�{�=��S�`!$@��w`���ճ���Pˠp6SQU��E��u��TERC����T=SUtB ����@hw&`gw�Q)�pOЌ���@IZ��{��^�PR�kюB1XsPU���E_DO���, XS�K~�AXiI�@���UR�p�GS�r� ^0�&��p_,) �ET�BPm��Jo��0Fo��0A|����Rԍ��a�<�SR�Cl>@P��b_�yUr��Y ��yU��yS��yS���U Ї�U���U���U�]���Ul[��Y�bXk�]C�m�����YRSC��� D h�D1S~0��Q�SP���eATހ���A]0,2~N�ADDRES<=B} SHIF{s��_2CH�p�I\��=q�TVsrI��AE"���a�CT�
���
;�VW�A��F 	\��q��0l|\A@�rC�_B"R{zp����q�TXSCRE�E�Gv��1TICNA���t{�@ �3Q_�b?�H T 1�ЂB�����I��Ap��BE�y RRO������� B���1UE�4I �g�!p�S���RSM]0�GU�NEX(@~Ƴ�j�S_S�ӆ��Á։񇣣��ACY�0� 2-H�pUE;�J���\��@GMT��Lֱ��A��O*BBL�_| W8���K �Լ0s�OM��LE�/r��� TO!�s�RwIGH��BRD
�%qCKGR8л�T�EX�@����WIDTH�� �B�|�<���I_��Hi� OL 8K���_�!=r���R:�_��HYґ��O6q�Mg0I紐U��h�Rm��LUMh��FpE#RVw��P���`��N��&�GEU�R��FP)�)� LIP��(RE%@�a)ק@�a�!��f �5�6�7�8Ǣ#B�à�@���tP�fW�Sv@M�USR&�OO <����U�Qs�FOC)��P�RI;Qm� :���T�RIP�m�U)N����Pv��0���f%��'���@�0 qQ����AG �0aT� �a>q�OSт%�RPo���8�R�/�A�H�L4����U¡�SU�g��¢5N��OFF���T��}�O�� 1R������S�GUN��-6�B_SUqB?���,�SRTN��`TUg2��mCOR�| D�RAUrPE�T<Z�#'�VCC��	3�V AC36MgFB1�%d�PG ��W (#��AST�EM�����0P�E��T3G�X �<\ ��MOVEz�A��AN�� ���M�>��LIM_X��2� ��2��7�,�����ı�
�BVF�`E�XQ�~��04Y��IB(�7���5S��_Rp� x2��� WİGp+@��}СP��3�Zx ���3A���A�ݠCZ��DRID����V�y08�90� De�MY_UBYd���6�ш@��!��X��P�_S��3��L�KB�M,�$+0DEY�(#EX`�����UM_MU� X����ȀCUS�� ���G0`PACI���а@�Հ:��:,�:����RaE/�3qL�+C���:[��TARGB��P�r ����R<�\ d`��A��$�i	��AR��SW2 $��-��@Oz�%qQA7p�yREU�U�0�1�,�HK�2]g0�qP� N� �sEAM0GWOR����MRCV3�^� ���O�0M�C��s	���|�REF_���x(�+T�  ���������3_RCH4(a�P@�І�hrj�NA�2��0�_ ��2����L@4��n�@@OU~7w�6���Z��a2[ư�RE�p�@;0\��c�a'2K�@SUL���]��C��0�^��� NT��L�3��@(6I�(6q�(3� L��@Q5��Q5I�]7q�}�)Tg`4D`�0.`0ПAP_HUC�5S]A��CMPz�F�6(�5�5�0_�aR��a��1I\!X�9��VG�FS��ad †M��0p�UF_`x��B� �ʼ,RO���Q��'����UR�3GR�`.�3IDp���)�D�;��A��~�IN��H{D���V@@AJ���S͓UW�mi=�����TYL�O*�5����bot +�cPA�{ �cCACH� vR�UvQ��Y��p�#�CF�I0sFR�XT8���Vn+$HO����P!A3�XBf�(01 ���$�`VPy� �^b_SZ313he6K3he12J�eh chlG�chWA�UMP�j���IMG9uPAyD�iiIMRE�$^�b_SIZ�$P�����0 ��ASYNB{UF��VRTD)u�5tqΓOLE_2�DJ�Qu5R��C��U���vPQuECCUlVEMV �U�r��WVIRC�aIuVTPG���rv1s���5qMPLAqa��v�ԂV0�cm� CKLAS�	�Q�"���d  �ѧ%ӑӠ@�}¾�$�Q���Ue A|�0!�rSr�T�# 0! �r�iI��ml�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f �� >֦3�@Sp�SgLOW>�RO��ACCE���!� 9��VR�#���p:���A1D�����PAV�j��� D����M_B8"���^�JMPG ���g:�#E$SSC@��F�vPq��hݲ�vQS�`qVN��L;EXc�i T`�s�r���Q�FLD �DEsFI�3�0�2���:���VP}2�Vj� �A���V�4[`MV_PIs��t���A�@&��FI��|�Z��Ȥ������A���A��~�G9Aߥ1 LOO��1 JCB���Xc��^`�#PLANE��R��1F�c�����pr�AM� [`�噴��S�� ��f����Af��R�Aw��״tU��pRKE<��d�VANC�A\���� k����ܲϡ�R_AA� l��2� ��p�#B�Gm h�@��O K�$�������kЍ0OU�&A�"A�
p�pSuK�TM@FVIEM 2l ��P=��҇n <<��dK�U�MMYK1P���`D��ACU���#AU��o $��TIT�$�PR����OP��?�VSHIF�r�p`J�Qsԙ�lfOxE$� _R�`U�#����s��q�������G�"G�޵'�T��$�SCO{D7�CNTQ i�l�>a�-� a�;�a�H�a�V���T1�+�2u1��D��ܲ��  � SMEO�Uq��a�JQЖ����a_�R[�r4�n�*@LIQ�AA^/`�XVR��s��n�TL�t�ZABC�t�t�c��
AZIP��u,���LVbcLn"��TED�ZMPkCFx�v:�$��� ���DMY_L�N������M�Ay�w� Ђ(a�u� MC�M�@CbcCART�_�DPN� '$J71D��=�NGg0Sg0�BUX�W� ��UXEUL|ByX��М	��H�Z��xC 	���m�YH�}Db  y 80<���0EIGH�3n�#?(� H����$�z ���|�����$%B� Kd'��_��L3�RVS�F`���OVC�2'�$|Ј>P&��
q���5D&�TR�@ �V�1��SPHX��!{ ,p� *<�$R�B�2 2 ����C!�  �@V+H�b*�c%g!`+g"�`�V*�,8�?� V+�/V.�/�/?�/�/V(7%3@/R/d/v/�/ 6?�/�/�?�?�?O4OOION;4]?o?�?�? �?SO�?�?�O_�O0_Q_8_f_N;5zO�O�O �O�Op_�O_o8o�_ MonoUo�oN;6�_�_ �_�_�_�oo%o4U@j�r�N;7�o �o�o�o�o� BQ��r�5���������N;8 �����Ǐ=�_� n���R���ş��ڟN;�G � џ�
����?��� W�i�{�������ï� .�������A��dW�<�N�|������� Ŀֿ�ޯ���0� B�_�R�d�꿤϶��� ����������*�L� ^��rτ�
������� �����&�8�J�l��~� `ҟ @ �з����ߩ��-����&�,���9� {�����a��������� ������A'Y �������@��a#1�
����N;_MODE � ��S "��[�Y�B���
/\/*	|/�/R4CWORK_AD��	�T1R  ����� �/� _?INTVAL�+$���R_OPTI[ON6 �q@�V_DATA_G�RP 27���D��P�/~?�/�?�9 ��?�?�?�?OO;O )OKOMO_O�O�O�O�O �O�O_�O_7_%_[_ I__m_�_�_�_�_�_ �_�_!ooEo3oioWo yo�o�o�o�o�o�o �o/eS�w �������+� �O�=�s�a������� ͏���ߏ��9�'��I�o�]�����$S�AF_DO_PULS� �~������CAN_TIM������ SCR ��������5�;#U! P"�1!��� �?E� W�i�{�����.�ïկ`�����'(~�ET"2F���dR�DI�Y��2�o+@a�@������)�u��� k0~ϴ��_ ��  T� � �2�D�~)�T D��Q� zόϞϰ��������� 
��.�@�R�d�v߈���/V凷������߽��R�;W�o �W�p���
�t��Di�z$� �0 � �T"1!������ ������������ *�<�N�`�r������� ��������&8 J\n����� ���"4FX ��࿁���� ���/`4�=/O/ a/s/�/�/�/�/�/�/�!!/ �0޲k�ݵu� 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  ok$o6oHoZolo~o �o�o�o�o1/�o�o  2DVhz�/5 ?�������� &�8�J�\�n������� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q�0c�u��� ���`� ��ϯ����)�;� M�_�q���������˿ݿ� ����3� ���&2,��	�1234567�8v�h!BW!��2�Ch���0�ϵ��������� �!�3�9ѻ�\�n߀� �ߤ߶���������� "�4�F�X�j�|�h�K� ����������
��.� @�R�d�v��������� �����*<N `r������ �&��J\n �������� /"/4/F/X/j/|/; �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�/�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_�?L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o =_�o�o�o�o�o�o  2DVhz�����h�������u�o.�@�R���C�z  B��  � ���2&� �� _�
���/  	�_�2�Տ�����_�p������ďi�{����� ��ß՟�����/� A�S�e�w��������� N������+�=�O� a�s���������Ϳ߿����'�9�K�_�������<v�_��$�SCR_GRP �1
� �� t ���� ��	 _����� �����������_���p���)�a����~&�DE� DW8����l�&�G�CR�-35iA 90�12345678�90��M-20���8��CR35 ��:�
��������������:֦� Ӧ�G���&������	��]�o����~:���H���>�����������&���ݯ:��j���`��g������B�t�!���������A�����  @�`��@�� ( ?�=��H�t�P
��F@ F�`z�y��� ��� �$H ��Gs^p��B��7��/� 0//-/f/Q/�/u/�/ �/�/8���P�� 7%?����"?W?-2?<���]? H�14�?t�ȭ7�������?-4A, �&E$@�<�@G�B-1A 3OZOlO-:HA�H��O�O|O P�B(��B�O�O_��EL_�DEFAULT � �����`SHOTS�TR#]JA7RMIP�OWERFL  �i�/UYTWFD�O$V /URRV�ENT 1�����NU L!DUM_EIP_�-8�j!AF_�INE#P�_-4!�FT�_->�_;o!���`o �*o�o!�RPC_MAI�N�ojh�vo�o�cV�IS�oii��o!7TPpPU�Y�dk!
PMON_PROXYl��VeZ�2r��]f���!RDM_'SRV��Yg�O�G!R��k��Xh>����!
�`M��\i����!RLSY3NC�-98֏3��!ROS�_-<�y4"��!
CE4p�MTCOM���Vk�n�˟!	��CON�S̟�Wl���!>��WASRC��V�m�c�!��US	Bd��XnR���Noӯ �������!��E���i�0���WRVICE_KL ?%�[� (%SVC�PRG1��-:Ƶ2�ܿ�˰3�	�˰4�,�1�˰5T�Y�˰6|ρ�˰7�ϩ�˰��$���9����ȴf� !�˱οI�˱��q�˱ ϙ�˱F���˱n��� ˱���˱��9�˱�� a�˱߉��7߱�� _��������)� ���Q����y��'� ���O����w���� ������˰�� İd�c����� �=(as^ ������/� /9/$/]/H/�/l/�/ �/�/�/�/�/�/#?? G?2?k?V?}?�?�?�? �?�?�?O�?1OCO.O gORO�OvO�O�O�O�O��O	_�O-_��_DE�V �Y��MC:5X�`>GTGRP 2SVK ���bx 	�� 
 ,�PK  5_�_�T�_�_�_o�_ 'o9o o]oDo�ohozo �o�o�o�o�o�o5 {�_g���� ������?�&� c�u�\�������Ϗ�� �J\)���M�4�q� ��j�����˟ݟğ� �%���[�B��f� �����ٯ������� 3��W�i�P���t��� ÿ���ο���A� (�e�L�ί��RϿ��� ������� ��O�6� s�Zߗߩߐ��ߴ��� ���'�~ϐ�]��� h����������� ��5��Y�@�R���v� ��������@�	�� ?&cu\��� �����;M 4qX������ �/�%//I/[/B/ /f/�/�/�/�/�/�/ �/�/3??W?�L?�? D?�?�?�?�?�?O�? /OAO(OeOLO�O�O�O��O�O�O�O�O_"Ud� �NLy�6� * 		S=>��+c"_VU@Tn_�Y_B���B�2��J�j~Q´�~_g_�_�Q%JOGGING�_�^7T�(?VjZ�Rf=��Y���/e�_%o7e�Tt�]/o�o{m �_�o�m?Qi�o�o`;)Kq%��o �}os����� �9�{`��)���%� ��ɏ���ۏ�S�8� w��k�Y���}���ş ���+��O�ٟC�1� g�U���y������� '����	�?�-�c�Q� ��ɯ����w���s�� ��;�)�_ϡ���ſ OϹϧ��������� 7�y�^ߝ�'ߑ�ߵ� ���������Q�6�u� ��i�W��{����� �=��M���A�/�e� S���w���������� ��=+aO� �����u��� 9']���M ������/5/ w\/�%/�/}/�/�/ �/�/�/=/"?4?�/? �/U?�?y?�?�?�?? �?9?�?-OO=O?OQO �OuO�O�?�OO�O_ �O)__9_;_M_�_�O �_�Os_�_�_o�_%o o5o�_�_�o�_[o�o �o�o�o�o�o!coH �o{���� ��; �_�S�A� w�e�������я��� 7���+��O�=�s�a� �����П����� '��K�9�o������� _���[�ɯ���#�� G���n���7������� ��ſ����a�Fυ� �y�gϝϋϭϯ��� ��9��]���Q�?�u� cߙ߇ߩ���%���5� ��)��M�;�q�_�� �߼��߅������%� �I�7�m������]� ����������!E ��l��5���� ���_D� we�����% 
//���=/s/a/ �/�/�/��/!/�/? ?%?'?9?o?]?�?�/ �?�/�?�?�?O�?!O #O5OkO�?�O�?[O�O �O�O�O_�O_sO�O j_�OC_�_�_�_�_�_ �_	oK_0oo_�_co�_ so�o�o�o�o�o#o Go�o;)_Mo� ���o���� 7�%�[�I�k������ ����ُ���3�!� W���~���G�i�C��� �՟���/�q�V��� ���w��������ѯ �I�.�m���a�O��� s�������߿!��E� Ͽ9�'�]�Kρ�oϑ� ����Ϸ����5� #�Y�G�}߿Ϥ���m� ��i������1��U� ��|��E������� ��	���-�o�T���� ��u����������� G�,k���_M�q ������ �%[Im�� �	���//!/ W/E/{/��/�k/�/ �/�/�/	???S?�/ z?�/C?�?�?�?�?�? �?O[?�?RO�?+O�O sO�O�O�O�O�O3O_ WO�OK_�O[_�_o_�_ �_�__�_/_�_#oo Go5oWo}oko�o�_�o o�o�o�oC1 Sy�o��oi�� ���	�?��f�x� /�Q�+���Ϗ���� �Y�>�}��q�_��� ����˟���1��U� ߟI�7�m�[�}���� ǯ	��-���!��E� 3�i�W�y�ϯ��ƿ� �������A�/�e� ����˿UϿ�Q����� ����=��dߣ�-� �߅߻ߩ�������� W�<�{��o�]��� �������/��S��� G�5�k�Y���}����� ����������C1 gU������{� ���	?-c� ��S����� �/;/}b/�+/�/ �/�/�/�/�/�/C/i/ :?y/?m?[?�??�? �?�?? O??�?3O�? COiOWO�O{O�O�?�O O�O_�O/__?_e_ S_�_�O�_�Oy_�_�_ o�_+oo;oao�_�o �_Qo�o�o�o�o�o 'ioN`9� �����A&�e �Y�G�i�k�}����� ׏���=�Ǐ1��U� C�e�g�y����֟� ��	���-��Q�?�a� ��ݟ��퟇��ϯ� �)��M���t���=� ��9���ݿ˿��%� g�Lϋ���mϣϑ� ��������?�$�c��� W�E�{�iߟߍ߯��� ���;���/��S�A� w�e���������� ����+��O�=�s��� ����c����������� 'K��r��;� ������#e J�}k��� ��+Q"/a�U/ C/y/g/�/�/�//�/ '/�/?�/+?Q???u? c?�?�/�?�/�?�?�? OO'OMO;OqO�?�O �?aO�O�O�O�O__ #_I_�Op_�O9_�_�_ �_�_�_�_oQ_6oHo �_!o�_io�o�o�o�o �o)oMo�oA/Q Se����%{�,p�$SERV�_MAIL  �+u!��+q�OU�TPUT��$�@�RV 2v�v  $� (�qx�}��SAVE7��(�TOP10 2�W� d 6' *_�π(_�� ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u�������0��Ͽݷ��YP��'��FZN_CFG ;�u$�~�����GRP 2��D� ,B �  A[�+qD;�� B\��  B�4~�RB21ފ�HELL��u��j�k�2�����%RSR������ �
�C�.�g�Rߋ�v� ���߬�����	���-��?�Q��  �_�%Q���_����,p�������g�2,pd�����HK 1�� ��E�@�R�d����� �������������*<e`r���OMM ������FTOV_ENB��_���HOW_R�EG_UI�(�IMIOFWDL� ��^�)WAIT����$V1��^�NTIM����VA�_)_�UNIT����L]CTRYB��
�MB_HDDNw 2W� 2� �:%0 �pQ/�qL/^/ �/�/�/�/�/�/�/�"�!ON_ALIA�S ?e�	f�he�A?S?e?w?�:/? �?�?�?�?�?OO&O 8OJO�?nO�O�O�O�O aO�O�O�O_"_�OF_ X_j_|_'_�_�_�_�_ �_�_oo0oBoTo�_ xo�o�o�o�oko�o�o ,�oPbt� 1������� (�:�L�^�	������� ��ʏu�� ��$�Ϗ 5�Z�l�~���;���Ɵ ؟����� �2�D�V� h��������¯ԯ� ��
��.�ٯR�d�v� ����E���п���� ��*�<�N�`�r�ϖ� �Ϻ���w�����&� 8���\�n߀ߒߤ�O� ����������4�F� X�j�|�'������� ������0�B���f� x�������Y������� ��>Pbt ������ (:L�p��� �c�� //$/� H/Z/l/~/)/�/�/�/ �/�/�/? ?2?D?V?�]3�$SMON_�DEFPRO ����1� *SY_STEM*0m6�RECALL ?�}9 ( �}�4xcopy f�ra:\*.* �virt:\tm�pback�1=>�147.87.1�49.40:93�08 �1 �815�172]?O+M}8��4s:orderfil.dat�<`�?�?O�O�O}/�2mdb:�?cO�0oO�O_$_7D3�5�?�? �5�O_�_�_;@�?O_ a_t_�_o)o<ONO�O �Oo�o�o�OUo�Opo �o%8_�_�_n_  ���_GY�_~��!�4g
xyzra?te 61 �� � �����6e?�_�?17516 _�q�����&�9btpdisc 0ɏہݏ�������7dtpconn 0 H�@Z�l�~��!�4g9?o�QoG�ہ������/l0 �oZ�Ҋp����%��|��Z�ֆ������� }5�P�b�u�����*�}<��γout�put\test�_server.�pcà: oY� �ߐ6279142�4:263469 ���ϟ�2�D�̟ͯ z��߰�¯����� �ߛ�.�@�ӿd�v߈� �߾��������ߊ� �������a�w��� -�?���c�������� ��P�]��߅�(;� ����q���9�K�]o�$��ߝ27168ޞ�� �����R�Sy
// /�A��T�/�/�/r8c6��empY�7680 v/�/?:�/.�&*.d�/�.`�/ ?�?�?�1 J? \?n?�?O#O6ȏ�2 �?�?O�O�O��T/ �(zO__0/B/�O�' �O_�_�_����YD u_�_o*o=�_�_tA �_+o�o-�?��)]ooo �o$���o�o�o�o����u�$SNP�X_ASG 2�����q�� P 0 �'%R[1]�@1.1��y?��s%�!��E�(�:� {�^�������Տ��ʏ ���A�$�e�H�Z� ��~���џ����؟� +��5�a�D���h�z� ����ů�ԯ���
� K�.�U���d������� ۿ������5��*� k�N�uϡτ��ϨϺ� �����1��U�8�J� ��nߕ��ߤ������� ���%�Q�4�u�X�j� ������������� ;��E�q�T���x��� ��������% [>e�t��� ���!E(: {^������ /�/A/$/e/H/Z/ �/~/�/�/�/�/�/�/ +??5?a?D?�?h?z? �?�?�?�?�?O�?
O KO.OUO�OdO�O�O�O �O�O�O_�O5__*_ k_N_u_�_�_�_�_�_ �_�_o1ooUo8oJo��ono�o�o�d�tPA�RAM �u}�q �	��jUP�d9p�ht���pOFT_KB_CFG  �c��u�sOPIN_S_IM  �{v�n��p�pRVQSTP_DSBW~�r"t�HtSR �Zy � &�!pOB195_S�ERV M����vTOP_ON_?ERR  uCy~8�PTN Zu�k�A4�R?ING_PR�D���`VCNT_GOP 2Zuq�!px 	r��ɍ����׏��wVD��RP' 1�i p�y ��K�]�o��������� ɟ۟����#�5�G� Y���}�������ůׯ �����F�C�U�g� y���������ӿ�� 	��-�?�Q�c�uχ� �ϫ����������� )�;�M�_�qߘߕߧ� ����������%�7� ^�[�m������� ������$�!�3�E�W� i�{������������� ��/ASew ������� +=Ovs�� �����//</ 9/K/]/o/�/�/�/�/ �/�/?�/?#?5?G? Y?k?}?�?�?�?�?�?��?�?OO)�PRG�_COUNT8vq�k�GuKBENB���FEMpC:t}O_UP�D 1�{T  
4Or�O�O�O_ _!_3_\_W_i_{_�_ �_�_�_�_�_�_o4o /oAoSo|owo�o�o�o �o�o�o+T Oas����� ���,�'�9�K�t� o���������ɏۏ� ���#�L�G�Y�k��� ������ܟן���$� �1�C�l�g�y����� ����ӯ����	��D� ?�Q�c���������Կ Ͽ����)�;�d��_�q�=L_INFO� 1�E�@ �2@����������� �ٽ`y*��d�h'����¬��=`y�;MYSDEBUG�U@�@���d�If�S�P_PASSUE�B?x�LOG U ���C��*�Α�  ��A��UD1:\�ԘΥ�_MPC�ݵE&�8A��V� �A�SAV !�����l��X���SVZ��TEM_TIME� 1"���@ �0  iX���������$T1S�VGUNS�@VE'��E��ASK_?OPTIONU@�Et�A�A+�_DI���qOG�BC2_GRP 2#�I�����?@�  C���<K~o�CFG %z�Ɠ� �����`��	�.>dO �s������ �*N9r]� ������/� 8/#/\/n/v$Y,�/ Z/�/�/H/�/?�/'? ?K?]�k?=�@0s?�? �?�?�?�?�?O�?O O)O_OMO�OqO�O�O �O�O�O_�O%__I_ 7_m_[_}__�_�_�X � �_�_oo/o�_So Aoco�owo�o�o�o�o �o�o=+MO a������� ��9�'�]�K���o� ��������ɏ���#� �_;�M�k�}������ ��ß�ן��1��� U�C�y�g��������� ������	�?�-�c� Q�s����������Ͽ ����)�_�Mσ� 9��ϭ�������m�� �#�I�7�m�ߑ�_� �ߣ����������� !�W�E�{�i����� ����������A�/� e�S�u�w��������� ����+=O��s a������� 9']Kmo �������#/ /3/Y/G/}/k/�/�/ �/�/�/�/�/??C? ��[?m?�?�?�?-?�? �?�?	O�?-O?OQOO uOcO�O�O�O�O�O�O �O__;_)___M_�_ q_�_�_�_�_�_o�_ %oo5o7oIoomo�o Y?�o�o�o�o�o3 !CiW��� ������-�/� A�w�e���������� я���=�+�a�O� ��s�������ߟ͟� �o�-�K�]�o�ퟓ������ɯ���צ���$TBCSG_G�RP 2&ץ�  ��� 
 ?�   6�H�2�l�V���z���@ƿ�������(��d�E+�?~�	 HC����>���G����C�  A�.�e�q�wC��>ǳ33��"S�/]϶�Y��=Ȑ� C\  Bȹ���B���>���X�P���B�Y�z�"�L�H�0�$���� J�\�n�����@�Ҿ ���������=�Z�%�07����?3������	V3.0�0.�	cr35��	*����
���0������ 3���4�   {�CaT�v�}��J2��)������CFG� +ץ'� �*������I����.<
 �<bM�q�� �����(L 7p[���� ��/�6/!/Z/E/ W/�/{/�/�/�/�/.� H��/??�/L?7?\? �?m?�?�?�?�?�? O O$O�?HO3OlOWO|O �O����Oӯ�O�O�O !__E_3_i_W_�_{_ �_�_�_�_�_o�_/o o?oAoSo�owo�o�o �o�o�o�o+O =s�E���Y� ����9�'�]�K� m�������u�Ǐɏۏ ���5�G�Y�k�%��� }�����ßşן��� 1��U�C�y�g����� ��ӯ������	�+� -�?�u�c��������� �Ͽ���/�A�S� ����qϓϕϧ����� ���%�7�I�[��� mߣߑ߳������߷� �3�!�W�E�{�i�� ������������ A�/�e�S�u������� ��������+ aO�s��e�� ���'K9o ]������ �#//G/5/k/}/�/ �/[/�/�/�/�/�/? ?C?1?g?U?�?y?�? �?�?�?�?	O�?-OO QO?OaO�OuO�O�O�O �O�O�O___M_� e_w_�_3_�_�_�_�_ �_oo7o%o[omoo �oOo�o�o�o�o�o !3�o�oiW�{ �������/� �S�A�w�e������� я�������=�+� M�s�a���������ߟ �_	���_ן]�K� ��o�������ۯɯ�� �#���Y�G�}�k� ����ſ׿������ ��U�C�y�gϝϋ� �ϯ��������	�?� -�c�Q�s�u߇߽߫� �������)��9�_� M����/����i�� ����%��I�7�m�[� ���������������� ��EWi{5� ������� A/eS�w�� ���/�+//O/ =/_/a/s/�/�/�/�/ �/�/?'?��??Q?c? ?�?�?�?�?�?�?�? O�?5OGOYOkO)O�O�}O�O�O�O�N  �@S V_R��$TBJOP_�GRP 2,�E��  K?�V	-R4S.;\{��@|u0�{SPU >�<�UT @�@LR	 �C� �Vf  C���U<LQLQ>�33�U�R�����U�Y?�@=��ZC��P���ͥR��P  Bq��W$o/gC��@g�dDb�^Ǚ��eeao�P&f�f�e=�7LC/�kaB o�o�P���P�efb-C�p���^g`�d�o�PL��Pt<�eVC\[  �Q@�'p�`�  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�ana�a`C�;�`L �w�aQoxp�x�p?:��XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb��� �X�	��1��)�W� ��c����������� �󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSocr35QT*��QT�A�� E��'E�i�F�V#F"wqF�>��FZ� F�v�RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG�G#
��D��E'
�EMKE����E�ɑE�ۘ�E��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF�u��<#�
<t���ٵ=�_��V �R�p�V�9� ]ESTPARbtp�HFP*SHR\�ABLE 1/;[I%�SG�� �W�G�G�G� WQ*G�	G�
G�GȖ�*QG�G�G�ܱNv�RDI~�EQ��@�Ϲ�������W�O_߀q�{ߍߟ߱���w�S]�CS !ڄ���� ��������&�8�J� \�n�������������  ]\�`��	��(� :�����
��.�@�w�~NUM  �E�EQ�P	P �۰ܰw�_CFG �0��)r-PIM?EBF_TTb��8CSo�,VERڳ-zB,R 11;[O 8��R�@2� �@&  �� �����//)/ ;/M/_/q/�/�/�/�/ �/?�/?J?%?7?M? [?m?>�@�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_H�_�_l_�Y@c�Y�MI_CHA�N8 c cDB'GLV��:cX��	`ETHERADW ?f�\`���?�_uo�oQ�	`R�OUTV!	
!��d�o�lSNMA�SKQhcba255.uߣ'9ߣ�Y�OOLOFS_�DIb��U;iOR�QCTRL 2$		�Ϸ~T�� ���#�5�G�Y�k� }�������ŏ׏������.��R�V�PE?_DETAI/h|z�PGL_CONF�IG 8�	����/cell/�$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c�u��� ��(���ϯ���� ��;�M�_�q�����$� 6�˿ݿ���%ϴ� I�[�m�ϑϣ�2��� �������!߰���W�@i�{ߍߟ߱�%}F� ������/�A�C�i�H�Eߞ������ ����?��.�@�R�d� v�������������� ��*<N`r� ������ &8J\n��! �����/�4/ F/X/j/|/�//�/�/ �/�/�/??�/B?T? f?x?�?�?+?�?�?�? �?OO�?>OPObOtO��O�O�O���U�ser View� ��}}1234?567890�O�O �O_#_5_=T�P��]_���I2�I:O�_�_��_�_�_�_X_j_�B3 �_GoYoko}o�o�o o�op^46o�o1 CU�ovp^5�o� ����	�h*�p^6�c�u����������ޏp^7R��)�;�@M�_�q�Џ��p^8� ˟ݟ���%���F��L� lCamera�J��@������ӯ���E~� �!�3��OM�_�q��������y  e��Yz� ��	��-�?�Q���u� �ϙ�俽���������>��e�5i��c�u� �ߙ߽߫�d������ P�)�;�M�_�q��*� <��i��������� )���M�_�q������ ����������<�û�� =Oas��>�� ��*'9K ]f�Q����� ��/�%/7/I/� m//�/�/�/�/n<� �^/?%?7?I?[?m? /�?�?�? ?�?�?�? O!O3O�/<׹��?O �O�O�O�O�O�?�O_ !_lOE_W_i_{_�_�_FOXG9+_�_�_oo (o:o�OKopo�o)_�o��o�o�o�o ��	g�0�oM_q�� �No����o�%� 7�I�[�m�&l�n� �Ə؏���� �� D�V�h��������� ԟ柍�g�ڻ}�2�D� V�h�z���3���¯ԯ ���
��.�@�R��� 3uF�鯞���¿Կ� �����.�@ϋ�d�v� �ϚϬϾ�e�w���U� 
��.�@�R�d�ψ� �߬����������� *���w���v��� �����w�����c� <�N�`�r�����=�w� �-�����*< ��`r�����������   ��1CUgy�������   -/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_�W_i_�  
��(�  �%( 	 y_�_�_�_�_�_ �_o	o+o-o?ouocoЙo�o�o�Z* �Q&�J\ n������o�� �9�(�:�L�^�p� ��������܏� � �$�6�}�Z�l�~�ŏ ����Ɵ؟���C�U� 2�D�V���z������� ¯ԯ���
��c�@� R�d�v�����᯾�п �)���*�<�N�`� �����ϨϺ������ ��&�8��\�n߀� �Ϥ߶���������E� "�4�F��j�|��� ����������e� B�T�f�x��������� ����+�,>P b��������� �(o�^p ������� / G$/6/H/�l/~/�/ �/�/�//�/�/?U/ 2?D?V?h?z?�?�/�`@ �2�?�?�?�3��7�P��!fr�h:\tpgl\�robots\m�20ia\cr35ia.xml�? ;OMO_OqO�O�O�O�O8�O�O�O ���O_ (_:_L_^_p_�_�_�_ �_�_�_�O�_o$o6o HoZolo~o�o�o�o�o �o�_�o 2DV hz������o �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟�ݟ��&� 8�J�\�n��������� ȯߟٯ���"�4�F� X�j�|�������Ŀ־:�8.1 �?@88�?�ֻ �ֿ�3�5�G�iϓ� }ϟ��ϳ�������� 5��A�k�U�wߡ߿���$TPGL_O�UTPUT ;|�!�! ��������,�>�P� b�t��������� ����(�:�L�^�p�Ђ����������23�45678901 ���������" ��BTfx��4������
} $L^p��,> ��� //$/�2/ Z/l/~/�/�/:/�/�/ �/�/? ?�/�/V?h? z?�?�?�?H?�?�?�? 
OO.O�?<OdOvO�O �O�ODOVO�O�O__ *_<_�OJ_r_�_�_�_ �_R_�_�_oo&o8o �_�_no�o�o�o�o�o `o�o�o"4F�o T|����\��}�����0�B�T��e�@������� ( 	 ��Џ�� ����<�*�L�N� `���������ޟ̟� ��8�&�\�J���n� ��������ȯ���"�������*�X�j�F� ����|�¿Կ��C��� ϱ�3�E�#�i�{�� �ϱ�S���������� /ߙ�S�e�߉ߛ�y� ����;�������=� O�-�s���ߩ��]� �������'����]� o������������E� ����5G%W} ������g��� 1�Ug	w� {��=O	//� ?/Q///u/�/��/�/ _/�/�/�/�/)?;?�/ _?q??�?�?�?�?�? G?�?O�?OIO[O9O O�O�?�O�OiO�O�O �O!_3_�O_i_{__��_�_�_�_�_�R�$�TPOFF_LI�M >�op:���mqbN_SV�`  l�jP_MON <6�Sdopop2l��aSTRTCHK' =6�f� b�VTCOMPAT�-h�afVWVAR� >Mm�h1d K�o �oop`b�a_DEFPR�OG %|j%�ROB195_S�ERV	�j_DISPLAY`|n"r�INST_MSK�  t| ^zI�NUGp�odtLCK��|}{QUICKM�EN�dtSCRE��p6��btpscdt�q��b�*�_.�ST�jiR�ACE_CFG �?Mi�d`	��d
?�u�HNL 2@|i����k r͏ߏ���'��9�K�]�w�ITEM� 2A�� �%�$1234567�890����  =�<��П��  !���p��=��c ��^���������� .���R��v�"�H�ί ��Я������*�ֿ ���r�2ϖ�����4� ޿�ϰ���&���J�\� n���@ߤ�d�v��ς� �����4���X��*� ��@�����ߨ�� ������T���x��� ���l��������,� >�P�������FX�� d������:� p"��o�� ���F6HZt ~��N/t/�/��/ / /2/�/V/?(?:? �/F?�/�/�/j?�?? �?�?R?�?v?�?QO�? lO�?�O�OO�O*O|O _`O _�O0_V_h_�O t_�O__�_8_�_
o o�_@o�_�_�_Lodo �_�o�o4o�oXojo3 �oN�or��o�(�s�S�B���z��  h��zq ��C�:y
 P��v�]����UD1�:\�����qR_�GRP 1C��� 	 @Cp ���$��H�6�l�Z��|�����f���˟x���ڕ?�  
� ��<�*�`�N���r� ������ޯ̯��&�`�J�8�Z���	�u������sSCB 2D� ���� �(�:�L�^�pς��|�V_CONFIGG E����}�����ϛ�OUTPU�T F�������6�H�Z�l�~� �ߢߴ���������� ��$�6�H�Z�l�~�� ������������� %�9�K�]�o������� ����������"�5 GYk}���� ���1CU gy������ �	/,?/Q/c/u/ �/�/�/�/�/�/�/? ?(/;?M?_?q?�?�? �?�?�?�?�?OO$? 7OIO[OmOO�O�O�O �O�O�O�O_ O2OE_ W_i_{_�_�_�_�_�_ �_�_oo._AoSoeo wo�o�o�o�o�o�o�o ������!�bt �������� �(�:�-o^�p����� ����ʏ܏� ��$� 6�G�Z�l�~������� Ɵ؟���� �2�D� U�h�z�������¯ԯ ���
��.�@�Q�d� v���������п��� ��*�<�M�`�rτ� �ϨϺ��������� &�8�J�[�n߀ߒߤ� �����������"�4� F�W�j�|������ ��������0�B�S� f�x������������� ��,>Pa�t ��������(:L/x���k}gV�K ���//&/8/J/ \/n/�/�/�/W�/�/ �/�/??1?C?U?g? y?�?�?�?`�?�?�? 	OO-O?OQOcOuO�O �O�O�?�O�O�O__ )_;_M___q_�_�_�_ �O�O�_�_oo%o7o Io[omoo�o�o�o�_ �o�o�o!3EW i{����o�� ���/�A�S�e�w� ������������ �+�=�O�a�s����� ����̏ߟ���'� 9�K�]�o��������� ȟۯ����#�5�G��Y�k�}�������ž��$TX_SCRE�EN 1G�g�}i�pnl/��gen.htmſ�*�<��N�`ϽPan�el setupd�}�dϥϷ����������ω�6�H�Z� l�~ߐ�ߴ�+����� ��� �2�߻�h�z� ������9�g�]�
� �.�@�R�d������ ����������}��� <N`r��; 1��&8� \��������QȾUALRM_�MSG ?��� �Ȫ-/?/p/ c/�/�/�/�/�/�/�/�??6?)?Z?%SEoV  -�6�"ECFG Iv��  ȥ�@�  A�1  w B�Ȥ
 [? ϣ��?OO%O7OIO�[OmOO�O�O�G�1G�RP 2J�; 0Ȧ	 �?�O �I_BBL_NO�TE K�:T?��lϢ��ѡ�0RDEFP�RO %+ (%N?u_Ѡc_�_�_�_ �_�_�_o�_o>o)o�boMo�o\INUSER  R]�O�o�I_MENHIS�T 1L�9  �( _P��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1`�oCUgy�)
13/�������*p381,2A3�L�^�p��'��~71�̏ޏ�����0���uedit~(rROB195t0RV��Y�k�}��|o ����ҟ������,� >�P�b�t�������� ί����9Rq�� B�T�f�x��������� ҿ����ϩ�>�P� b�tφϘ�'�9����� ����(߷�L�^�p� �ߔߦ�5������� � �$����Z�l�~�� ���C�������� � 2��/�h�z������� ��������
.@ ��dv����� _�*<N� r�����[� //&/8/J/\/��/ �/�/�/�/�/i/�/? "?4?F?X?C�U��?�? �?�?�?�?�/OO0O BOTOfO�?�O�O�O�O �O�O�O�O_,_>_P_ b_t__�_�_�_�_�_ �_�_o(o:oLo^opo �oo�o�o�o�o�o  �o$6HZl~i? {?������ 2�D�V�h�z����-� ԏ���
����@� R�d�v�����)���П ���������N�`� r�������7�̯ޯ� ��&���J�\�n�����������$UI�_PANEDAT�A 1N����ڱ  	��}/frh�/cgtp/si�ngldev.stm���&�8�J�Y�)priρ�@�}�ϩϻ�������� )�)��M�4�q� ��jߧߎ�����������%�7��[�7����q}��#�flextree���?_fontsize=14e�����x����j�dual��"����i��%�]� o�������������� ��#
G.k} d������n�ܳ��<N`r ��������/ /&/8/�\/n/U/�/ y/�/�/�/�/�/?�/ 4?F?-?j?Q?�?�?s� �?�?�?OO%O 7O�?[O�O�O�O�O �O�O@O�O_�O3__ W_>_i_�_t_�_�_�_ �_�_o�_/oAo�?�? wo�o�o�o�o�o$o�o hO+=Oas�o �������� '��K�]�D���h��� ����ۏNo`o�#�5� G�Y�k�������ş ן�������C�*� g�y�`�������ӯ�� ��ޯ��-�Q�8�u� �������Ͽ��� �j�;Ϯ�_�qσϕ� �Ϲ� ���������� 7��I�m�Tߑ�xߵ� �߮������!�� W�i�{������� H�����/�A�S��� e���p����������� ��+=$aH� �~�.�@���� "4FX)�} ��l�����/ j'//K/2/D/�/h/ �/�/�/�/�/�/�/#?�5??Y?��C�=��$�UI_POSTY�PE  C�� 	 e?��?�2QUICKM_EN  �;�?��?�0RESTOR�E 1OC�  �L?B��6OCC1O��maO �O�O�O�O�OuO�O_ _,_>_�Ob_t_�_�_ �_UO�_�_�_M_o(o :oLo^oo�o�o�o�o �o�oo $6H �_Ugy�o��� ��� �2�D�V�h� �������ԏ�� ��w�)�R�d�v��� ��=���П������ *�<�N�`�r����� ���ޯ���&�ɯ J�\�n�������G�ȿ�ڿ�����7SCR�E�0?�=�u1sc+@u2�K�3K�4K�5K�6�K�7K�8K��2UScER-�2�D�ksMê��3��4��5��6ʬ�7��8���0ND�O_CFG P�;� ��0PDAT�E ����None�2��_I�NFO 1QC�@��10%�[���I� ��m߮��ߣ������� ���>�P�3�t��i�����<-�OFFSE/T T�=�ﲳ $@������1�^�U� g�������������� ��$-ZQcu����?�
����U�FRAME  ���*�RTOL_ABRT	(�!�ENB*GRP� 1UI�1Cz  A��~��~ ���������0UJ�9MS�K  M@�;N%8�%��/�2oVCCM��V��V�#RG�#Y�9����/����D�BH��p71C����3711?�C0�$MRf2_�*S�Ҵ��	���~XC�56 *�?�6����1$�5���A�@3C��. ��8�?��OOKOx1FOsO�5�51���_O�O�� B����A2�DWO�O 7O_�O8_#_\_G_�_ k_}_�__�_�_�_�_�"o�OFoXo�%TCC��#`mI1�i������� GFS��2�aZ; �| 23�45678901 �o�b�����o�� !5a�4BwB�`56� 311:�o=L�Br5v1�1~1�2�� }/��o�a��#� GYk}�p��� ����ُ�1�C�U� 6�H���5�~���ߏ����	���4�dSEL#EC)M!v1b3��VIRTSYNC��� ���%�SI?ONTMOU�������F��#b�����(u FR:\H��\�A\�� �߀ MC��LO�G��   UD�1��EX����'� B@ �����̡m��̡  O�BCL�1�H� ��  =	 �1- n6  G-������[�,S�<A�`=��͗���ˢ��TRAIAN⯞b�a1l�
0�d�$j�T2cZ; (aE2ϖ�i��;� )�_�M�g�qσϕϧπ�������	��F�S?TAT dm~2!@�zߌ�*j$i߾߮�_GE�#eZ;��`0�
� 02���HOMIN� f������ P~�����БC�g�X����JMPERR {2gZ;
  �� *jl�V�7�������� ������
��2�@�q�hd�v�B�_ߠRE� �hWޠ$LEX��i�Z;�a1-e��VM�PHASE  �5��c�!OFFX/�F�P2n�j�0�㜳E1@���0ϒE1!1?s33�����ak/�k�xk䜣!W�m[�� ���[����o3;� [i {����/ �O�?/M/_/q/� �/��//�/'/9/�/ =?7?I?s?�/�?�/�/ �?�??Om?O%O3O EO�?�?�O�?�O�O�? �O�O�O__gO\_�O E_�O�_�O�O/_�_�_ �_oQ_Fou_�_|o�o �_�oo�o�o�o�o;o Mo?qof-�oI� ����7�[ P���������ˏ ��!�3�(�:�i�[��ŏg�}������TD�_FILTEW�n��� �ֲ:��� @���+�=�O�a�s� ��������֯��� ��0�B�T�f�x����SHIFTMENoU 1o[�<��%��ֿ����ڿ�� ��I� �2��V�hώ� �Ϟϰ�������3�
��	LIVE/S�NAP'�vsf�liv��E��^��ION * Ub�h�menu~߃��`���ߣ���p����	����E�.�5T0�s�P�@� ���AɠB8z�z���}��x�~�P��c  ���MEbЩ��<�0���M�O��q���z�W�AITDINEN�D������OK�1�OUT���S�D��TIM����o�G���#���C����b������REL�EASE������T�M�������_A�CT[�����_D?ATA r���%L����xRDI�Sb�E�$XV�R�s���$ZA�BC_GRP 1Ut�Q�,#�0�2���ZIP�u�'�&����[M�PCF_G 1v��Q�0�/� wx�ɤ� 	�>Z/  85�/0�/H/�/l$?��+�/ �/�/?�/�/???r?>�?  �D0�? �?�?�?�?�;����x�]hYLINuD֑y� ��� ,(  *VO�gM.�SO�OwO�O�M i?�O�O^PO1_�O U_<_N_�_�O�_�_�_ _�_�_x_-ooQo8o`�_�o�oY&#2z�� ���oC�e?�a?>N|�oq�����qA�$DSPHE_RE 2{6M��_ �;o���!�io| W�i��_��,��Ï�� �Ώ@��/�v���e� ؏��p���������l�ZZ�� �N