��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SF�TVER����_�GRP6� �2$FS_FOR�C� ��P�S_GMEA2'%� 1G�F#2G0 �GTS_K_CHKY%O �RIc"]!APP��$PS_AA�ML��$�"�	]$/!_MI2�$AS�!!�#'#�#�!��3  2 RO�M_RU2$Jn� EST2!$� ��N_NU�$�u �  
$SBn*BSCNCTO�INS29FS� _�NG$GAG�Ex� � CUToFREQY#LR*�REAL%� �2M�OMEN�T�V�C�F�C��2N�C�K1DT��1D�EVIDS�7 {	�3PATH�0]A�3FNA� 6!�	AEX� �5O �8BUF�7TDP�Y�FLGEJ5�� � � N IU�
@!(UF*����4OS/� ��DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� !�ARE-  ? � �0�BB{F S{T� M�D|TRS$STD6XlQCWFA� 7X�QCW��"YV�"eS/ �A7 �  $�@TI�Nd@�0SULگ �R_@ g $}@ SW�@�RO�RR%	� �P�T� �@J�U� �SqFS4DN6
 �2P�0_@�cFOL[d!$�FIL� jjE�P��C�S�aDIG4R_C_SCA��c�INTTHRS�_BIdA�dSMA9L�bCOL�b9G�`� �� ��_IVTIM��$!0B"$S�?0xCCBDDN���-qI2wT2wDE�BUdA\!SCHN�"TOfa0�! �  Q0mr<0V� �;!�r~AUTTUN�� TRQa�uE�40N �qFS3A	XG  � 1eb}tj�rI�v,	"G_gr>7 l �!�3>@WEIGH�q�2� uS_5QF(�T�2�WA� 	pEsNTERVA�; -  Q�� S!�t�AS0S��$J-_STAF�p JQg���1(�U��2��3��W����� hqx��"COG+_X�Y�Z�ҁCM�p?�p�܂RSLT�4��D��D��	"_�p_�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDBH	"I%�0 ,$M"Pp30f��� d��:pG p"��HCDv�GV�#GVY��Z�JDO5�,q���S��$R��E_�8@{٣�pAP�HBC��$VF6�P��2L��蘨@IL[����;����;�d@���RG���NGEW_���r�Q}�8��ڡ�5OBOA@fQY�sW2/�G<�	����ȴ\�2�E�KP��NUCNPRGOVp����@`d_TW�cj,�G�E^!NV2#�C�c0@�WTS�T�RL_SKI2!�$SJ�Q��NQpG�W���q��7 o\ ;0FR]b3� � CMDC��`�T�b���TO?@��� �5گ���_�A�h 0 '��ALARqM�_�*�TOT6�GFRZn l�,!Y 3 ��X!��mӥ�X �Œ`�X �ʕ�U#��2��2p
�X#Z���FIX�8"��F�"��IT�`�IB�PN_d��CH8�%��_DFL _�GBF2N�ڶ�3����� ��3�"���@��ʷ�� ����3���3
��X��DIA ����/#� ���%�����[1��g1� [���Z��#��!���%���$0�@
p��d7F��D�� HA�p�U�5����v�FSI]W6 �2PN@�`R>!�PHMP�`HCK%���>0G�'*#e A����p�NT��^H	��HU�FRzs3��A��U�gvCa�$v0Q O����@p@p3 �  SI0��  �=5�IRTU_��|� %SV 2���   �6>0]@]	Q�EF@ �oP��  @p�  � �//'/9/K/U%*@pd@p
m hK�/ w/�/�/�(��$��/ � �/�/?.8e"�/? J?\?r?8?�?|?�?�? �?�?�?�?>O4ObOO �OTO�O�OjO|O�O�O �O_�O(__\_f_�_ B_�_�_�_�_ o�_$o �_Ho>oo^b�/�ot���%�/�o�o�k	�MC: 5678�  Afsdt�1 789012�34q#5w  �	q 6xz.�Ops�'��j !l�o�o����������,�5�DMM �)5�A ��x�������|=���OR 2	Q� ��m���_� tuB?�)DN�S4D7 
Q�!tY�d�!Ls|�q`rƈ̀[?�l�B𴐠��$ ONFIG ��(�� � 2�����i!��� 2�,
�Hand gui�de��?�3�?��  �X��с쿏ь�g#�=���A��ύ��� ����p�ݯ�(���L�7�p�[����m*������ʿܿ�  ��$�6�H�Z�lɌ� �ό��ϰ���������
�C�E�I 2jQ�(�0� -�hzՀ�Fտ��_`�πB����d�C� y ��uq=#�
_a�Nnk(��K�y���̥@��e���=D����_a;�{���8I��^_aIt$ �$Fݟ>���k"��{�Q�Fۀ3]� ��ѯǯ���!�/�``�+�����.��y���_a$敕��(4$�����>��E��B<~w�%�_a8E�y5�;�jA��Ҝ��Q�>��]�_a? ��m��箑����~u1Џ?�33����0�:�o����0�����LSB��~uq@�ӻ��m�S]�}��8��� ���t�	eF|����]��߯�����n��;ӽ.����3�'	c�����B���4* 2/V��<%D�DH  *%v�+��^-��
�/1��/u/~u�J/l/�)AI��/�/�?/G A��n5��p�� 4vO?;)�7�?�?�o�?�8Jhq�?�?zyj�G�_FSIW Q��9��O�O�Ou�