��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SF�TVER����_�GRP6� �2$FS_FOR�C� ��P�S_GMEA2'%� 1G�F#2G0 �GTS_K_CHKY%O �RIc"]!APP��$PS_AA�ML��$�"�	]$/!_MI2�$AS�!!�#'#�#�!��3  2 RO�M_RU2$Jn� EST2!$� ��N_NU�$�u �  
$SBn*BSCNCTO�INS29FS� _�NG$GAG�Ex� � CUToFREQY#LR*�REAL%� �2M�OMEN�T�V�C�F�C��2N�C�K1DT��1D�EVIDS�7 {	�3PATH�0]A�3FNA� 6!�	AEX� �5O �8BUF�7TDP�Y�FLGEJ5�� � � N IU�
@!(UF*����4OS!	 D�MM�A@  �@ $�AbERE�G_OF�B�BME��HAS�C1�A ��DRE-  � � �0�B{F S{T� M�DTRS$STD6XlQCWFA� 7X�QCW�"YV�"eS/ �A7  w $�@TINd@��0SUL� ��R_@  $}@ SW@�R�O�RR%	 h�P�T� �@JU� z�SO/ FS4D6'
 �2P�0_@c�FOL[d!$FCIL� jjE�P��C�S�aDIG4RC�_SCA��cI�NTTHRS_�BIdA�dSMAL��bCOL�bG��`� �� ��_�IVTIM�$t!0B"$S?0~xCCBDDN���-qI2wT2wDEByUdA\!SCHN�"TOfa0�! � Q0 mr<0V� �;!�r�AUTTUNN� TRQa�uE40�N �qFS3AXG  � 1eb}t�r5I�v	"G_gr7 l �!�3@�WEIGH�q�2 UuS_5QF(�T2��WA� 	pEsNTERVA�; - Q��� S!�t�AS0S�{$J-_STA�p� JQg���1(�*��2��3��W���� hqx��"COG_�X�Y�Z�ҁCM�p?�p�܂RSLT�4��D�P�D��	"_�p_�q�7  �~�b#0V�ROUNDCMVP�ERIODA�1P�UU3F2D�'TM01� �Ƒ_D���GAMMc1�TWRXI�K�K�MK��CLbP�&O00�ADJ�GAu�U�PDB#I%0/ ,$M"P30f��� d�:pG �p"��HCD�G]V�#GVY��Z�GJDO5�,q��S��7$R��E_8@{t٣�pAPHBCy��$VF6��P��2L��蘨@IL [����;���;�d@���RG���NEW_���r�Q}���ڡN�5OBOA@fY�sW2/�G<�	����ȴ�\�2�E�KP�NUC?NPRGOV��Ŝ�@`d_TW�c,�G�E^!NV2#C�c0�@�WTS�TRL�_SKI2!$SiJ�Q��NQpGW���	"��7 \ m;0FR]b� � CMDC���T�b���TO?��� �5گ���_�Ah 0 '�>�ALARM�_��*�TOT6�FRZn l�,!Y 3��X!�� mӥ�X �Œ`X �ʕ�U#��2��2
�X#Z�N��FIX�8��F�"d��IT�`IB�PN_d��CH�%���_DFL _�BF2N�ڶ�3����� ��3�"�����ʷ�(� ����3��3
��X��DIA����/#� ���%��� ��[1��g1�[���Z���#��!���%����$0�@
p��7F��D,�� HA�pU�5����v�FSIW6K �2PN@�`R>!��PHMP�`HCK%���>0G�'*#eb A����pNT��p^H	��HUFRzs�3��A��UgvM���$v0Q ��i��@p@p � � SI0��  �5�I�RTU_��� %S�V 2���  � �6>0]@�]	Q�EF@� �oP�  �p�p � �/@/'/9/K/U%@pd@p
m hK�/w/�/�/ �(��$��/� �/�/ ?.8e"�/?J?\?r? 8?�?|?�?�?�?�?�? �?>O4ObOO�OTO�O �OjO|O�O�O�O_�O (__\_f_�_B_�_�_ �_�_ o�_$o�_Ho>o o^b�/�ot��%�/�o��o�k	MC:� 5678  A�fsdt1 78901234qx#5w  	q 6xz.Ops�1'O�O��h l�o�o����������,�5�DMM c�)5�A ���x�������=���O�R 2	Q� "��m��_� tu�B?)D�N�S4D 
FQ�!tY�d�!Ls`|�q`rƈ̀?�l��B𴐠�$ ON�FIG �}(�[ � ������i!�� 2��,
Hand guide���?�3��� � �X��с��ь��g#�=���A��ύ�������p �ݯ�(��L�7�p�x[����m*�� ����ʿܿ� ��$� 6�H�Z�lɌ��ό��� ���������
�C�E�]I 2Q�(�0� -�zՀ�F�M���_`πB��<��d�C�  ��#��=#�
_aNnk=(��K����̥�@��e��=D�y���_a;�����8I��_aIt�$ �$F�>�s��k"���Q�Fۀ3]儢ѯǯ����!�/�``+��=���.�����_a�$敕��(4$������>�E���B<~w%�_a8�E�y5�;�j�A��Ҝ�Q�>��]�_a?��m���஑����~u1�?�3�3����0�:�o ����0�����LSB��~uq�ӻ���m�S]���/8��� ��� t�	eF|���P]��߯���x�n��;�.��z��3�'	���,��B���4*� 2/V��%D�DGH  *%v�+� �^-��
�/��/u/F~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?�;)�7�?�?�o�?�8J�hq�?�?zyjG�_F?SIW Q��9 ��O�O�Ou�