��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER��q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OSu?  �DMM�A@�  @ $��AbEREG_OFl�B�BME�HAS�C�1�A �DRE�-   � �0�B{F S{T� �M�DTRS$ST1D6XlQCWFA� 7X �QCW�"YV�"eS/ �A~7   $�@�TINd@�0SkUL� �R_@�  $}@ S�W@�RO�RR�%	 �P�T� Ɔ@JU� �SqFS;4D6
 �2P�0�_@cFOL[d!$FIL� jjEʄP�C�S�aDI~G4RC_SCA���cINTTH�RS_BIdA�dS�MAL�bCOL��bG�`� �� ��_IVTIM��$!0B"�$S?0xCCBDSDN��-qI2wT2w�DEBUdA\!SCHN�"TOfa0�!  � Q0mr<0V� ��;!�rAUTTUuN� TRQaʤuE40N �qFS'3AXG  � 1eb}t�rI�v �bgr>7 l �!�3>@WEIGH�q�2� uS_5QF(�T�2�WA� 	pEsNTERVA�; -  Q�� S!�t�AS0S��$J-_STAF�p JQg���1(�U��2��3��W����� hqx��"COG+_X�Y�Z�ҁCM�p?�p�܂RSLT�4��D��D���r_�p_�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDB�rI%�0 ,$M"Pp30f��� d��:pG p"��HCDv�GV�#GVY��Z�JDO5�,q���S��$R��E_�8@{٣�pAP�HBC��$VF6�P��2L��蘨@IL[����;����;�d@���RG���NGEW_���r�Q}�8��ڡ�5OBOA@fQY�sW2/�G<�	����ȴ\�2�E�KP��NUCNPRGOVp����@`d_TW�cj,�G�E^!NV2#�C�c0@�WTS�T�RL_SKI2!�$SJ�Q��NQpG�W���r��7 �\ ;0FR]b� � CMDC���T0�b���TO?�� � �5گ���_�Ah �0 '��ALARM��_�*�TOT6�F#RZn l�,!Y 3�� X!��mӥ�X �Œ`X P�ʕ�U#��2��2
�8X#Z���FIX�8�ґF�"��IT�`IeB�PN_d��CH��%��_DFL _�B#F2N�ڶ�3����� ��3�"�����ʷ�� ����3��3p
��X��DIA����/#� ���%�����[1��g1�[� ��Z��#��!���%���$0�@
p��7F���D�� HA�pU��5����v�FSIW.6 �2PN@�`uR>!�PHMP�`HCK%���>0G�'�*#e A����pN�T��^H	��HUFARzs3��A��Ugv�Ca�$v0Q ����@p�p� � � SI0��P��5�IRT�U_��� %SV �2��   ��P4>0]@]	Q<�EF@ �o|P�  @pP�� �//'/9/�K/U%@pd@p
m h K�/w/�/�/�(��$ ��/� �/�/?.8e" �/?J?\?r?8?�?|? �?�?�?�?�?�?>O4O bOO�OTO�O�OjO|O �O�O�O_�O(__\_ f_�_B_�_�_�_�_ o �_$o�_Ho>oo^b�/��ot��%�/�o�o�k�	MC: 56�78  Afs�dt1 78901234q#5w� ��	q 6xz.�Ops�'��j !l�o�o����������,�5�DMM �)5�A ��x�������|=���OR 2	Q� ��m���_� tuB?�)DN�S4D7 
Q�!tY�d�!Ls|�q`rƈ̀[?�l�B𴐠��$ ONFIG ��(�P� � 2�����i!��� 2�,
�Hand gui�de��?�3�?��  �X��с쿏ь�g#�=���A��ύ��� ����p�ݯ�(���L�7�p�[����m*������ʿܿ�  ��$�6�H�Z�lɌ� �ό��ϰ���������
�C�E�I 2jQ�(�0� -�hzՀ�Fտ��_`�πB����d�C� y ��uq=#�
_a�Nnk(��K�y���̥@��e���=D����_a;�{���8I��^_aIt$ �$Fݟ>���k"��{�Q�Fۀ3]� ��ѯǯ���!�/�``�+�����.��y���_a$敕��(4$�����>��E��B<~w�%�_a8E�y5�;�jA��Ҝ��Q�>��]�_a? ��m��箑����~u1Џ?�33����0�:�o����0�����LSB��~uq@�ӻ��m�S]�}��8��� ���t�	eF|����]��߯�����n��;ӽ.����3�'	c�����B���4* 2/V��<%D�DH  *%v�+��^-��
�/1��/u/~u�J/l/�)AI��/�/�?/G A��n5��p�� 4vO?;)�7�?�?�o�?�8Jhq�?�?zyj�G�_FSIW Q��9��O�O�Ou�