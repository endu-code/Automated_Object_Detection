��   �A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����CCSCB3�_GRP_T �  � $FS�_TYP3  �$PS_SBF�RAME3��$�J  $INIT_TOL^�RANGE3_F�_uT~FTR/ATIO^c ��P_H_LIMA��L�FSOF�ST_S^JM3�_f _ �$$�CLASS  O������[���[� VERSIO�N�  ��5IRTU�AL��' 2 [� 6 � � �����b@� � B ��B A�x���Cp  ��� Y��B�z��m