��   P�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����PM_CFG�_T   � �$NU( HNL�  $IOD�_KEEP?ER�R_SEV?DE_V_FLG?CG	�CT
SCAN_M�ULT?CH1_wENB>CH2��SPARE1�2�3�e�   G ��i�2����  &ST�AT- \ �$BD$?UPD�ATE_FW?P�MTK_DBGL�V>PMUIQE�XPE_VERS�? $CURp ��$$CLASS  �������b��b�tIO�N�  ��5�IRTU�AL��'/ �bw � � � //0/B/ T/f/x/ 
 ���/�/ �/�/�/�// ?2?D? V?h?z?�/�?�?�?�?`�?�?���6����:@