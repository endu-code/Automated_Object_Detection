��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SF�TVER����_�GRP6� �2$FS_FOR�C� ��P�S_GMEA2'%� 1G�F#2G0 �GTS_K_CHKY%O �RIc"]!APP��$PS_AA�ML��$�"�	]$/!_MI2�$AS�!!�#'#�#�!��3  2 RO�M_RU2$Jn� EST2!$� ��N_NU�$�u �  
$SBn*BSCNCTO�INS29FS� _�NG$GAG�Ex� � CUToFREQY#LR*�REAL%� �2M�OMEN�T�V�C�F�C��2N�C�K1DT��1D�EVIDS�7 {	�3PATH�0]A�3FNA� 6!�	AEX� �5O �8BUF�7TDP�Y�FLGEJ5�� � � N IU�
@!(UF*����4OS^� ��DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�Ag 	 �ARE-   � �0��B{F S{T� M��DTRS$STD6XlQCWFA� 7X�Q CW�"YV�"eS/ �A7 �  $�@T�INd@�0SU�L� �R_@ � $}@ SWP@�RO�RR%G	 �P�T� �@�JU� �SqFS4�D6
 �2P�0_�@cFOL[d!$FIL� jjE�eP�C�S�aDIG4�RC_SCA��cINTTHR�S_BIdA�dSMsAL�bCOL�rbG�`� �� v��_IVTIM��$!0B"$�S?0xCCBDD�N��-qI2wT2wD�EBUdA\!SCHN�"TOfa0�!  � Q0mr<0V� �;!��rAUTTUN:� TRQa�u�E40N �qFS3AXG  � 1eb�}t�rI�v	"G_|gr7 l �!|�3@WEIGH�qV�2 uS_5QF(�MT2�WA� 	pEs?NTERVA�; @- Q�� S!�t�AS0�S�$J-_ST�A�p JQg���1�(���2��3��W����� hqx��"COWG_X�Y�Z�6ҁCM�p?�p<�܂RSLT�4�@�D��D��	"_�p9_�q7  �~�b#�0VROUNDCM?VPERIODA�w1PUU3F2D�'�TM1� �Ƒ_D<��GAMMc1^�TRXI�K�5K�K��CLbP�&�O00ADJ�GAVu�UPDBh	"I%0 ,$M"�P30f��� �d�:pG p"��HC�D�GV�#GVY:��Z�JDO5�,q���S��$R��E�_8@{٣�pA�PHBC��$#VF6�P��2L����@IL[����;� ��;�d@���RG����NEW_���r�Qp}���ڡ�5OBOA@�fY�sW2/�G<�	 ����ȴ\�2�E�KP��NUCNPRGO�V����@`d_TWԔc,�G�E^!NV02#C�c0@�WTS�TRL_SKI2!O$SJ�Q��NQp�GW��	"��7 o\ ;0FR]b3� � CMDC��`�T�b���TO?@��� �5گ���_�A�h 0 '��ALARqM�_�*�TOT6�GFRZn l�,!Y 3 ��X!��mӥ�X �Œ`�X �ʕ�U#��2��2p
�X#Z���FIX�8"��F�"��IT�`�IB�PN_d��CH8�%��_DFL _�GBF2N�ڶ�3����� ��3�"���@��ʷ�� ����3���3
��X��DIA ����/#� ���%�����[1��g1� [���Z��#��!���%���$0�@
p��d7F��D�� HA�p�U�5����v�FSI]W6 �2PN@�`R>!�PHMP�`HCK%���>0G�'*#e A����p�NT��^H	��HU�FRzs3��A��U�gvCa�$v0Q O����@p@p3 �  SI0��  �=5�IRTU_��|� %SV 2���   �6>0]@]	Q�EF@ �oP��  @p�  � �//'/9/K/U%
@pd@p
m P�M� y/�/�/�&��$��/ � �/�/?.8e"�/? J?\?r?8?�?|?�?�? �?�?�?�?>O4ObOO �OTO�O�OjO|O�O�O �O_�O(__\_f_�_ B_�_�_�_�_ o�_$o �_Ho>oo^b�/�ot���%�/�o�o�k	�MC: 5678�  Afsdt�1 789012�34q#5w  �	q 6xz.�Ops�'��j !l�o�o����������,�5�DMM �)5�A ��x�������|=���OR 2	Q� ��m���_� tuB?�)DN�S4D7 
Q�!tY�d�!Ls|�q`rƈ̀[?�l�B𴐠��$ ONFIG ��(�� � 2�����i!��� 2�,
�Hand gui�de��?�3�?��  �X��с쿏ь�g#�=���A��ύ��� ����p�ݯ�(���L�7�p�[����m*������ʿܿ�  ��$�6�H�Z�lɌ� �ό��ϰ���������
�C�E�I 2jQ�(�0� -�hzՀ�Fտ��_`�πB����d�C� y ��uq=#�
_a�Nnk(��K�y���̥@��e���=D����_a;�{���8I��^_aIt$ �$Fݟ>���k"��{�Q�Fۀ3]� ��ѯǯ���!�/�``�+�����.��y���_a$敕��(4$�����>��E��B<~w�%�_a8E�y5�;�jA��Ҝ��Q�>��]�_a? ��m��箑����~u1Џ?�33����0�:�o����0�����LSB��~uq@�ӻ��m�S]�}��8��� ���t�	eF|����]��߯�����n��;ӽ.����3�'	c�����B���4* 2/V��<%D�DH  *%v�+��^-��
�/1��/u/~u�J/l/�)AI��/�/�?/G A��n5��p�� 4vO?;)�7�?�?�o�?�8Jhq�?�?zyj�G�_FSIW Q��9��O�O�Ou�