��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP������8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGDsEV��RCM+ ;$Z <��QSIZ�X|�� TATUSW�MAILSERV~ $PLAN� �<$LIN<�$CLU���<${TO�P$CC�&sFR�&�JEC�!}�%ENB � �ALARl!B�TQP�3�V8 S��_$VAR9M �ON
6��
6APPL
6PA� 5B 	7'POR��#_�!�"�ALERT�&�2U�RL }�3A�TTAC��0ER�R_THRO�3UaS�9z!�800CH- �Y�4MAXNS_�1�AMOD4�AI� $B� �(APWD  �� LA �0�ND�ATRYQFDEL�A_C@y'>AERS�I�A�'ROtIC�LK�HMR0�'� X�ML+ :3SGFReM�3T� XOU�3�PING_�_COAPA1�Fe3�A�'C�25�B_AU�� k �6R,2COU�!H!U�MMY1RW2?��RDM*� $�DIS�� SMeB�	"�BCJ@b"CI2AIP�6EXPS�!�P�ARQ$�RCL��
 <(C�0�S�PTM�E� PWR���X�V�RoC l5��!�"%�7�ICC�%� kf�R�0leP� _DLIV��YNo3 �<oNbX_�P~#Z�_INDE
C�`O�FF� ~UR�iD���c�   �t �!�`MON��%sD�&rHOU�#EWA,vSq;vSqJv�LOCA� Y$�N�0H_HE����@I"/ 3 �$ARPz&�1FF�W_\ �I!F�`�;FA�Dk01#�H{O_� INFO�s;EL	% P K � !k0WO` $ACCE� �LVZk�2H#IcCE�L��P�$�s�# ���k���
���
`�K`SQi���P�5|�I�0ALh�z�'0 ��+
���F����P��܅�$� 2ċT"�w��� ���� č��!r�Z����4���Ċ!�147.87.2�24.20h�S���96����܁܁3�u_{p_  ċ�� bfh.ch̟�1�C�U�g�y����������ӯ^�� _?FLTR  ��πW �������!�n�nxč2n��r{SH�PD 1ĉ�  P!
r�obstatio�n֯՚!k�. �Q�ſ�������� ޿?��c�&χ�Jϫ� �π��Ϥ����)��� M��"߃�Fߧ�j��� ���߲���%���I�� m�0��T��x���� �����3���W��{� ��P���t��������� ����Sw:� ^������@= a$Zׯ$ �_L�A1��x!�1.�ğP�1|�Q255.%L�S���2���E �//*/<&3 F/�� l/~/�/�/<&4�/�50�/�/??<&56?��0\?n?�?�?<&6�?�%@�?�?��?
O1�?P��M�Y� MY���c��� 'Q� �VN<�O�O _�O+_=_O_"_s_�_NPd_�_�_�_�_�_ o!o3o�_Woio{oVNLoM��o�l�oAo�
.@U}i�RConnect�: irc\t//?alertsE� ���Pu���P�1�C�UуP_R8�d��H�~����� ��Ə؏���� �2��D�V�S$���8�( p����o͟ߟ��QIA8��d�A�B 4��j�h9�Q+��@7DM_�A+��?SMB 	X�8%�ğVO��߯���_C�LNT 2
X� 4C�ɯ0��l� c�B�T���x���Ͽ�� ����)�;��_�q��Pϕ��MTP_C�TRL ��% ���ϙdc���ߋ�� ?�*�c߳l��N���@C{�Vߵ�Ƥ��������ѓC��USTOM {�2��}�@ }�D_TCPIPu�{�q�h�E�TEL��{��A���H!�Ta�t�çrooblolr�  �~��!KCL�����F��!CR�T��������!CONS&����	n+���