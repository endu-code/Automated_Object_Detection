��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�#J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA R�!R�	� � $TIT�!$I��N �D@d�Dd �Dc@�D5�FU6�F7�F8�F9�G0�G�GJA�E�GbA�E
�G1�G1�G �F�G�2�B!SBN_C�F>"
 8F CN�V_J� ; �"�!_�CMNT�$F�LAGS]�CH�EC�8 � ELL�SETUP ރ $HO30IO��0� %�SMAC{RO�RREPR�X� D+�0��R{�T� UTOBACK�U�0 ��)DEVIC�CT	I*0�� �0�#��`B�S$INTE�RVALO#ISP�_UNI�O`_D�O>f7uiFR_F�0AIN�1���1<c�C_WAkda^�jOFF_O0N�DEL�hL� ?aA�a1b?9a�`C#?��P�1E��#s�ATB�d��MO<� �cE D [�M�c��^qREV��BILrw!XI�� QrR  �� OD�P�q�$NO^PM�#  �s�r/"�w@� �u�q�r�0D`S� p E R�D_E�pCq$F�SSBn&$CHK�BD_SE^eAG� G�"$SLOCT_��2=�� V�d¾%��3 a_E�DIm   �S �"��PS�`�(4%$EP�1�1'$OP�0�2�a�p�_OK�UST1P_C� ��d��U �P/LACI4!�Q�x4�( raCOMM� ,0$D����0�`���EOWBn�IGALwLOW� (Kt�"(2�0VARa�Є@�2ao�L�0OUy� ,Kvay��P9S�`�0M_O]�����CCFS_UT~p0 "�1�3�#�ؗ`X"�}R0 � 4F IMCM�`O#S�`��upi R�_�p�BA�!t���M/ h�pIMPEE_F� N��N���@O��r��D_�~�n�Dy�F� dCC_�r0 � T� '��'�DAI�n0"��p�P�$I�������F�t X� G�RP0��M=qNF�LI�7��0UIR�E��$g"� SWI�TCH5�AX_N��PSs"CF_LI�M� � �0EED��!��qP��t�`PJ_dVЦMODEh�.Z`�PӺ>�ELBOF� � �����p� ���3���� FB/��0��>�G� �� WOARNM�`/���qP��n�NST� C�OR-0bFLT�Rh�TRAT�PT|1�� $ACC1a��N ��r$OR�I�o"V�RT�P_�S� CHG�0I���rT2��1�I���T�I1��� x i#�Q��HDRBJ; CQ�U2L�3L�4L�5L�E6L�7L� N�9s!���O`S <�F +�=�O��#92��L�LECy�"MULTI�b�"N��1�!t���0T�� �STY�"�R`�=l��)2`����*�`T  |� �&$��۱m�a�P�̱�UTO��:�E��EXT����pÁB���"2� (䈴![0������p<�b+�� "D" ���ŽQ��<煰kc!(�9�#���1��ÂqM�ԽP��" '��3�$ L� E���P<��`A�$JO�Bn�T���l�TRIG3�% dK����� ��<���\��+�Y����_M��& tf�pFLܐBNG AgTBA� ���M� �
�!��p� �q��0��P[`��O�'[���0tna*���"MJ��_R���CDQJ��IdJk�D�%�C�`�Z���0��Pq_�P��@ ( @F �RO.��&�t�IT�c�NOM�
��T��Sp�P`T)w@���Z�P�d���RA�0��2b"�����
$T����MD3�T��`U31���pe(5!HGb�T1�*	E�7�c�KAb�WA8b�cA4#YNT����PDBGD�� *(��PUt@X�܌W���AX��a��eT;AI^cBUF��|0!+ � 7�n�PIW�*5 P��7M�8M�9
0�6F>�7SIMQS@>wKEE�3PATn��^�a" 2`#�"�L6�4FIX!, ���!d��D�2Bus=CsCI�:FPCH�P:BAD�aHCEhAOG�hA]HW�_�0>�0_ h@�f�Ak���F�q\'�M`#�"�IE3�- l�p3G��@FSOES]FgHBSU�IBS�9WC��. ` ��MARG쀳���FACLp�SLEWxQe�ӿ���MC�/�\pSM_JBM����QYC�	g�e#��0� ā�CHN-�MP�$G� Jg��_� #��1_FP$�!TCuf!õ#�� ���d�#a��V&��r��a;�fJR���rSoEGFR�PIO�^ STRT��N���cPV5���!41 �r��
r>İ�b�B�~O�2` +� [���,qE`&�,q`y��Ԣ}t��yaSIZ%���t�vT�s� �z|�y,qRSINF} Oбc���k��`��`��`L�ĸ T`7�CRCf�ԣCC/�9��`�a�uah�ub'�MIN@��uaDs�#�G�D�YC��C�����e�q0���� �EV�q�F*�_�eF��N3�s�Pah��Xa+p,5!��#1�!VSCA$?� A��s1�"!3 ��`F/k��_�U ��g��]��C�� a�s��.bR�4� @����N����5a�R��HANC��$LG؆�P�f1$+@ND,P�t�AR5@N^��a0�q���c��ME�18����}0��RAө�A�Z 𨵰�%O��F�CTK��s`"�S\�PFADIJ�OJ� ʠ�ʠ���<���Րļ�GI�p�BM�P�d�p�Dba��AE�S�@	�K�W_��B�AS�� �G�5 � M�I�T�CS�X[@@�!62�	$�X���T9�{sC➠N�`�a~P_HE�IGHs1;�WIDl�0�aVT ACϰ��1A�Pl�<���E�XPg���|��CU��0MMENU��7n�TIT,AE�%)�a2��a��8� P� a�ED�E�  ��PDT��R�EM.��AUTH?_KEY  ������ �b�O	ь}1�ERRLH� �9 1\� �q-�OR�DB��_ID�@l �PUN�_O��Y�$SY�S0��4g�-�I��E�EV�#q'�PX�WO�� �: $CSK7!f2��(�Td�wTRL��; �'�AC�`��ĠIND&9DJ.D��_��f1���f���PL�AF�RWAj���SD�A���A+r|��UMgMY9d�F�10d��&���J�<��}1PR�� 
3�POS���J�= �M$V$�q�PL~�!>���SܠK�?�����CJ�@����ENE�@T��A���S_��RECOR��B�H 5 O�@=$LA�>$~�r2�`R��`�q�b`�_Du�&�0RO�@�aT[�Q� �b������! }У��PAUS���dETgURN��MR�U�  CRp�EWyM�b�AGNAL:�s2$LA�!�?$PX�@$P��y A �Ax�C0 #ܠDO�`X�k��W�v�q�GO_AWAY��MO�ae����]�CSS_CCwSCB C �'N��CERI��гJ`u�QA0�}�\�@�GAG� R�0��`��{`��{`O�F�q�5��#M5A��X���&ш�LL�D� �$���sU�D)E%!`|���OVR10W��,�OR|�'�$E�SC_$`�eDSB#IOQ��l ��B.�VIB&� �c,������f�=pSSW����f!VL��PL|���ARMLO
���`����d7%SC� �bALspH�MPCh �Ch �#h �#
h 5�UU���C�'��C�'�#�$'�d�#C \4�$�pH��Ou��!Y��!�SB���` k$4�C�P3Wұ46�$VOLT37$$`�*�^1���$`O1*�$o��0R�QY��2b4�0DH_THE����0S�<�4�7ALPH�4�`����7�@ �0�qb7
�rR�5�88� ×@���"��Fn�	MӁVHBPFUAF�LQ"D�s�`�THR��i2dB�����G
(��PVP�����������1�J2�B�E�C�E�CPSu�Y@��F b3���H�(V�H:U�G��
X0��FkQw�[�N�a�'B���C INH=BcFILT��� $��W�2�T1�[ @��$���H YАAF�sDO��Y�R p� fg�Q�+�c5h`�Q�iSh�QPL��x�Wqi�QTMOU�# c�i�Q\��X�gmb��Hvi�h�bAi�fI�aCHIG��ca	xO��hܰ��W�"vAN-uX!��	#AV�H!Pa8$P�ד#p�RE_:�A�a��B�qN0�X�MCN�0��f1[1�qVE�p��Z2;&f�I�QO�u�r�x�wGldDN{G|d��aF>!�9��a9M:�U�FWA�:�Ml���X�Lu��$!����!l�ZO����0%�O�lF�s�13�DI�W�@��Q����_��!CURVAL԰0rCR41ͰZ�C <�r�H�v���<�`��<�(�f�CH�QR3��S���t���Xp�VS!_�`�ד�F��ژ����!?NS�TCY_ E 	L����1�t�1��U���24�2B�NI O�7������DEVIn|� F��$5�wRBTxSPIB�P���BYX����yT��HNDG��G H tn����L��Q�C���5�:�Lo0 H���閻�FBP�{tFE@{�5�t��T��I��DO���uPMCS��v>�f>�t�"HO�TSW�`s��҈E;LE��J T���e �2��25�� O� ��HA7�E��344�0�ܘ�A�K �� MD�L� 2J~PE ��	A��s��tːÈ�s�JÆG!��rD"��0������\�TO��W��	��/��SLAV��L  \0IN�Pڐ���`%ن_C�Fd�M� $n��ENU��OG��`b�ϑ]զP�0`�<��]�IDMA�Sa��\�WR�#��"]�sVE�$a�SKI�S!Ts��sk$��2u���J�������	��Q����_SVh�EXC�LUMqJ2M!ONLD��D�Y��|�PE �ղI_V�APPsLYZP��HID-@�Y�r�_M�2��VRFY�0��r�1�c�IOC_f�� 1�������O��u�LS����R$DUMMKY3�!���S� L_TP/Bv�"����AӞ�ّ N ����RT_u��� ��G&r[�O{ D��P_BA�`g�3x�!F R��_5���H������� �� P $<�KwARGI��� �q�2O N�_wSGNZ�Q �~P/�/PIGNs�l��$�^ sQANNUN�@�T<�U/�ߴ�LAzp]	Z�d~
��DEF�wPI�@ R @��F?IT�	$TOTA%��d����!�M�NI�Y�S+���E�A�[�
DAYS\�A�Dx�@��	� �EFF_AXI?�1TI��0zCOJA� �ADJ_RT+RQ��Up��<P$�1D �r5̀Ll�T�p? ]P�"p��pmtpd��V 0w��G��������S�K�SU� ��CT�RL_CA�� }W�TRANS��6PIDLE_PW����!��A�V��V�_�l�V �D�IAGS���X�w /$2�_SE�#TAC���t!�!0�z*@��RR��vPAh���p ; SW�!@�!�  ��ol�U��foOH��PP� ���IR�r��BRK'#��"A_Ak���x  2x�9ϐZs2��%�l�W�pt*�x%RQ�DW�%MSx�t5A�X�'�"��LIFEgCAL���10��N�1{"�5Z�3{"dp�5�ZU`}�MOTNr°Y$@FLA�c�ZOVC.p�5HE|	��SUPPOQ�ݑ/q� Lj (C�1S_X6�IEYRJZRJWRJ�0TH�!UC��6�XZ_AR�p��YM2�HCOQ��Sf6�AN��w$X��I{CTE�Y `��CACHE�C9øM�PLAN��U7FFIQ@�Ф0�<�1	��6��M�SW�EZ 8�K�EYIM�p��TM~�SwQq�wQ#���}�OCVIE� ��[ A�BGLx��/�}�?� 	��?��D\p�ذST��!�R� �T� �T�� �T	��PEMAI�f�ҁ��_FAKUL�]�Rц�1��U�� �TRE��^< $dRc�uS�% IT�ӇBUFW}�W��N�_� SUB~d��C�|��Sb�q�bSAV �e�bu �B��� �gX��^P�d�u+p�$�_p~`�e�p%yOTT����sP��M��OtT�FLwAX � ��X~`�9#�c_G�3
�YSN_1�_�D��T1 �2M���T�F��H@ g�?`� 0p���Gb-sC_R�AIK ���r�t�RoQ�u�7h�qDSPq��rP��A�IM�c6�\��Ä�s2�U�@�A�sMF*`IP���s�!DҐ�6�TH�@n�)�OT��!6�HSDI3�AGBSC���@ Vyİ�� �_D�CONVI�G���@$3�~`F�!�pd��p�sqSCZ"���sM3ERk��qFB��k��pET���aeRFMU:@DUr`����x�CD,���@p;cH%R�A!��bp�ՔXՔ+PSԕCN�%�C��pN�ғ|Sp�cH *�LX�:cd�Rqa�| �� ��W��U��U��U�P	�U�OQU�7R�8R��9R��0T�^�1k�1�x�1��1��1��1���1��1ƪ2Ԫ2T^�k�2x�2��2��U2��2��2��2ƪ�3Ԫ3^�3k�x�3P���o���3��3���3ƪ4Ԣ�AEXTk!0�d <� 7h�p��6�pO��p����NaF{DRZ$eT^`�V�Gr����䂴2R�EM� Fj��BOV�M��A�TRO�V�DT�`-�MX�<�IN��0,�W!INDKЗ
w�׀�p$DG~q36��P�5�!D�6�RIVx���2�BGEAR�KIO�%K�¾DN�p���J�82�PB@�CZ_MCM�@�1��@9U��1�f ,②aO? ���PI�.�!?I�E��Q�!����`m���g� _05Pfqg RI9ej��k!UP2_ h � �cTD�p����! a��壓�BAC�ri T�P�b�`Z�) OG��%�8��p��IFI�!�p0m�>��	�PT�"���FMR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4�@��Uk��� �T�FS#p�Tl �P���e�qP�p$GEX_���1M�2��2� 3�5��9G ���m ��Ѝ��SW�eOe6DEBcUG���%GR���pU�#BKU_�O�1'� �@PO��I5�5MSf��OOfswSM���E�b֐��0�0_E n �p C _�TERM�o���0�ORI+�p���"�SM_����b�q�!&��TA�r�UP>�Rs� -�1�2�n$�' o$S�EG,*> ELTO���$USE�pNFIAU"4�e1��|�#$p$UFR����0ؐO!�0����OT��'�TAƀU�#N;ST�PAT��P��"PTHJ����Ep�P rF�V"ART�`�`%B`�abU!REL<:�aSHFT��V!\�!�(_SH+@M$�D��� ��@N8r�����OVRq��rSH�I%0��UN� �aAGYLO����qIl�����!�@��@ERV ]��1�?:�¦'�2`��%��5�%�RCq��EASYM�q�EV!#WJi'��}�E���!I�2��U@D��q�%Ba��
5Po��0�p6�OR�MY� `GR��t2b5n� � p��UPa�Uu Ԭ"�)���TOCO!S�1POP ��`�p(C�������Oѥ`KREPR3��aO�P,�b�"ePR�%WU�.X1��e$PWRf��IMIU�2R_	S��$VIS��#(AUqD���Dv" v���$H���P_AD+DR��H�G�"�Q��Q�QБR~pDp1�w H� SZ�a��e`�ex�e��SE�l�r��HS��MNv?x ���%Ŕ��OL���p<Px��-��ACROlP<_!QND_C��גx�1�T �ROUPT���B_�VpQ�A1 Q�v��c_��i���iр�hx��i���i��v�AMCk�IOU��D�g�fsu^d�y $|�P_D��VB`boPRM_�b��A�TTP_אHaz{ (��OBJEr�l�P��$��LE�#��s`{ � \��u�AB_x�T~��S�@�DBGL�V��KRL�YHIoTCOU�BGY �LO a�TEM���e�>�+P'�,PSS�|�P�JQUERY�_FLA�b�HW(��\!a|`u@�3PU�b�PIO��"��]�ӂ/dԁ=dԁ�� _�IOLN��}�����CXa$SL�Z�$INPUTM_g�$IP#�P��L'���SLvpa~���!�\�W�C-�B �y
���pF_ASv��$L ��w �DF1G�U�B0m!���0HY��ڑ���$���UOPs� `������[�ʔ[�і"�[PP�SIP�<�і�I�2��P_MEM�B��i`� X��I1P�P�b{�_N�`����R�����b�SP��p$FOC�USBG;��UJ�Ƃ �  � o7�JOG�'�DISf[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A��oAPHIb�Q�:]�D� J7J\���޷ _KEYt� ��KՀLMONza���$XR���ɀ��WATCH_0��3���EL��}S1y����s� �Ю!qV�g� �CTR3�򲓥��LG�D� ��R��I�
LG_SIZ���J�q I�,��I�FDT�IH�_� jV�GȴI�F�%SO� ��q �Ɩ���v��ƴ��K�S����w�k�)N����E� �\���'�*�U�s5�r�@L>�4�DAUZՃEA�pՀ�Dp�f�G�H�B�OGBO}O��� C����PIT���� ��R{EC��SCRN��ⵖD_p�aMARGf�`��:���T�$L���S�s��W�Ԣ��Iԭ�JGMO�MN3CH�c��FN��R��Kx�PRGv�UF���p0��FWD��H]L��STP��V��+���Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*�a2�8����Gh�0P!O��������M8�Ģv��EX��TUIv�	I��(�4�@� t�x�J0J�~�P���J0��N�a�#ANA8��O"�0VAIA��d�CLEAR�6DCS_HI"�/c�5O�O�SI��9S��IGN_�vp�q�uᛀT�d� DE�V-�LLA �°B�UW`��x0T6<$U�EM��Ł�����"Qa���x0�σ�a�@OS1��2�3���_�`� �ࠜh�ApN%-���-�IDX�D	P�2MRO��Գ!�+ST��Rq�Y{b!� �$E&C +��p.&A&��a� L��ȟ%Pݘ���T\Q�UE�`�US:�c��_ � ��@(��`�����# �MB_PN@ R`r�y�R�w�TRIN��P��BASS�a	6gIRQ6�qMC(��� ��CLD�P�� ETRQLI`��!D�O9=4FLʡh2�Aq3zD�q7���LDq5[4q5ORG �)�2�8P�R��4�/c�4=b-4�t� ��rp[4*�L4q5S�@T�O0Qt�0*D2FRCLMC@D�?�?RIAtr,1ID`�D� d1���RQQprpDS3TB
`� �FᆻHAXD2���G�LE�XCES?R��BMhPa�͠�BD4Y!��B�q`�`�F_�A�J�C[�O�H� K���� \���bTf$�� ��LI�q�SRE�QUIRE�#MOx�\�a�XDEBU���,1L� M䵔 @�p���P�c�AA,1N��
Q�q�/�&���f-cDC��B�IN�a�?�RSM�Gh� Np#B��N�iPST9�� � 4��LO�C�RI���EX��fANG��A,1O�DAQ䵗�@$��9�ZMF�����f���"��%u#ЖVS�UP�%�qFX�@I{GGo�� �rq �"��1��#B��$���p%#by��rx���vbP�DATAK�pE�;����R��M��*�[ t�`MD�qI��A)�v� �t�A�wH�`���tDIAE��sANSW��th���u�D��)�bԣ(@$`�[ PCU_�V6��ʠ�d�PLOr�$`�HR���B���B�p���������MR�R2�E�  ���V�A/A d$OCALI�@��G~��2��!V��<$R�SW0^D"���ABC�hD_J2�SE�Q�@�q_J3:M�
G�1SP�,��@PG�n�3m�u�3p
�@��JkC���2'A�O)IMk@{BCS�KP^:ܔ9�wܔJy�{BQܜ������`_AZ.B��?�E�L��YAOCMP0�c|A)��RT�j�ƚ�1�ﰈ��@1�茨`��Z��SMG0��pԕ� ER!��L� �INҠACk�p����b�n _������h�D�/R��DIU�F�CDH�@
�#a�q�$V�Fc�$x�$���`@���bʺ�� Rc�׀�H �$BELP�|���!ACCEL����kA°IRC_)R�p\�T!�O$PS�@B2LY ���W3�ط9� ٶPATH��.�γ".�3���p�A_���_�e�-B�`C���_{MG�$DD��<ٰ��$FW�@�p`����γ����DE���PPABN�ROTSPEEu��8O0��DEF>Q��~Y $USE_��JJPQPC��JY�����-A 6qYN�@A��L�̐�L�MOUf�NG��|�OL�y�INCU��a�¢��B��ӑ�AENCS����q�B�����D�IN�I�����pzC��VE�����23_�U ��b�LOWL����:�O0��0�D�i�B�PҠ� ��PRC�����MOS� gTM�Opp�@-GPERC�H  M�OVӤ  �����!3�yD!e� ]�6�<�� ʓA����LIʓdWɗ��:p3�.�I�TRKӥ�AY����?Q^���m�b���`p�CQ�� MOM �B?R�0u��D���ay�0Â��DUҐ�Z�S_BCKLSH_C����o�n���TӀ���
c��CLALJ��A��/PNKCHKO0�Su�'RTY� �q��M�1�q_
#c�_UM�CP�	C���SCLܵ��LMTj�_L �0X����E��  �� ���m�hј��6��PC����H�� �P�ŞCN@�"X�T����CN_��N�^C�kCSF����V 6����ϡj���n7CAT�SHs�� ���ָ1���֙�����̭���PA���_P���_P0� e���O1u�$xJG� P{#��OG���TORQU(�p�a�~����R0y������"_W��^􀖡��4t�
5z�
5I*;I ;Iz�F�`�!���_8�1��VC��0�D�B�21�>	P�?�B�5JRK�<�2�6i�?DBL_SM�Q&B�MD`_DLt�&BGRV4
Dt�
Dz��1�H_���31�8JCO1SEKr�EHLN�0hK �5oD��jI��jI<1�J��LZ1�5Zc@y��1M1YqA�HQBTHWMY�THET09�NK�23z�/Rn�r@CB�4VCBn�CqPAS�faYR<4gQt�gQ4VSqBt��R?UGTS���Cq��a��P#���Z�C$DUu ��R@䂥э2�Vӑ��Q�rN�f$NE�+pIs@H�|� �$R�#QA'U�PeYg7EBHBALPHEE.b�.bS�E�c�E �c�E.b�F�c�j�FR�EVrhVghd��lV�jUV�kV�kV�kV�kV�kV�iHrh�f�rP�m!�x�kH�kH�kUH�kH�kH�iOcl�OrhO��nO�jO��kO�kO�kO�kO
�kO�FF.bTQ���E���egSPBALAgNCE��RLE�PH_'USP衅F���F��FPFULC��3��3��E��1��l�UTO_p �%Tg1T2t���2NW �����ǡ��5�`�擳�T�OU���� �INSEG��R�R�EV��R���DIF�H��1���F�1��;�OB��;C��2�� �b�4LCHW3AR��i�ABW!��?$MECH]Q�@Xk�q��AXk�Pp��IgU�i�� 
����!����ROB��C�R��ͥL� ��C��_s"T �� x $WEI3GHh�9�$cc�2� Ih�.�IF ќ�'LAGK�8SK��nK�BIL?�OD��LU��STŰ�P�@; �����������
�Ы�L��  2y�`�"�DEBU.��L&�n��PMMY�9��NA#δ9�3$D&���$��� �Q   �D�O_�A��� <@	���~��L�BX�P�N��+�_7�L�t��OH  �� E%��T���ѼT��<���TICK/�C��T1��%������N��c�Ã�R L�S���S�����PROM�Ph�E� $IR� X�~ ���!҇MAI�0��j���_�9����t�l�Rn�0COD��FU`�+�ID_" =����~�G_SUFF<0G 3�O����DO��ِ��R��Ǔـ��S����!{�������	�H)�_FI���9��ORDX� ����36��X������GR9�S��Z�DTD���v�ŧ�4 *�L_N�A4���K��DEF_I[�K���g��_����i��Ɠ�š���IS`i �萚����e����4�0i��Dg����D� O|��LOCKEA!�uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ�{� ���}��v�Ա�� g������^���K‒Փ����!w�N�P@'���^���,`�W\�l[R��7�TEF�Ĩ �OULOOMB_u�0�wVISPITY��A�!OY�A_FR1Id��(�SI��B�R������3��
�W�W��0��09_,�EAS%��@�!�& "���4p�}G;� h ���7ƵCOEFF_AOm���m�/�G!2%�S.�߲CA5�����u�GR` � � $R� �X]�TME�$R�s�XZ�/,)�ER�T;��:䗰�  ]�LLt��S�_SV�&�($~����@�� "SETU��MEA��Z�x0��u������ � �� �� ȰID@�"���!*��&P���$*�F�'����)3��#���"�5;`:*��REC���!=�MSK_���� P	�1_USER��,��4���D�0��VEL,2�0��ȯ2�5S�I�|��M�TN�CFG}1� � ���Oy�N�ORE��3��2�0S�I���� ��\�UaX-�ܑPDE�A� $KEY_�����$JOG<EנSVIA�WC�� 1DSWy���
��CoMULT�GI�@�@C��2� 4 ��#t�+�z�XYZ���|�����z� �@_7ERR��� ��S L�-���@��s0BB_$BUF-@X1�7ࡐMOR�� H	�CU�A3�z�1Q��
��3���	$��FV��23��A�bG�� � �$SI�@ G�0VOx B`נOBJE&��!FADJU�#EEGLAY' ���SD�W�OU�мE1PY���=0QT i�0�W�DIR$ba�pےʠDYNբHe	T�@��R�^�X����OPWORK}1��,�SYSB9U@p 1SOP�aR$�!�jU�k�PR��2�ePA�0�!�cu� 1+OP��UJ��a'�zD�QIMAG�A1	��`i�IMACr�IN,�bsRGO�VRD=a�b�0�aP �`sʠ� �^uz��LP�B�@��!PMGC_E,�Q��N@�M�rǱ��1Ų7�=q�SL&�~0���$OVSL\G*E��"*E2y�Ȑ�_=p�w ��>p�s���s	�����y�z=q�#}1� @h�@;���OE�RI#A��
N��X�s�f�ՠ����PL}1�,RT�v�m�ATUSRBT�RC_T(qR��B  �����$ �Ʊ��,�~0� D��`-CSALl`�SA���]1gqXE���%���C�1�J�
���UP(4�����PX��؆�q��3��w� �PG�5�� $SUBࠁ����t�JMP�WAITO��s��L�OyCFt�!D=�CV!F	ь�y���R`�0~��CC_CTR�Q��	�IGNR_P�Lt�DBTBm�P���z�BW)����0UL@���IG�a��Iy�OTNLN��Z�R]a�K� N��`B�0�PE��s���r��f�SPD.}1� L	�A�`g����S��UN�{���r]�R!�`BDLY��2���7�PH_�PK�E��2RETRIEt��2�b6��v��FI�B� ��м�8� 2��0D�BGLV�LOGgSIZ$C�KTؑ�Uy#u�D7�_�_T,1@�EM�@C\1aAě���R��D�FCHgECKK�R�P�0ʳ���@&�(bLE,c�" PA9�T���PJ�C߰PN�����ARh�0���Ӯ�P�O�BORMATTnaF�f1h���2�LS��UXy`	����LB��4�  rEITCH�B7�9�PL)�AL_ G� $��XPB�q�� C,2D�!��+2�wJ3D��� T�pPDCKyp��oC� �_ALPH���BaEWQo���� ��|I�wp � �b@?PAYLOA��m��_1t�2t���J3AR��؀դ֏�la�TIA4��5��6,2MOMCP������h�����0BϐAD��p������PUBk`R��;���;�������z4�` I$PI\Ds�oӓ1yՕ�w�T2�w�Z��I��I��I���p����n���y�e`�9S)bT�S/PEED� G��(� Е��/���Е�`/��e�>��M��ЕSAMP�6V��/���Е#MO�@ 2@�A�� QP���C��n������� ����LRf`kb�ІE9h�EIN09��7 S.В9
yPy�/GAMM%S���D$GET)bP�ciD]��2
�IB�:q�I�G$HI(0;�A��LREXPA8)LWVM�8z)��g���C�5�CHKKp]�0�I_��h`eT��n� q��eT,����� �$�� �1�iPI� RCH�_D�313\��30L�E�1�1\�o(Y�7 ¾t�MSWFL �M.��SCRc�7�@�&���%n�f�SV���PB``�'�!�B�sS_SAV&0ct5B3NO]�C\�C2^� 0�mߗ�uٍa��u� ��u:e;��1���8��D�P��������� )��b9��e�GEX�3��V�4�f�Ml��� � �YL(��QNQSRlb fqXG�P�RR#dCQ�p� �S:AW70�B �B[�CgR:AMxP�K�CL�H���W�r�(1�n�g�M�!o�� �8F�P@}t$WP�u �P r��P5�R<�R C�R��%�6�`��� (��qsr X��OD�q�Z�Ug�ڐ>D� ��OM#w�J?\? n?�?�?��9�b"���tg�]�_��� |� �X0��bf��qf��q`��ڏgzf��Eڐ� S�Ag�"ɵ��кFdPB��PM�Q}U�� � 8L��QCOU!h QT�HI�HOQBpHY�SY�ES��qUE��`�"�O���  b�P�@\�UN��ʄCf�O�� �P��Vu��!����O�GRAƁcB2�O��tVuITe �q:pINFO�����{�q�cB�e�OI�r� =(�@SLEQS��q���p�vgqS����� 4L�ENAB|DRZ�PTIONt������Q���)�GCF:��G�$J�q^r�� R���U�|g�d�OS_ED��N��� �F��PK��j��E'NU߇�وAUT$1܅CO�PY�����n�00M�N���PRU�T8R �Nx�OUN��$G[rf�e�_RGADJ���*�3X_:@բ$�����P��W��P��} ���)�}�EX�YCZDR|�NS.��F@�r�LGO�#�NY�Q_FREQR�W`� �#�h�TsLAe#�����ӄ �CRE�� s�IF��sNmA��%a�_Ge#STATUI`e#MAIL�����q �t�������ELE�M�� �/0<�FEASI?�B��n��ڢ�vA�]� � I �p��Y!q]�t#A��ABM���E�p<�VΡY�BASR�Z���S�UZ��0$�q���RMS_TR ;�qb ���SY�	�ǡ���$���>C�Q`	~� 2� _ �TM������̲�@ ��A��)ǅ�i$DOUd�s]$Nj���PR+@z3���rGRID�q�M�BARS �TY�@��OTO�p��� Hp_}�!����d��O�P/�� � �p�`POR�s��}�.��SRV��)����DI&0T����� �#�	�#�4!�5!�6J!�7!�8�6AF��2��Ep$VAL�Ut��%��ֱ��/��� ;�.1�q��1���(_�AN�#��ⓡRɀ(���TOTcAL��S��PW��Il��REGEN�1�cX��ks(��a����`TR��R��_!S� ��1ଃV�����⹂Z�E��p�q���Vr���V_H��DqA�S����S_Y,1��R4�S� AR�P2�� ^�IG_S!E	s����å_Zp���C_�Ƃ�ENHA�NC�a� T �;�������IN�T�.��@FPsİ_OVRH�P�`p�`��Lv��o��7�}���Z�@�SLG�AA�~�25�	��D��YS�BĤDE�U�̦���TE�P���G� !Y��
�J��<$2�IL_MC�x r#_��`TQ�`��q����'�BV�C�P�_� 0�M�	V1V�
V1�2�2�U3�3�4�4�
 �!���� � m�A�2;IN~VIBP����1�2�2�3*�3�4�4�A@p-�C2���p� �MC_Fp+0B�0L	11d���M501Id�%"E� S`�R�/�@KEEP__HNADD!!`$$^�j)C�Q���$��"	��#O�a_$A�!pK��#i��#REM�"��$��½%�!�(U�}�e�$HPWD � `#SBMSUK|)G�qU2:��P	�COLLAB � �!K5�B�� ��g��pITI1{9p#n>D� ,�@FLAP>��$SYN �<�M�`C6���UP�_DLYAA�ErDGELA�0ᐢY�`�AD�Q��QSwKIP=E� ���XpOfPNTv�A�0P_Xp�rG�p�RU@ ,G��:I+�:IB1:IG� 9JT�9Ja�9Jn�9J{к9J9<��RA=s� X���4�%1�Q}B� NFLIC�s��@J�U�H�LwNO�_H�0�"?��RIT�g��@_PA�pG��Q� �K�^�U�W��LV�d�NGRLT�0_q��O�  p" ��OS��T_JvA� V	�APPR_W�EIGH�sJ4CH?pvTOR��vT���LOO��]�+�tVJ�е�ғA�Q�U�S�X�OB'�'�2��J2TP���7�X�T� <a43DP=`Ԡ\"<a�q�\!��RDC��L�+ �рR��R�`� ��RV��jr�b�R�GE��*��cN�FL�G�a�Z���SPC��s�UM_<`^2�TH2NH��P.a �1� m`EFv11��� lQ `�!#� <�p3AT�  g�S��Vr�p�tMq�Lr���HOME(wr�t2'r�-?�Qcu��w3'r逪������w4'r�'�9�K�]�o���
�w5'r뤏��ȏڏ(����w6'r�!�3��E�W�i�{��w7'r퀞���ԟ����w8'r��-�?�Q�c�u�R�uS$0�q�p�� sF��`la�!`P�����`/���-�IO[M�I֠��q�POWE�� ���0Za*��� ��5��$DSB� GNAL���0C�p��OF�RS2;323�� �~`��9� / ICEQP��cPEp��5PIT�����OPBx0��FLOW�@TRvP��!�U���CU�M��U�XT�A��w�ERF�AC�� U���p�SCH��� t�Q  _��>�Q$L����OM��A�`�T�P#UPD7 Ad�ct�T��UEX@8�ȟ�U EFA: X"΁1RSPT����)�T ��PPA�0o�l���`EXP�IOS���)ԭ�_���%Ќ�C�WR�A��ѩD�ag֕`ԦFRIE3NDsaC2UF7P��ޤ�TOOL��MY�H C2LENGT_H_VTE��I�<�Ӆ$SE����?UFINV_����RGI�{QITI5B��Xv��-�G2-�G17�w�S�G�X��_��UQQD�=#���AS��d~C��`��q�� �$$�C/�S�`������S0)�����VERsSI� ��)��5��I��������AAVM_Y�2� � �0  �5���C�O�@�r� r�	 ����S0�!����������������
?QY�B�S���1��� <-�� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O�OiCC�@XLM�T��C�  ��DIN�O�A�Dq�EXE�HPV_���ATQz
��L�ARMRECOV� �RgLM_DG *�5���OLM_IF 	*��`d�O�_�_�_ �_j�_'o9oKo]onm, 
��odb���o�o�o�o^��$� yz, A   2�D{�PPINFO7 u[ �Vw��������`� ������*��&��`�J���n�����DQ� ���
��.�@�R��d�v���������a
P�PLICAT��?��P��`�Handlin�gTool 
� �
V8.30P�/40Cpɔ_LI
883��ɕ$ME
F0G��4�-

39�8�ɘ�%�z�
?7DC3�ɜ^
�NoneɘVr����ɞ@6�d� Vq_ACT#IVU��C죴�MODP���C�I��?HGAPON����OUP�1*�� i�m�����Қ_����1*� ) �@������� ��Q���Կ�@�
������ ���5�Hʵl�K�HTTHKY_� �/�M�SϹ������� ��%�7ߑ�[�m�� �ߣߵ���������� !�3��W�i�{��� ������������/� ��S�e�w��������� ������+�O as������ �'�K]o �������� /#/}/G/Y/k/�/�/ �/�/�/�/�/�/?? y?C?U?g?�?�?�?�? �?�?�?�?	OOuO?O QOcO�O�O�O�O�O�O �O�O__q_;_M___ }_�_�_�_�_�_�_k�ƭ�TOp��
�DO?_CLEAN9�ꤾpcNM  !{ 衮o�o�o�o�o��DSPDRYRwo&��HI��m@�or ����������&�8�J���MAX@ݐWdak�H�h�XWd��d���PLUG�GW�Xgd��PRC*)pB�`�kaS��Oǂ2DtSEGF0�K� �+��o�o�r����������%�LAPOb�x�� �2� D�V�h�z�������¯�ԯ�+�TOTAL�����+�USENU
O�\� e�A�k­��RGDISPMM�C.���C6�z�@I@Dr\�OMpo�:��X�_STRING� 1	(�
�kM!�S�
���_ITEM1Ƕ  n������+� =�O�a�sυϗϩϻπ��������'�9��I/O SIG�NAL��Tr�yout Mod�eȵInpy�S�imulated�̱Out���OVERRLp =� 100˲In� cycl�̱�Prog Abo�r��̱u�Sta�tusʳ	Hea�rtbeatƷMH Faul	��Aler�L�:� L�^�p��������� ScûSaտ ��-�?�Q�c�u����� ����������)�;M_q��WOR .�û������ +=Oas� ������//'.PO����M � 6/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l?�~?�?�?�?�?H"DEVP.�0d/�?O*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_>n_PALT	��Q �o_�_�_�_�_oo )o;oMo_oqo�o�o�o��o�o�o�o�_GRIm�û9q�_as �������� �'�9�K�]�o�������'�R	�݁Q�� ��)�;�M�_�q��� ������˟ݟ����%�7�I�ˏPREG �^����[�����ͯ߯ ���'�9�K�]�o� ��������ɿۿ�Oݿ�$ARG_� D ?	���0���  �	$O�	[�D�]D��O�e�#�S�BN_CONFIOG 
0˃����}�CII_SA_VE  O������#�TCELLSETUP 0��%  OME_I�OO�O�%MOV�_H������REP���J��UTOBA�CK�����FRA:\o�c Q�o���'`��qo��ҟ�� �� f�o������*�!�3�`�Ԉ�� f����������o� {��&�8�J�\�n��� ���������������� "4FXj|�������끁�  ��SYSUI�F.SV V T�.TP D MP� 6.VD GIF 7N`r�o��N.E#��f�INUI�Po���c�?MESSAG������8��ODE_D����z��O�0�c�oPAUSM!!�0�? (73�U/g+(Od/�/x/�/ �/�/�/�/�/???�P?>?t?1�0$: TSK  @-��T�f��UPDT��d��0
&XWZD_E�NB����6STAp�0��5"�XIS��?UNT 20Ž�� � 	 �I�20�e���� ��?�z⶙�E� �2�џ��HsM�Oo��}C��� �D�O�O�O _�?5C�MET߀2CMP�TA@4;?����?�/�@5���@��@��]4��4���%4cG.5q��24h�@4����8]SCRDC�FG 1�6��Ь�H  _�_oo(o:oLo��o�Q���_�o�o�o�o �o�o]o�o>Pb�t���o9�i�G�R<@M/�sUP_kNA�/�	i�n�v_ED�1�Y�� 
 �%-BCKEDT-��'�GETDATAU�o�9��?�j�H�o�f�\��A�^�  ���2�0&�!�E���:IB����~�ŏ׏m����3 ��&۔��D��ߟJ� ����9�ǟ�4��� ϯ�(����]�o�����5N������(��w��)�;�ѿ_��6 ϊ�gϮ�(�CϮ���ϝ�+��7��V�3� z�(��z�����i���B�8��&���~�]����F�ߟ�5����9~������]����`Y�k�����CR� !ߖ���W�q���#�5����Y��p$�NO_D�EL��rGE_U�NUSE��tIG�ALLOW 1z��(**�TEM*S	$SERV_GR��V� : REG�q$�\� NUM�
<��PMUB U�LAYNP\PMPAL�>CYC10#6� $\ULSU`�8:!�Lr~�BOXORI��CUR_��PoMCNV��10L�T4DL!I�0��	����B N/`/r/�/�/�/�/�/����pLAL_OU�T �;���qW?D_ABOR=f��q;0ITR_RT�N�7�o	;0NON�S�0�6 
HCC�FS_UTIL s#<�5CC_@�6A 2#; h� ?�?�?O#O6]CE�_OPTIOc8�qF@RIA_IIc f5Y@�2�0�F�Q�=2q&}ނA_LIM�2�.� �K �]B���KXK 
K �,2O�Q��B�r�qFK Q5T1)TR�H�_:JF_PA�RAMGP 1�<g^&S�_�_�_��_�VC�  C��d�`�o!o`��`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?���2HE ONFI�� E?�aG_P�1#; ���o 1CUgy�a�KPAUS�1�yC ,���� �����	�C�-� g�Q�w���������я4���rO�A�O�H~�LLECT_�B1�IPV6�EN. QF܍3�NDE>� ��G�71234567890���sB�TR����%
 	H�/%)����� ��W���0�B���f�x� ��㯮���ү+���� �s�>�P�b������� ���ο��K��(Ϡ:ϓ�^�|��B!F�� �I|�IO #��<U%e6�'��9�K���TR�P2$���(9X�t�Y޼`�%�̓ڥH��_MO�R�3&�=�K XB2�a��A� $��H�6�l�~���~S"��'�=�r_A?�a�a�`��K K��R�dP�)F�ha�- �_�'�9�%
�k���G� ��%Z�%���`K c.�PD�B��+���cpmidbg��	3 F:��D����p��|N  �K ğ1���]�`��{<�^�K čzg�$� o�sfl�q��ud1:��:J��?DEF *ۈ���)�c�buf.txt�����_L64FIX ,������l/[Y/ �/}/�/�/�/�/
?�/ .?@??d?v?U?�?�?��?�?�?�?,/>#_E -���<2ODO`VOhOzO�O6&IM���.o�YU>����d�
�IMC��2/�����dU�C��20��M�QT:Uw�Cz � B�i�A����A�jA@���B3�*CG��B<�=w�i�B.���B�v1B����B�$�D��%B���ezVC�it&C��C��n�D-lE?\D�n�jlJ��22o�D|���0�0 �0�'��C����
�x�Obi�D4cdv`D��`/�`v`s]E�D� D�` E4��F*� Ec���FC��u[F����E��fE���fFކ3FY_�F�P3�Z��@��33 ;��>�L���Aw�n,a@:�0@e�5Y���a����`A��w�=�`<#���
��?�ozJ�RSMOFST c(�,bIT1��eD @3��
д���,�a��;��bw�?���<�M^�NTEST�1O��CR@�4��>VCF5`A�w�Ia+a�a�ORI`CTPB�U�C��`4���r�0:Sd����qI?�5���qT_�PRO'G ��
�%$/ˏ��t��NUSER � �U������KE�Y_TBL  �����#a��	
��� !"#$%�&'()*+,-�./��:;<=>�?@ABC�GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~��������������������������������������������������������������������������������͓���������������������������������耇��������������������������LCK��
����STAT�/��s_AUTO_�DO �	�c�INDT_ENBP�b��Rpqn�`�T2�����STOr`���X�C�� 26���8�
SONY XOC-56�"b�����@��F( ����HR50�w���>�P�7b�t�A�ff����ֿ�  Ŀ����C�U�0�y� ��fϯ��Ϝ������ϸ�-ߜ�TRL��L�ETEͦ ��T�_SCREEN ���kcs����U�MMEN�U 17�� <ܹ���w������ ����K�"�4��X� j������������ 5���k�B�T�z��� ������������ .g>P�t�� ����Q( :�^p���� /��;//$/J/�/ Z/l/�/�/�/�/�/�/ �/7?? ?m?D?V?�? z?�?�?�?�?�?!O�? 
OWO.O@OfO�OvO�O��O(y��REG 18�y����`�M�����_MANUAL��k�DBCO��R�IGY�9�DBG_oERRL��9��q��_�_�_ >^QNUMLI�pϡ���d
�
^QPXWORK 1:���_5oGoYoko}oӍ�DBTB_N� �;������ADB_AWAYzfS�qGCP 
�9=�p�f_AL�pR���bbRY�[�
�WX_��P 1<{y�n�,��%oc�P��h_MM��ISO��k@L���sONTIMX�M�
���vy
���2sMOTNEND��1tRECORDw 1B�� ���sG�O�]�K��{ �b��������V�Ǐ� ]����6�H�Z��� ������#�؟���� ��2���V�şz����� ���ԯC���g��.� @�R���v�寚�	��� п���c�χ�#ϫ� `�rτϖ�Ϻ�)ϳ� M���&�8ߧ�\�G� Uߒ�߶�����I������4�� �p7�n� ���ߤ�������� �"���F�1���|��� ������[�����i����BTf���bTOLERENC�dsB�'r�`L��^P�CSS_CCSCOB 3C>y�`IP�t}�~�< �_`r�K�����/�{��5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O_�~ֽLL� D���&qET�c�a C[C�`ZP^r_W A� p� �s�p��QGPt[	 !A�p�Q�_�[? �_h�[oU�p��p�pSB�V�c�(a@�PWoio{h+�o�Xa�o�oY��[�	r�hN�>������AAs�<�h8<K��c���aD@VB���|�G����+��K� A�otGhXGr�S�o����eB  _ =��Ͷa>�t&YB�� �pC�p�q
�aA"�H�S�Q-��q ���ud�v�����Af�P ` 0����D^P��p@�a
�QXTHQ����a� aW>� �a9P� �b�e:�L�^�h�Hc�́PQ�RFQ�PU�z �֟�o\^��-�?���c�u����zCz�ů�b2�Щ�RoD�������Z� ����S̡0��]�0� .��@���EQ�p�� F�X�ѿUҁп�VS�ȺNSTCY S1E��]�ڿ ��K�]�oρϓϥϷ� ���������#�5�G��Y�k�}ߏߒ��DEVICE 1F5� MZ�۶a��	�@ ��?�6�c���	{�𰟗��_HNDGD G5�VP���R>�LS 2H�ݠ� �/�A�S�e�w������ ZPARAM �I�FgHe�RBoT 2K��8р�<��WPpC�C�,`¢P��|}���%{�C*  � 2�jMTLU,`"nPB, s��M� `}�gT�g��
B��!�bcy�[2D chz����/���/gT#I%D��C�` b!�R���A��A,�ͿBd��A��P���_C4kP�!2�C���$Ɓ�]�ffA��À��B�� ��| ���/�/�T ( �P54a5�}%/7/ d?/M?_?q?�?�?�? �?�?O�?OO%O7O IO�OmOO�O�O�O�O �O�O�OJ_!_3_�_�_ 3�_�_�_�_�_o�_ (ooLo^oЁ=?k_Io S_�o�o�o�o�o�o �o#5G�k} �������H� �1�~�U�g�y�ƏAo �Տ���2�D�/�h� S���go����ԟ���� ϟ���R�)�;��� _�q����������ݯ �<��%�7�I�[�m� ��������}�&�� J�5�n�YϒϤϏ��� ��ѿ������F�� /�Aߎ�e�w��ߛ߭� ��������B��+�x� O�a��������� ��,���%�b�M���q� ������������� �L#5�Yk} ��� ��6 1CUg��� �����	//h/ ���/w/�/�/�/�/�/ 
?�/.?@?I/[/1/ _?q?�?�?�?�?�?�? �?OO%OrOIO[O�O O�O�O�O�O�O&_�O _\_3_E_W_�_?�_ �_�_�_�_"ooFo1o joE?s_�_�om_�o�o �o�o�o0f= Oa������ ����b�9�K��� o���Ώ��[o��(� �L�7�I���m�������$DCSS_S�LAVE L����ё���_4D  �љ��CFG MMѕ��������FRA:\�ĐL-�%04d.wCSV��  }��� ���A i�CH
q�z������|�����"������Ρޯx̩�Ґ-��*�����_CRC_OU/T N�������_FSI ?>њ ���� k�}�������ſ׿ � ����H�C�U�gϐ� �ϝϯ��������� � �-�?�h�c�u߇߰� �߽���������@� ;�M�_������� ��������%�7�`� [�m������������ ����83EW� {������ /XSew� ������/0/ +/=/O/x/s/�/�/�/ �/�/�/???'?P? K?]?o?�?�?�?�?�? �?�?�?(O#O5OGOpO kO}O�O�O�O�O�O _ �O__H_C_U_g_�_ �_�_�_�_�_�_�_ o o-o?ohocouo�o�o �o�o�o�o�o@ ;M_����� �����%�7�`� [�m��������Ǐ�� ����8�3�E�W��� {�����ȟß՟�� ��/�X�S�e�w��� �����������0� +�=�O�x�s������� ��Ϳ߿���'�P� K�]�oϘϓϥϷ��� ������(�#�5�G�p� k�}ߏ߸߳����� � ����H�C�U�g�� ������������ � �-�?�h�c�u����� ����������@ ;M_����� ���%7` [m����� ��/8/3/E/W/�/ {/�/�/�/�/�/�/? ??/?X?S?e?w?�? �?�?�?�?�?�?O0O +O=OOOxOsO�O�O�O��O�C�$DCS_�C_FSO ?�����A? P �O�O _?_:_L_^_�_�_�_ �_�_�_�_�_oo$o 6o_oZolo~o�o�o�o �o�o�o�o72D Vz����� ��
��.�W�R�d� v������������ �/�*�<�N�w�r��� ������̟ޟ��� &�O�J�\�n������� ��߯گ���'�"�4� F�o�j�|�������Ŀ ֿ������G�B�TϾ�OC_RPI�N _jϳ����ς��O��`��1�Z�U��NSL��@&�h߱��������� "��/�A�j�e�w�� ������������ B�=�O�a��������� ��������'9 b]o����� ���:5GY �}������ ///1/Z/U/g/y/ �/�/�/�/�/�/�/	? 2?-???Q?z?u?��� �߆?�?�?�?OO@O ;OMO_O�O�O�O�O�O �O�O�O__%_7_`_ [_m__�_�_�_�_�_ �_�_o8o3oEoWo�o {o�o�o�o�o�o�o /XSew� �������0� +�=�O�x�s������� ��͏ߏ���'�P��K�]�o����� �PR�E_CHK P�۪�A ��,�8�2��� �	 8�9�K��� +�q���a�������ݯ �ͯ�%��I�[�9� ���o���ǿ��׿�� �)�3�E��i�{�Y� �ϱϏ��������� ��-�S�1�c߉�g�y� ���߯����!�+�=� ��a�s�Q����� ���������K�]� ;�����q��������� ����#5�Ak {����� �CU3y�i ������/-/ G/c/u/S/�/�/�/ �/�/�/??�/;?M? +?q?�?a?�?�?�?�? �?�?�?%O?/Q/[OmO O�O�O�O�O�O�O�O _�O3_E_#_U_{_Y_ �_�_�_�_�_�_�_o /ooSoeoGO�o�o=o �o�o�o�o�o= -s�c��� ����'��K�]� woi���5���ɏ���� ����5�G�%�k�}� [�������ן�ǟ� ���C�U�o�A����� {���ӯ����	��-� ?��c�u�S������� Ͽ῿�����'�M� +�=σϕ�w�����m� �����%�7��[�m� K�}ߣ߁߳��߷��� �!���E�W�5�{�� �ϱ���e�������	� /��?�e�C�U����� ����������= O-s����] ����'9] oM������ �/�5/G/%/k/}/ [/�/�/��/�/�/�/ ?1??U?g?E?�?�? {?�?�?�?�?	O�?O ?OOOOuOSOeO�O�O �/�O�O�O_)__M_ __=_�_�_s_�_�_�_ �_o�_�_7oIo'omo o]o�o�o�O�o�o�o !�o1W5g� k}������ /�A��e�w�U����� ��я��o����	� O�a�?�����u���͟ �����'�9��]� o�M���������ۯ�� ǯ�#�ůG�Y�7�}� ��m���ſ�����ٿ �1��A�g�E�wϝ� {ύ�������	�߽� ?�Q�/�u߇�e߽߫� ���������)��� _�q�O�������� ������7�I���Y� �]������������� ��!3WiG� �}����%� A�1w�g� �����/+/	/ O/a/?/�/�/u/�/�/ �/�/?�/9?K?�/ o?�?_?�?�?�?�?�? �?O#OOGOYO7OiO �OmO�O�O�O�O�O_ �O1_C_%?g_y__�_ �_�_�_�_�_�_o�_ +oQo/oAo�o�owo�o �o�o�o�o);U_ _q����� ���%��I�[�9� ���o���Ǐ����� ۏ!�3�M?�i��Y� ������՟�ş�� ��A�S�1�w���g��� �������ӯ�+�=���$DCS_SG�N QK�c���7m� 12�-FEB-19 �10:06   |O�l�4-JANt��08:38}������ N.D������������h�x�,rWf*σ��^M��  O�VE�RSION �[�V3.5.�13�EFLOG�IC 1RK���  	����P�?�P�N�!�P�ROG_ENB � ��6Ù�o�U?LSE  TŇ��!�_ACCLI�M����Ö���WRSTJNT��c��K�EMO�x̘��� ���INIT S.�G�Z����OPT_SL ?�	,��
 	�R575��Y�74j^�6_�7_�50��1��2_�@ȭ��<�TO  Hݷ���V�DEX��d�c����PATHw A[�A\��g�y��HCP_CLNTID ?��6� @ȸ�����IAG_GRP� 2XK� ,`����� �9�$�]�H������1234567�890����S�� |�������!�� ��H���;�dC�S���6�� ���.�R v�f��H�� //�</N/�"/p/ �/t/�/�/V/h/�/? &??J?\?�/l?B?�? �?�?�?�?v?O�?4O FO$OjO|OOE��O y��O�O_�O2_��_�T_y_d_�_,
�B^ 4�_�_~_`Oo�O &oLo^oI��Tjo�o.o �o�o�o�o �O'�_ K6H�l��� ����#��G�2� k�V���B]���Ǐُ �������(��L�B\�B_�
Ĥ��GC*��@�b�.f� >���:�����ߟʟܟ����CT_CON�FIG Y��|Ӛ�egU����STBF_TTS��
��b����Û�:u�O�MAU��|�~�MSW_CF6��Z��6��OCVI�EW��[ɭ������-�?�Q�c�u� G�	�����¿Կ��� ���.�@�R�d�v�� �ϬϾ�������ߕ� *�<�N�`�r߄�ߨ� ����������&�8� J�\�n���!���� ���������4�F�X��j�|����RC£\�e��!*�B^�������C2g{�SB�L_FAULT �]��ި�GPM�SKk��*�TDI�AG ^:�ա�I��UD1:� 6789012�345�G�BSP �-?Qcu�� �����//)/�;/M/� �
@�q��/$�TREC	P��

��/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO�0OBOi/{/xO�/UM�P_OPTIONk���ATR¢l��	��EPMEj��OY�_TEMP  ?È�3B�J�Ps�AP�DUNI���m�Q��YN_BR�K _ɩ�EMGDI_STA"U��aQK�XPNC_S1`ɫ �FO�_�_
�^
�^dpOoo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{�E���� �y�Q��� �2�D� V�h�z�������ԏ ���
��.�@�R�d� �z�������˟�� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i������� ��ÿݟ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�{�iߗߩ߻�տ�� ����'�9�K�]�o� ������������� �#�5�G�Y�s߅ߏ� ����i������� 1CUgy��� ����	-? Qk�}������� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?u? �?�?�?��?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_m?w_�_�_�_�? �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9Ke_W ����_�_��� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�]oy������� �ӟ���	��-�?� Q�c�u���������ϯ ����)�;���g� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�_�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�W� E�s������ߧ����� ��'9K]o �������� #5O�a�k}� E������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-?G Yc?u?�?�?��?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_Q?[_m__ �_�?�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ I_Sew��_�� �����+�=�O� a�s���������͏ߏ ���'�A3�]�o� ������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 9�K�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� �����ߑ�C�M�_� q߃ߝ��߹������� ��%�7�I�[�m�� ������������� !�;�E�W�i�{��ߟ� ����������/ ASew���� ���3�!O as������� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?+=G?Y?k?!?� �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	_#?5??_ Q_c_u_�?�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o -_7I[m�_ �������� !�3�E�W�i�{����� ��ÏՏ����%/� A�S�e�q������� џ�����+�=�O� a�s���������ͯ߯ ����9�K�]�w� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������'� 1�C�U�g߁��ߝ߯� ��������	��-�?� Q�c�u������� ����m��)�;�M�_� y߃������������� %7I[m �������� !3EWq�{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/�/+?=?O? i_?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O?� �$ENETM�ODE 1aj5��  
0054_F[P�RROR_PRO/G %#Z%6�_��YdUTABLE  #[t?�_�_�_�gdRSEV_NU�M 2R  ��-Q)`dQ_AU�TO_ENB  qPU+SaT_NO>a� b#[EQ(b�  *��`��`��`��`4`+�`�o�o�oZdHIS%c1+P�Sk_ALM 1c.#[ �4�l0+�o;M_q���o_b``  �#[aFR�zPTC�P_VER !�#Z!�_�$EXTLOG_REQ�fs�Qi,�SIZ5��'�STKR�oe��)�TOL  �1Dz�b�A '�_BWD�p��Hfܻ�D�_DI�� dj5SdDT1KRņSTEPя�P>��OP_DOt�Q�FACTORY_�TUN�gd<�DR_GRP 1e#YNad 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ� ԟ���1��U�@�y� d�v�����ӯ����LW
 J%�,�,��tۯ�j�U���~y�B�  B୰}���$  A@��s�@UUUӾ����|���E�� E�`�F@ F�5U�/�,��L���M���Jk�L�zp�JP��F�g�f�?�  �s��9�Y9}��9��8j�
�6��6��;��	�\��鉵 �� �
H 	ȥ��ma͜[FEAT?URE fj5���JQHan�dlingToo�l � "
P�Englis�h Dictio�nary�def�.4D St��ard�  
�! hAnalog I/OI׿  !
IX�g�le Shift�I�d�X�uto �Software� Update � rt sѓ�ma�tic Back�up�3\st���ground� Edit��f�d
CamWera`�Fd�e���CnrRndIm����3�Comm�on calib� UI�� Eth�e�n��"�Mon�itor�LOA�D8�tr�Relgiaby�O�ENS��Data Acq�uis>��m.f�dp�iagnos���]�i�Docum�ent ViewyeJ��870p��ual Chec�k Safety�*� cy� �han�ced Us��F�r����C �xt�. DIO :�f�i�� m8���en]d��ErrI�L���S������s  t� Pa�r[�� ����J944�FCTN Men�u��ve�M� J9�l�TP InT�f�ac{�  744���G��p Mas_k Exc��g�� R85�T��Proxy Sv��  15 J�i�gh-Spe��S�ki
� R738�Г��mmuni�c��ons�S R7��urr�T�d��022��aю�connect 2�� J5��Incr���stru,Қ�2� RKARE�L Cmd. L���ua��R860~hRun-Ti��EnvL�oa��K^U�el +��s���S/Wѹ�7�Li�cense���r�odu� ogBo�ok(Syste�m)�AD p�MACROs,>��/Offs��2�NDs�MH��9 ����MMRC�?�ޙ�ORDE� ec_hStop��t? n� 84fMi$�,|� 13dx��]�p��׏���Modz�_witchI�VP��?��. sv<��2Optm�8�2��fil��I ��z2g 4 !+?ulti-T������;�PCM gfunY�Po|����4$�b&Regir� r �Pri���FK+7���g Nu�m SelW  �F�#�� Adj9u���60.��%�|� fe���&tatu�!$6���%���  9 J6�RDM Robo}t)�scove2�� 561��Rem�U�n@� 8 (|S�F3Servo���ҩ�)SN�PX b�I�\d�cs�0}�Libr<1��H� �5б f�0��58��S�o� tr�ssag�4%G 91�p Ȓ�&0���p/Iތ�  (ig TM�ILIB(MӋ�Fgirm����gd7����s�Acc�����0�XATX�Hel	n��*LR"1���Spac�Arqu>z�imulaH��ѹ Q���Tou�Pa��I��T��c���&��ev. f.�svUSB �po��"�iP�a��  r"1Unexcept��`0i$�/����H59� VEC&�r��[6����P{��RcJPRIN<�V�; d T@�TSP CSUI՚� r�[XC��#W�eb Pl6�%d# -c�1R�@4dp�����I�R66?0�FV�L�!FVGrid~K1play C�`lh@����5RiR�R�.@���R-35i�A���Asci�i���"��� 51�f�cUpl� � �(T����S��@r�ityAvoid�M �`��CE��r9k�Col%�@�GuF� 5P��j}P�����
 B�L�t� W120C C� o���!J��P��y��� �o=q�b @DCS- b ./��c��O��q��`�; ���q�ckpaboE4�D�H@�OTШ�mai'n N��1.�H��Gan.��A> aB!GFRLM���!i ��~�MI Dev� s (�1� h8j��spiJP��� �@��D�Ae1/�r���!hP� M-2� i��߂^0i�p6�P}C��  iA/'�?Passwo�qT�ROS 4����q�eda�SN��ClAi����G6x Ar��� 47�!���5s��DER��Tsu�p>Rt�I�7 (9M�a�T2DV�
�3D Tri-���&��_8;�
�A�@Def?����{Ba: deRe p 4t0��e�+��V�st64MB �DRAM�h86�΢FRO֫0�A;rc� visI���n��7| ), <�b�Heal�wJ�{\h��Cell`�2�p� �sh[���� Kqw�c� - ��v���p	VCv�t�yy�s�"Ѐ6�ut��v�m��"�xs ���TD_0��XJ�m�` 2��a[��>R tsi�MA3ILYk�/F2�h�|�ࠛ 90 H��(F02]�q�P5'����T1C��5��@FC��U�F9�Gig�EH�S�t�0/A� cif�!2��boF��dri=c ��OLF�S����" {H5k�OPT �򆧊49f8���cCro6��@��l�A�pA�Syn.(RSS) 1L�\1y�rH�L� (2x5�5��d�pCVx9����e�st�$SР��> \�pϐSSF�e$�tex�D o���A��	� BP���a�(R;00�Qirt��:���2)�D��1�e�V}Kb@l Bui, 9n��WAPLf�į0��Va�kT�XCG�M��D��L����[CcRG&a�YBU��YKfL��pf��k�7\sm�ZTAf�@�О�Bf2�и��V�#�s���� r���CB���
f���W�E��!��
���T�p��DT�&4 1Y�V�`��EH�����
�61Z��
�R�=2�
�E (Np��F��V�PK�B���#��GHf1`?G���H��р?I�e ����L�D�L��N��7\@s@���`���M��Odela<,��2�]M�� "L[P� �`?��_�%�����5S��-F�TSO��W�J57��VG�F�|�VP2֥ 5\b�`0&�cV:����T;T� �<�c�e,?VPD���$
T;F��DIu)�<I�a\so<"��a-�6Jc6s6�4L��M�V9R�h���T�ri�� ���5�` �f@�@�������P
� �����`��Img PdH�[l��I/A  VP�S��U��Ow��!%S�Skast�dpn)ǲt�� S�WIMEST�BFfe�00��-Q� �_p�PB�_�Rued�_�T�!�_�S ��_bOH573o2c2��-oNbJ5N�Iojb)�	Cdo�cxE��o�_�l p��o�TdP�o�c�B�o r�2.rٱ(Jsp�EfrSEo�f1�}Ξr3 RGoeEL	S��sL����s�� ���B	��S\ $�F�3ryz�ftl�o~�g�o���������?�����P  �n�&�"�l ��T�@<�^�蒐Y��e�u8Z���alib��Γ��ɟ3����埿�\v ��e\c�6�Z�f�T�v�'R VW���8S��UJ91����i�ů[c�91+o�w8���847�:��A4�j���Q��t6�m���vrc.����HR����ot�0ݿ��  d��8ޯ�460�f>eS0L�97��0�U�ЄϦ�60.� g �н�+��'�ܠ�Ϻ��8co��DM߱U"������ߕpi�߲T!� ��na;�� @���u%��ⅰI�loR�d��1a5a9gϱŭ���95����R����1��?��o��#��1A�/���vt{�UWeǟ���ￇ�73[���7�ρ�C3 W��62K�=f	R���8��������d����2�ڔ�����@�@" "http�����t87 �� v R7��78����4�� ��TTPT�#	���ePCV4/v߀�jL�Q�Fa7��$N�0�/2�rIO�)/;/M/N6.sv3�64i�o|S�l? torah?p*�|`�?��AM/�?�
??.?0�k/��1 �JO��� ,O�tro����[P��OB4c.0K?�g'�)�24g?��� (B�Od�\i�OA5sb�?U_�?vAi�/i��/�/Wn��`�o%�Fo�4l�$opf��oXF I)xoΚcmp\7��mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@����naO��4*O0wi��%P�?"�bsg@?�]7�YEM���8wo2VJ�/ե11?o��3DMs�BC��!7J�\���(�52�XFGa AP�ڟ<�v�`/şaqs����'/Of��1�	9�VRK���ph�fքH5+�=�IN/�¤SkiW�/�I�F��_�%��fsH�I�O�l����"<�`���$�`����\jԿ8z5bO�vrouς�93(�ΤH (DϮ� �?sG��|��F�Ou��������D)O��*�3 P$�FӅ�k��ϻ���럴� �PL��ʿ���pbox�ߦeboL���Sh �>�R.�b0wT{����fx6 ��P��D��3��#_&I\m;YEe�OԆ�M�hxW�=Ete,���dct\���O$AkR������Xm*���ro3��D�l��j9��V'�  FC���|@�քy f?6KARE0�_�~ (Kh��.ccf���WpoO�_K�up��a���<H/j#- Eqd/�384���$qu�o�@�/ o2o?Vo<�7C�)�s�NJԆ�|?�3l\sy�?�40�?�Τwio�u]?�w58�?,F�$OJ�
?&Ԇ"io�!�V��u&�A��PR�ߩ5,� s��v1\  H552B��Q21p0R{78P510.R�0  nel �J614Ҡ/WATUP��\d8P545*�H8R�6��9VCAuM�q97PCRImP�\1tPUIF�C8Q2?8  ingsQy0X��4P P63P @P� PSCH��D�OCVڀD �PCS�U���08Q0=PqpV?EIOCr���v P54Pupd�P�R69aP���PSET�pt\hPQ`Qt��8P7`Q�!MA�SK��(PPR�XY���R7B#PO�CO  \pppb36���PR�Q��b�1Pd60Q$cJ53�9.eHsb��v�LCH-`(�O�PLGq\bPQ0t]`��P(`HCR��t4`S�aund�P'MCSIP`e0aPle�5=Ps�p(`DSW � �  qPb0`�aPa��(`PRQ`Tq�RE`(P�oa601P<cPCM�PHcR0@q\j23b�V�`E`�S`UPvisP`E` c�`�UPcPRS	a�bJs69E`sFRDmP�sRMCN:eH9y31PHcSNBARan�rHLB�USM�q�c�Pg52�fHTyCIP0cTMIL�eh"P�`eJ �PA�P�dSTPTX6p967PTEL�p��P�`h�`
Q8P8$Q48>a0"PPX�8P95�P`�[�95qqbUEC�-`F
PUFRhmPfahQCmP90ZQ�VCO�`@PVI�P%�537sQSU�IzVSX�P�SWE�BIP�SHTTIPthrQ62aP�!tP�G���cIG؁�`c��PGS�eIRC�%��cH76�P�e� Q�Q|�Ror��R5�1P s:P�P,t53�=P8u8=Py�C�Q6�]`�b�PI��q52]`sJ56E`s��L�PDsCL�qPt5�7\rd�q75UP c�R8���u5P sR55]`,s� P8s���P�`CP�PP�SJ7]7P0\o�6���cRPP�cR6�ap0�`�QtaT�79P`�364�Pd87]`�d90P0c��=P,����5�9ta�T91P�� ��1P(S���Qpa�i�P06=P- C
�PF�T	���!aLP� PTS�pL�CABR%�I БIQ` ;��H�UPPaintPM�S�Pa��D�IP|�S{TY%�t\patP�TO�b�P�PLSR76�`�5�Q��Wa�NN�Paic�qN9NE`�ORS�`�cwR681Pint'�'FCB�P(�6x�-�W`M�r��!(`OB^Q`plug�`L�awot �`OPI-���PSPZ�PPGڤQ7�`73ΒPRmQad�RL��W(Sp�PS��n�@��E`�� �PTS-�� W��P�`�apw�`��P`cFsVR�PlcV3D%��l�PBVI�SAP�L�Pcyc+PAP�V1�pa_�CCG^IP - U��L�Pwrog+PCCR�`��ԁB�P �PԁK�=�"L�P��p��(h�<�P��h�̱�@g�=Bـ
TX�%�n��CTC�ptp��<2��P927"0ҝP�s2�Qb��TC-�r�mt;�	`#1ΒT�C9`HcCTE�Peurj�EIPp.p/��E�P�c��I�useZ��Fـvrv�F%���TG�P� CP��%��d -h�H-�Tr�a�PCTI�p��T=L� TRS���p��@נ��IP�PTh�Mn%�lexsQTMQ`�ver, �p�SCp:���F��Pv\e�PF�IPSV"+�H�$c�j�ـtr�aCTW8-���CPVGF-��S�VP2mPv\fx����pc�b��e��bV=P4�fx_m��-���SVPD-��SVP]F�P_mo�`V�Z cV��t\��LmP�ove4��-�sVKPR�\|�tPV�Qe5.W`V6�*u"���P}�o`���`��CV�K��N�IIP��CV�����IPN9�Gene���D��D�R�D(����  ��f谔��pos.��inaEl��n��DeR��d�`��d�P��omB���on,���R�D�R��\��TXf��D$b���omp�� "NȔ�P��m���! ��=C-f����=�FXU�����g �F��(��Dt IIД�r�D��u�� "x����Cx_ui 0X������f2��h	Crl2��D,r9�ui�Ԣ� it�2c�0co��e�"����ا(.{)� ���� ﯶ� IQn�Q �I[ ���_= wo���,bD� ���|GG� �����4 ��e� vʷ�� ��&� 2��Z uz������� ��TW�&q~q 5��޷&�o? ;0{��  �2� ��y� ����W&��� ?Ȼ3� A��ew�/> �\�3&�T��� 77߽� ���� �w��� ֵ��&8 �l1���S�) ��{�d *J� �F's ~���� 6:0� ���,��s�- Q��v� ���� �,�T �Z�BLx6���6 ݀�6���Pa�r ��s>�E��j�6dsq��F  ��������ЁDhel������ti-�S�� �Ob��Dbc`f�O�����t OFT��P<A�_�V �ZI��D��V\�qWS|��= dtle�E�an�(bzd��t�itv�Z�z�Ezt XWO H6�6܋��5 H�6H6�91�E4܀TofksqtF� Y682��4�`�f804�E9�1�g�`30oBkmo�n_�E��eݱ�� wqlm��0 J�f�h��B�_  ZD�TfL0�f(P7�EcklKV� �6|�ƁD85��ّ�m\�b����xo�k�ktq��g2.g���y�LbkLVts��IF�bk������I�d I/f��GR8� �han�L�`�Vy��%��%ere�����io�� ac.�- A�n�h��.�cuACl�_�^Cir��)�g��	.�@�& G��R630���p v�p�&H�f���un��R57v�OJavG�`Y���owc��-AS�F��O��7���S�M�����
afN��rafLa�Qvl�\F c�w a�`��?VXpoV �30���NT "L�FFM ��=����yh	a�G-�uw�� �m2.��,�t��̹�6lԯ��sd_�MC'VČ���D���fsl�m�isc. � H552�2��21&dc.pR78�����0�708J�614Vip OATUu�@�OL�w545ҴINTL��6�t8 (V�CA���sse�CRI��ȑ��U�I���rt\rL�2�8g��NRE��.�f,�63!��,�S�CH�d Ek�DO#CV���p��C,�<��L�0Q�isp��EcIO��xE,�54�����9��2\sl,�SET���lр�7lt2�J7�Ռ?MASK��̀?PRXY҇�ҹ7���OCO��J�6l�3�l�� (SVl�A�H�L�@Օn��539Rsv�v��#1��LCH����OPLGf�ou�tl�0��D��HC]R
svg��S@��h��CSa�!�{�50��D�l�5!�lQ��DSW��S����̀���OP����7��P�R���L�ұ�(Ssgd���PCM�Զ�R0 \s��5P՝���0���n�qԋ AJ�1��N�q�2���PRSa���69��� (AuF�RD�Խ��RMC�N���93A�ɐC�SNBA�F9N� HLB��� M���4���h�2A�95�z�HTCaԈ�TM;IL6�j95,��o857.,PA1��ito��TPTXvҴ JK�TEL���piL�� XpL�80�I)��.�!��P;��J95��s "N����H�UEC��77\cs�FR��<Q���C��57\{VcCOa�,���IP1�jH��SUI�	C�SX1�AWE9Ba��HTTa�8�R62��m`��G�P%�IG %tut�KIPGSj�| R�C1_me�H7�6��7P�ws_�+�?x�R51�\�iw�N���H�53�!��wL�8!�h�R66��H���Ԡ�8��@;J56��1�P��N0��9�j��L�F��R5`%�A|�5qԉr�`,�8 5��{16�5!��@�"5��H84!�29��0��P�J���n B[�J377!Ԩ�R6�5h3�n���y36P��3R6 ��-`;о Ԩ@��wexeKJ87���#J90!�stu�+�~@!䬵�k90�kop�B���D�@!�p�@|BA�g*�0n@!��Q��06!�@"[�F�FaP�6��́v,�TS� NC[ЗCAB$iͰl1I��R7��@q�y�wCMS1�rog+Q1M�� �� TY$x�wCTOa�nv\+���1�(�,�6�co�n�~0��15��JNN�%e:��P��9GORS%x���8A�w815[�FCBaUnZQ�P!��p{��C�MOB��"G��O�L��x�OPI�$\�lr[�SŠ�T	D7��U��CPRQR9R	L���S�V�~`����K�ETS�$1��0����3�Ԩ�FVuR1�LZQV3D$� ���BVa�SAP�L1�CLN[�PV��	rCCGaԙ��sCL�3CCRA�/n "W!B�H�7CSKQn\0�pX��)�0CTPn����Qe��p!$bCt�aT0U�pCTC��yЋRC1�1 (<�s��trl,�r��
TX��TCaersrm�r�MC"�sܡ�#CTE��nr5r�REa�XPj�^���rmc�^�a"��P�QF!$���$p� "�rG1�tTG�$c8��QH�$SC�TI�! s��C;TLqdACK�Rpt)��rLa�R82���M��YPk�.���OF ��.���e�{�CN���^�1�"M�^�aԀС�Q`US��!$��M�QW�$m�VGFޑ$R MH��P2�� H5� ΐq���ΐ�$(MH[�VP��uoY����$)��Dv��hg��VPF��"MHG̑`e!�+�V/vpcm�N���p��N��$�VPRqdL)��CV�x�V� `"�X�,�1�($TIa��t\mh��K��eCtpK�A%Y�VP%�ɠ�!PN���Ge{neB�rip�����8��extt���Y�m�"� (��HB���)�� x�������Ȣ�res.�yA�ɠ�n����*���p��@M�_�NĀ6�L���Ș�yAv`L�Xr�Ȉ2��"R;ʎȽ\ra��	P�� 7h86��Gu+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr�Ȩ2��L�1��n2�h� �0XL�XR}�RI{�e� L�x���c�Ș����N�vx�L��"��2\�r�]�N�82�d ���b�ɉa��y1��/��k�@���A��ruk8�ʘ L�sop��H��}�ts{�����sx��9��j965���Sc��h��5 JI9�{�
�PL�J	ween��t I[
.x�com��Fh�L��4 J��fo.��DIF+�6�Q����rati|��p�ڙ1�0�
R8l߾�M �����P��8� �j�mK�X�HZ��$��N�oڠ�ș3�q��vi���890�~�l Sl�yQ���tpk�xb�j �.�@�R�d������,/n(�8�8�0����
:�O8�<�Q}�C�O���PT��O (��.�Xp|�~H���?��v �wv���8�22�pm���7322��j7�^Ϙ@ƙ���cf�=Yv9r���vcu�� �O�O�O�O_#_5_7�93Y_��wv4{_��_w�ʈ�ust_�_�cus�_�Z�� oo,o>oPo�io���nge��(pLy747�jWelʨHM;47ZKEq {����[m�MFH�?�(wsK�8J�n����o��fhl;��wmf���? :�}(�4	<g J{��I�I)̏މw��X�7c74kﭏ/7ntˏ2݊e+���se�/�Caw��8�ɐ��EX �\�!+: �p��~�0e0��nh�,:Mo+�<xO��1 "K�O��\a��#0��.8����{h�L?�j+�mo�n�:��t�/�st�?-�w�:���)�;੬(=h�;
d Pxۻ�{:  ���c �J0��re��}��STD�!�treLAN�G���81�\tq�d�������rc�h.������htwv�WWָ�� R79��"Lo�51 (�I�W�ph�Ո�4�aww�� �vy �62�3c�h a?�ctAi�֘!�X�iؠ�t ��n,�։�����j��"AcJP@�3p�vr{��H�6��!��- S�eT� E3�) G�J�934��LoW�4 (S������ <���91 ��8!4�jA9�所+���y�
��v	�btN�ite{�R ��I@Ո����� P�������	 ����Z�vol��X ��9�0<�I�p���ld*���F�864{��?��K�	�k扐�֘1^�wmsk��M�q�Xa�e�����p��0RBT��1ks.OPCTN�qf�U$ RTCamT��y�� U��y��U��UlU6L�T�1Tx��D��SFq�Ue�6T���USP W�b# DT�qT2h�T��!/&+��TX�U\j6&�U U�UsfdO&�&ȁ�T���662DPN�bi��%�Q�%62V��$���%�� �#(�(6To6eG St�%��#5y��$�)5(To�%tT0�%5�W6T���%�#�#orc��#I��8�#���%cct�6ؑ�?�4\W6965q"p6}"�#\j536����4�"�?kruO O,Im?Np�C ��?t�0<O�;�ea �%���?
;gcJ7� "AV�?�;av�sf�O__&_8WtpD_V_0GT�F|_:U�cK6�_�_r�O�3e�\s�O2^y`O:�m�igxGvgW! m��%��!�%T�$E �A{6�po6��#37N�)5R5_2E���$�0���$Ada�Vd ���V�?;Tz7�_�e7�DDTF9���#8��`�%��4y�ted Z@�A}�@�}�04N�}�}���}�#dc& }����u �6�v��v1�u1\�b�u$2}���}� R�83�u�"}��"}�v�alg���Nrh �&�8�J�Y�o�ue��� j70�v=1���MIG�uerfa ��{q���E�N�ءEYE�ce A���񁏯pV�e�A! ���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b��T��/E In�B�  8W�|��537g��.��(MI�t�Ԇ1r��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y��ac���2���Rɏ �jo��2�� dj�d�8r}� og\�k�0��g��wm�f�Fro/� E�q'�4"}�3 J8��oni[���0�}Ĵ�� o� ��$ʛ��m@�R�e��{n�Д�V�o�������  ����=裆"POS\��<��ͯ menϖ��6��OMo�43��� ��(Coc� An`[�t���"e�a\�v�p��.��cflx$�le��8�hr�trv�NT� CF+�x E/�t	qi�M��ӓxc��p�f�lxX����Z�cx��
0 lh��h8��mo���=� H���)� (�vSER,���g�0߆0\r�vX�= ���I � - �t�i��H��VC�8�28�5��L"�RC��n G/���w��P�y�\v�vm "o�lϚ�x`��=e�:ߠ-�R-3?������vM [�AX/2��)�S�rxl�v#��0��h8߷=� RAX�A�����9�H�E/Rצ�����h߶"RXk��F��˦85��2L/��xB885_�q�R�o�0iA��5\rO�9�K��v����q8���.�n "�v��88��8s�i ?� 9 ��/�$�y O�MS"���&�9�R H74&�`�745�	p��p��y'cr0C�c�hP0� j�-�a%?o��6D9;50R7trl��wctlO�APC����j�ui"�L��� � ����^棆!D�A��qH��&-^7����� λ�616C�q�7914h���� M�ƔI��99��(���$FEAT_�ADD ?	����Q%P  	�H._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������������ &8J\n���������TD�EMO fY   WM _������� �//%/R/I/[/�/ /�/�/�/�/�/�/�/ ?!?N?E?W?�?{?�? �?�?�?�?�?�?OO JOAOSO�OwO�O�O�O �O�O�O�O__F_=_ O_|_s_�_�_�_�_�_ �_�_ooBo9oKoxo oo�o�o�o�o�o�o�o >5Gtk} �������� :�1�C�p�g�y����� ��܏ӏ���	�6�-� ?�l�c�u�������؟ ϟ����2�)�;�h� _�q�������ԯ˯ݯ ���.�%�7�d�[�m� ������пǿٿ��� *�!�3�`�W�iϖύ� ������������&�� /�\�S�eߒ߉ߛ��� ��������"��+�X� O�a��������� ������'�T�K�]� ���������������� #PGY�} ������ LCU�y�� ����/	//H/ ?/Q/~/u/�/�/�/�/ �/�/???D?;?M? z?q?�?�?�?�?�?�? 
OOO@O7OIOvOmO O�O�O�O�O�O_�O _<_3_E_r_i_{_�_ �_�_�_�_o�_o8o /oAonoeowo�o�o�o �o�o�o�o4+= jas����� ���0�'�9�f�]� o���������ɏ��� ��,�#�5�b�Y�k��� ������ş����(� �1�^�U�g������� ��������$��-� Z�Q�c����������� ��� ��)�V�M� _όσϕϯϹ����� ����%�R�I�[߈� ߑ߫ߵ�������� �!�N�E�W��{�� ������������ J�A�S���w������� ������F= O|s����� �B9Kx o������/ �/>/5/G/t/k/}/ �/�/�/�/�/?�/? :?1?C?p?g?y?�?�? �?�?�? O�?	O6O-O ?OlOcOuO�O�O�O�O �O�O�O_2_)_;_h_ __q_�_�_�_�_�_�_ �_o.o%o7odo[omo �o�o�o�o�o�o�o�o *!3`Wi�� ������&�� /�\�S�e�������� ������"��+�X� O�a�{���������� ߟ���'�T�K�]� w����������ۯ� ��#�P�G�Y�s�}� �������׿��� �L�C�U�o�yϦϝ� ���������	��H� ?�Q�k�uߢߙ߫��� �������D�;�M� g�q���������� 
���@�7�I�c�m� �������������� <3E_i�� �����8 /A[e���� ����/4/+/=/ W/a/�/�/�/�/�/�/ �/�/?0?'?9?S?]? �?�?�?�?�?�?�?�? �?,O#O5OOOYO�O}O �O�O�O�O�O�O�O(_ _1_K_U_�_y_�_�_ �_�_�_�_�_$oo-o GoQo~ouo�o�o�o�o �o�o�o )CM zq������ ���%�?�I�v�m� ��������ُ��|�;�  2� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as��������'9  :>Ugy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w����� ����я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ �������(/=C6Y k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ������/�A��$FE�AT_DEMOIoN  E��q���>�Y�INDE�Xf�u��Y�IL�ECOMP g�������t�T���SETUPo2 h����?�  N ܑ���_AP2BCK �1i��  �)B���%�C�>���1�n�E����)� ��M�˯�������<� N�ݯr������7�̿ [��ϑ�&ϵ�J�ٿ Wπ�Ϥ�3�����i� �ύ�"�4���X���|� ��߲�A���e���� ��0��T�f��ߊ�� ����O���s����� >���b���o���'��� K���������:L ��p����5�Y �}�$�H�l ~�1��g� � /2/�V/�z/	/ �/�/?/�/c/�/
?�/ .?�/R?d?�/�??�? �?M?�?q?O�?O<Ot���P� 2�*.VRCO�O�0*�O�O�3�O�O�5�w@PC�O_�0F'R6:�O=^�Oa_�KT���_�_&U�_�\�h�R_�_�6*.F�zOo�1	(SoElx�_io�[STM �b��o�^+P�o�m�0�iPendant? Panel�o�[H�o �g�oYor�ZGIF|��e�pOa��ZJPG ��*��e���z��JJS�����0@���X��%
JavaSc�riptُ�CS�ʏ1��f�ۏ %�Cascadin�g Style ?Sheets]��0�
ARGNAME�.DT���<�`\@��^���Д៍�АDISP*ן���`�$�d��V�e��C?LLB.ZI��=��/`:\��\������Collabo�鯕�	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V� 9���ϝ�$�4i����V���zό�!ߘ�TP�EINS.XML�(�@�:\<����C�ustom To�olbar}��PASSWORD��~�>FRS:\���� %Pass�word Config��?J���C� ��"O��3�����i��� ��"�4���X���|�� ���A���e����� 0��Tf���� �O�s��> �b�[�'�K ���/�:/L/� p/��/#/5/�/Y/�/ }/�/$?�/H?�/l?~? ?�?1?�?�?g?�?�?  O�?�?VO�?zO	OsO �O?O�OcO�O
_�O._ �OR_d_�O�__�_;_ M_�_q_o�_�_<o�_ `o�_�o�o%o�oIo�o �oo�o8�o�on �o�!��W�{ �"��F��j�|�� ��/�ďS�e������ ���T��x������ =�ҟa������,��� P�ߟ񟆯���9��� �o����(�:�ɯ^� ����#���G�ܿk� }�ϡ�6�ſ/�l��� ��ϴ���U���y��  ߯�D���h���	ߞ� -���Q߻��߇��,���$FILE_D�GBCK 1i������� ( �)
�SUMMARY.�DG,���MD:�`����Dia�g Summar�y���
CONSLOG��y����$����Consol�e log%���	?TPACCN���%g�����TP �Accounti�nF���FR6:�IPKDMP.ZIP����
��)�����Excepti�on-����MEMCHECK�������8�Memor?y Data���LN�)�RI�PE���0��%� Pack�et LE���$ySn�STAT*�#� %~LStatus�i	FTP�/��/�:�mmen�t TBD=/� �>)ETHERNE�/o�/�/���Ethern�U<�figura�L��'!DCSVRAF1//)/B?�0� verify �allE?�M(=5DIFF:? ?�2?�?F\8diff��?}7o0CHGD�1�?�?�?LO X�?sO~3&�
I2BO8)O;O�O bO�O�OGD3�O�O�OT_� �O{_
VUPDATES.�P��_��FRS:\��_�]��Upda�tes List��_��PSRBWLOD.CMo���R�o�_9�PS_RO�BOWEL^/�/:GIG��o>_�o��GigE ��n�osticW�N��>�)�aHADOW�o�o�ob��Shadow ?Change���*8+"rNOT�I?=O��N?otific�"���O�A�PMIO�o��h��f/���o�^U�*�UI`3�E�W��{�UI������B���f��_� ������O������� ��>�P�ߟt������ 9�ί]�򯁯�(��� L�ۯp������5�ʿ ܿk� Ϗ�$�6�ſZ� �~��wϴ�C���g� ��ߝ�2���V�h��� ��߰���Q���u�
� ���@���d��߈�� )��M��������� <�N���r����%��� ��[����&��J ��n��3�� i��"�X� |��A�e� /�0/�T/f/��/�/�/=/�/�/�$�$�FILE_�PPR��P��� �����(MDONLY 1i5~�  
 �z/ Q?�/u?�/�?�?t/�? ^?�?O�?)O�?MO_O �?�OO�O�OHO�OlO _�O_7_�O[_�O_ �_ _�_D_�_�_z_o �_3oEo�_io�_�oo �o�oRo�ovo�o A�oew�*� �`����&�O�~�*VISBCK,8|1;3*.VDV�|���FR:\o��ION\DATA�\��/��Vi�sion VD filȅ��&� <�J�4�n������3� ȟW������"���F� ՟�|������m�֯ e������0���T�� x������=�ҿa�s� ϗ�,�>���b��� ϗϼ�K���o��� ��:���^����ϔ��*�MR2_GRP �1j;�C4�  B�}�	 �71������E�� �E�  F@ F�5U�������L���M���Jk�Lzp��JP��Fg�f�?�  S�����9�Y9}��9��8j
��6��6�;֞�A�  ���BmH��B���B���!$����������<���@UUU#��� ��Y�D�}�h������� ��������
C��_CFG k;T M����]�NO :�
F0� � \�R�M_CHKTYP  0�}�00�0��OM_MsIN	x���5v0X� SSBd]l5:0���bx�Y���%TP_DEF_OW0�x�9�IRCO�M��$GENOVRD_DO*�62�THR* �d%d�_ENB�� �RAVCr��mK�� ��� ��/3�/��/�/n�� �M!OUW -s��}��ؾ��8�g�;?�/�7?Y?[?  D�Cý���(7�?�<B�?B����2��*9�.N SMTT#t[)���X}�C�f�HOS�TCd1ux�s��?�� MCx���;zOx� _ 27.0�@1�O  e�O�O	__ -_;Z�O^_p_�_�_�L�N_HS	anonymous�_�_�_oDo1o yO��FhFk �O�_�o�O�o�o�o�o J_'9K]�o �_�����4o� XojoG�~�o^����� ��ŏ�����1� T���y��������� ��,�>�@�-�t�Q� c�u���������ϯ� ��(�^��M�_�q� ����ܟ� �ݿ�� H�%�7�I�[Ϣ�ϑ� �ϵ����l�2��!� 3�E�Wߞ���¿Կ�� ��
�������/�v� S�e�w������� ������+�r߄ߖ� s�����߻������� ���'9K]��� ������4�F� X�j�l>��}�� ����//1/ T��y/�/�/�/�/�.D\AENT 1v�
; P!J/?  ��/3?"?W? ?{?>?�?b?�?�?�? �?�?O�?AOOeO(O �OLO^O�O�O�O�O_ �O+_�O _a_$_�_H_ �_l_�_�_�_o�_'o �_Koooo2o{oVo�o �o�o�o�o�o5�o Y.�R�v���zQUICC0 ���3��t14��"����t2��`�r�ӏ�!ROUTER�ԏ��#�!PC�JOG$���!�192.168.�0.10��sCA�MPRTt�P�!bd�1m�����RT�🟱���$NAME� !�*!RO�BO���S_CF�G 1u�) ��Auto�-started^FTP&�� =?/֯s����0� B��f�x��������� S������,���� �����ϼ�ޯ������ ���ʿ'�9�K�]�o� ��ߥ߷��������� (:~�k�Ϗ� ������������ 1�C�f���y������� �����,�>�R�? ��cu��`��� ��(�$M_ q������  /H%/7/I/[/m/4 �/�/�/�/�/�~/? !?3?E?W?i?��� �?�/�?/�?OO/O �/�?eOwO�O�O�?�O RO�O�O__+_r?�? �?�?�O|_�?�_�_�_ �_o�O'o9oKo]ooo �_o�o�o�o�o�o�o F_X_j_~ok�_� �����o��� 1�TU��y����������U�)�_ERR �w3�я�PDU�SIZ  g�^ڀp���>�WR�D ?r�Cq� � guestb�Q�c�u��������"�SCDMNG�RP 2xr����Cqg�\��b�K� 	P0�1.00 8(q _  �5p�5p�z�5pB  ��{ ���H����L��L��>L�����O8������l�����a4� �x��Ȥ�x��8��U�\���)�`蠍;�������d��.�@�R�ɛ_GR�OUېy���⽒	ӑ���QUPOD  ?u����VİTYg�����TTP_AUTH� 1z�� <!�iPendan䷗-�l���!KAREL:*-�6�H�KC]�m���U�VISION SET���ϴ�g� G�U������R�0�� H�Bߏ�f�x��ߜ߮����CTRL {�����g�
S�?FFF9E3��At�FRS:DEF�AULT;�F�ANUC Web Server;� )����9�K��ܭ����������߄WR_�CONFIG �|ߛ ;��I�DL_CPU_P5CZ�g�B�Dpy�w BH_�MINj��)�}�GNR_IO���g���a�NPT?_SIM_D_������STAL_S�CRN�� ���T�PMODNTOL8������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMAST�E��ɾeSLAV�E ~��c�O�_CFGٱBU�O�O@CYCL�En>T�_ASG� 1ߗ+�
  ����//+/=/ O/a/s/�/�/�/�/���NUM��
�@IPCH�^R?TRY_CNZ��@�@��������1 @kI�+E��z?E�a�P_MEMBERS 2�ߙ�� $���2����ݰ7�?�9a�SDT�_ISOLC  �����$J23�_DSM+�3J?OBPROCN���JOG��1�+��d8�?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSRE�QO��KANJI_����a[�MONG ����b�yN_ goyo�o�o�o�Y�`3	�<� ��e�_ִ���_L���"?`EY�LOGGINL�E�������$L�ANGUAGE Y��<T� {q��LGa2�	�b����g�xP��  *��g�'��b����>�MC:�\RSCH\00�\<�XpN_DISP �+G�J��O��O߃LOCp�D�z���AsOGB?OOK ����`��󑧱����X� ����Ϗ����a�*��	p������!�m��!���=p_B�UFF 1�p��2F幟���՟�D� Collaborativǖ ���F�=�O�a�s��� ����֯ͯ߯����B�9�K���DCS ��z� =��� '�f��?ɿۿ���H@�{�IO 1��# ~?9ü��9�I� [�mρϑϣϵ����� �����!�3�E�Y�i� {ߍߡ߱��������-E��TMNd�_B� T�f�x�������� ������,�>�P�b��t�������L��SE�VD0��TYPN1�$6���Q�RS"0&��<2FLg 1�"�J0��� �����G�TP:pOF�NGNAM1D�mr�t7UPS�GI"5�a�O5�_LOAD�N@G %�%��pIND�`5SE�� ��$MAXUALRM�'���(��'_PR"4F0d��1��B_PNP� V� 2�C	M�DR0771ߕz�BL"8063%�@ �_#?�ߒ|/�C��z�6��/􈃟/Po@P 2���+ �ɖ	~T 	t  ��/ �%W?B?{?�k?�? g?�?�?�?O�?*OO NO`OCO�OoO�O�O�O �O�O_�O&_8__\_ G_�_�_u_�_�_�_�_ �_o�_4ooXojoMo �oyo�o�o�o�o�o �o0B%fQ�u �������� >�)�b�M�����{��� �����Տ��:�%��^�p�S�������D�_LDXDISA�pB�MEMO_{APjE ?C
 �,�(�:��L�^�p������IS�C 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%� �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A����??��4[���ཌ���qϿ��j]�Q_D���^�PL_NA_ME !3%,��!Defau�lt Perso�nality (�from FD)� �RR2� 1��L6(L?y�,0	l d� �������/ /(/:/L/^/p/�/�/@�/�/�/�/�/ZX2u ?0?B?T?f?x?�?�?�?�?\R<?�?�?O  O2ODOVOhOzO�O�O\�OZZ`\R�?"�N
�O_\TP�O:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHo_ )_~o�o�o�o�o�o�o �o 2DVhz �[omo����
� �.�@�R�d�v�����𬏾�Џ� E�f  Fb� F�7���   ��!��d��@�R� 6�t������l���pʝ����� ݘ ����"�@�F�d����� "𩯹�ݐA�#  ϩU[�$n��B�E ��� � @D7�  �?�� ��?�@��A@�;f���FH� ;�	l>,�	 |��j�ys�d�>���� ��� K(��K�d$2K ��J�7w�KYJ˷�ϜJ�	�ܿ��� @I���_�f�@�z���f�γ�N��}����	Xl��������S��ĽÔ��I �����5���  �����A?oi#��;��A��� o���l� �π��-���ܛG�G�Ѳ���@n�@a �  �  ���ܟ*�͵	'�� � H�I� �  �Р�n�:�Èl�È�=��̈́�в@�ߚЕ����/������̷NP� � ',���-�@�
�@���?�=�@A���B� � Cj�a�Be�Czi��@#�B�޸�ee��^^ȹBР��P��`��̠�����ADz՟ �n�3��C�i�@�R�pR�Yщ��  �@O� ��Ż���?�ff������n� ɠ#ѱy9�G
(���I�(�@uP@~����t�t���>�����;�Cd;���.<߈<�g�<F+<L�������,�d�,�̠�?fff?��?&�&��@��@x���@�N�@�?��@T�H�� ��!-�ȹ�|�� 
`�������/ /</'/`/r/]/�/��eF���/�/�/�/@m?��/J?�(E���G�#�� F Y�T?�?P?�?�?�?�? �?O�?/OO?OeOk� ��O�IQOG�?�O1?��OmO_0_B_T_������A_�_	_�_P�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�ol�o���W�����o;C�E� q�H�d��؜a@q��e��F�BµWB]��NB2�(A����@�u\?��D�������b�0��|�uR�����
x~�ؽ���Bu*C���$�)`�$ ����GC#����rAU�����1�eG��D�I�mH��� I:�I��6[F���C��I��J�:�\IT�H
~�QF�y��p���*J�/ I8�Y�I��KFjʻCe�o��s��� ��Џ���ߏ�*�� N�9�r�]��������� ���۟���8�#�\� G�����}�����گů ���"���X�C�|� g�����Ŀ������ �	�B�-�f�Qϊ�u� ���ϫ��������,� �P�b�M߆�qߪߕ� �߹�������(��L� 7�p�[����������s($���3:�����$���3���d�,�4��x@�R��񴲚�l�<~�wa���e����wa4 �{����@��(L:ueP�	P~�A�O�������	���� G2W}h� �����/�� �O�O7/m/[(d=�s/ U/�/�/�/�/�/?�/�1??U?C?y?�=  �2 Ef9gFb-��77�9fB)aa�)`C9A`�&`w`@ -o�?9de�O-OOQOpn�?�?�O�O�O�O�9c?�0�A7ht4Rw`w`!w`xn
 �O9_K_]_o_ �_�_�_�_�_�_�_�_po#ozzQ ��h���G���$MR�_CABLE 2}�h �a:�T� @@�0�A�e��a�a�a��`���0�`C�`�aO8��tB����bo}GT D�D�F��o�f�#��0���0�DO���`����0��CbD�%���o�h8  ����C�07�d�4�`���P�}�T D��R"�4��`y`By`C\�p�bHE��`�,�w��И5D��#z�lҠ`��0�q�pήb0��abr3E}�T D�R��y /o�c-���H� �2��� V�����������'��"���D���^q��o <�\���������������*,�**} \cOM �ii�����r���%% 23456�78901i�{� �f�����������1�����
��`��not sen�t 5���;��TESTFECoSALGupeg`���1d.�š
:��� �DCbS�Q�c�u���� 9UD1:�\mainten�ances.xm�l��ֿ�`Z�DEFAULT-���4\bGRP 2��M�  =�U[ � �%Forc�e�sor ch�eck  �����Bz��p����h5-���ϻ��������%!�1st clea�ning of cont. v�ilation��}�Rߗ+��[�ߔ��߸���mec�h�cal`�������0��h5 k�@�R�d�v����(�rolle_Ƶ����/���(�:��L��Basic� quarterCly�������,������������MH��:(�"GpP(�X_h5�������#C���M"��{Pbt����Suppq�greasq� ��?/&/8/J/\/���C+ ge��. batn�y`/��/h5	/�/�/�/? ?X_�ѷen'�v��/�/��/��?�?�?�?�?�G=?O�aEp"CrB1O��0�/ `OrO�O�O�O�t$��Lf��C-(��A�O:�OO$_6_H_Z_l_z�t*cabl�O(���S<(��Q�_:�
_�_�_oo0o@o)(Ӂ/�_�_���_��o�o�o�o�o�O�@hau1�l��2r x(�<qC:���op������R/eplaW�fUȼ2�:�._4�F�X�j�|�(�$%���ߟ�� ��#���
��.�@��� d���ŏ׏����П� ���U�*�y�����r� ��������	�q��?� ߯c�8�J�\�n���ϯ �����ڿ)����"� 4�Fϕ�jϹ�˿��� ���������[�0�� ��fߵϊߜ߮����� !���E�W�,�{�P�b� t����߼����� A��(�:�L�^���� ����������  $s�H������q� ����9]o �Vhz���U �#�G/./@/R/ d/��/�/��//�/ �/??*?y/N?�/�/ �?�/�?�?�?�?�??? Oc?u?JO�?nO�O�Op�O�O+Jkb	 H�O �O__6M2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�op*<ND@ �bA�?�  @!Q _���Fw��� �H* �** @A>F�pRT�f��x�:�������ҏ��eO^C7�Տ#�5�G� 	�k�}���ُ���c� ����W��C�U�g� ��ß)�����ӯ��� 	��-�w�����9��� ����m�Ͽ��=�O��E!Q�$MR_HIST 2�>E}N�� 
 \
B�$ 2345678901^�f�#��]�9O���φϸ� O�)�;����q߃� ��L�^߬����ߦ�� ��7�I� �m�$��� Z���~������!��� E�W��{�2�����h������:�SKCFM�AP  >E�Q��r5�!P�����ONREL  .�3���EXCFENB8q
��QFNCX�JJOGOVLI�M8dNá ��KE�Y8��_P�AN7����RU�N����SF?SPDTYPxC���SIGN8JTO1MOT�G���_CE_GRP 1�>EV��@ �����/Ⱥ� �/�/U//y/0/ n/�/f/�/�/�/	?�/ ???�/c??\?�?P? �?�?�?�?�?O)OO�MO,���QZ_ED�IT5 )TCO�M_CFG 1����[�O�O�O 
>�ASI �y3�!
__+[_O_ċ�>O�_bHT_/ARC_U.Ń	�T_MN_MOD�E5�	UAP�_CPL�_gNO�CHECK ?^�� �� o .o@oRodovo�o�o�o �o�o�o�o*!�NO_WAIT_�L4~GiNT�A���EUwT_ERMRs2���3��Ʊ J�����>_)�V�|MO�s��}x:O�v���8�?������ l��rPA�RAM�r�����j���5�5�G� = ��d�v�~�X� �����������֟�0����b�t������SUM_RSPACE�����Aѯۤ��$ODRDSP��S7cOFFSET_CARt@�_��DIS��PEN_FILE:�7�A�F�PTION_�IO��q�M_P�RG %��%$�*����M�WORK� �yf C��춍���  '� �������G	 ������It���RG_DS�BL  ��C��{u��RIENTkTO7 �C� �A �UT_S/IM_Dy����V�LCT ���}{B �٭��_P�EX�P=��RAT��W dc��UOP ���`����e�w�]ߛߩ��$��2r�L6(�L?���	l d������&�8� J�\�n������� �������"�4�F�X���2�߈���������@����*�<w� Tfx��������J` [ˣG���Tz��Pg������ /"/4/F/X/j/|/�/ �/�/���/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?�/�/,O>O PObOtO�O�O�O�O�O �O�O__(_:_��O���y_�]2ӆ� �_�^�_�_�W^]^]��/ooSog��Hgro hozo�o�o�o�o�oF`��#|`�A� � 9y����OK�1��+k�+�����<�E�A�nq @D�C  �q����nq?���C��s�q1� ;��	l��	 �|�Q�s�r�q>���u
��qF`H<�zH~�H3�k7GL�zH?pG�99l7�0k_B�T�F`C4��k��H���t��-�Ae����k�����~s���  �ሏ�����EeBVT����dZ=���ڏ ���q�-�Fk�y�{FbU��= n@6�  ���z�Fo���Be	'� � ���I� � � �:p܋=��q�ڟ웆�@�@��B�,���B����g�AgN����  '�|���g��B��
p�BӀC׏����@?  #�Bu�&��ee�^^މB:p2���>�m�06p�Z�=Dz?o}� ܏������׿�������Ǒ��� f�  ȧ �M���*�?��ff�_8�J�ܿ !3pϑ�ñ8= �ϐ�ʖq.·�(= ��P@���'��s�tL�>���/�;�Cd;���.<߈<�g�<F+<L ��^oiΚrd@��r6p�?fff?�?&��п�@��@x���@�N�@�?��@T싶�Z ���ћtމ�u�߈w	� x��ti�>�)�b�M�� q����������� ��:�%�^�������W����S�E�  G}�=F�� Fk� ��������1U@ yd������q ��	��{�A��h@�����a��ird��A{/w/J/(5/n/	�A��A���":t�/ C^/�/Z/ ލ?���/�/1?,?���W����g��pE� ~1�?0�4�0
1�1@I�Ӏ��BµWB]��NB2�(A���@�u\?����������b��0�|�uR�����
�>�ؽ���Bu*C��$�)`�?� ���GC#����rAU�����1�e�G���I�mH��� I:�I��6[F���C�4OI��J��:\IT�H
?~QF�y�Ol@��*J�/ I�8Y�I��KFjʻC��-?�O�O __>_)_b_M_�_�_ �_�_�_�_�_o�_(o o%o^oIo�omo�o�o �o�o�o �o$H 3lW�{��� ����2��V�h� S���w�����ԏ���� ���.��R�=�v�a� ������П����ߟ� �<�'�`�K�]����� ����ޯɯ��&�8��#�\��3(J���3�:a������J�3Ï�c4�����������������xڿ�n����e�<�n�4 �{2�2ɀr�`ϖτϺϨ��%PR�P���!�h��!�K�6�o�Z�����u�|ߵߠ������� ���3��W�B�{�f�@4���������d�A ����!��1�3�E�{��i������������� � 2 Ef�7F[b�7��6B�!,�!� C9� �� n�@�/`r������#x��+D=�3?, V�8v�n�n��n��.
 D��� ��//%/7/I/[/�m//�/�:� ���ֻ�G���$P�ARAM_MEN�U ?2���  �DEFPULSE��+	WAITT�MOUT�+RC�V? SHE�LL_WRK.$�CUR_STYLv� 4<OPTJNJ?PTB_?Y2C/?R_DECSN 0 �Ű<�?�?�?�?�?O O?O:OLO^O�O�O�O��O�O�!SSREL?_ID  .�����EUSE_PR_OG %�*%�O0_�CCCR0�B���#CW_HOST !�*!HT�_=ZAT��O_�Sh_zQ�S|�_<[_TIME
2��FXU� GDEB�UG�@�+�CGINP_FLMSKo�5iTRDo5gPGA�b` %l�tkCH�Co4hTYPE�,� �O�O�o#0 Bkfx���� �����C�>�P� b���������ӏΏ�� ���(�:�c�^�p������7eWORD �?	�+
 	�RSc`n�PNS2��C4�JOv1���TE�P�CO�L�է�2��gLP �3��n��OjTR�ACECTL 1�2��! .��m n����|��q�DT Q�2��Ǡ��D � _: Ԡؤؤ��ڢׯ� ����1�C�U�g�y����������ӿ���':�����X}`���1�<���&�@.�K�uJ�qJ�H�EH�	H�?�K�H�UH�H�H�H�T�@J�H�H�H��E�W�i�{ύϟϰ�������;��a�ߞ߰����� ���'��������� ������'���/��� 7���?���G�3�ݿ� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������С �*<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6@ubt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀�V�߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z?��?�?�?�?�1�$P�GTRACELE�N  �1  ����0���6_UP �����A@�1�@�1_CFG ��E�3�1

@�<D�3UOaHSO��0$BDEFSPD� �/L�1�0���0H_CONF�IG �E�3� �0�0d�D�&�2 �1�APpDsAl�A�0��0IN'@?TRL �/MOA�8pEQPE�E��G�A<D�AIWLID(C�/M	bT�GRP 1ýI� l�1B � �����1A��33FC� F8� E�� @eN	�A�AsA�Y�Y�A�@?� 	 vO�Fg�_ ´8cokB;`baBo,o>oxobo��o�1>о�?B�/�o�o~�o =%<��
 C@yd��"�������  Dz@�I�@A0�q� � ������ˏ���ڏ� ��7�"�4�m�X���|����Ú)ґ
V7�.10beta1�HF @�����Aq��Q�  �?� �B���P�p �C��~&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@p���f������ҡr�R�ܣ�Rљ����1�i�������t<B!CeQKNO?W_M  lE7F�bTSV ĽJ�BoC_�b�t��������������1�]aSM��SŽK ���	�NB�0����ĿK���-�bb��A�RP���`�0�Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1=�K
 4MU�iǨj� K�]�oߠ� �ߥ߷�������2�� #�h�G�Y��}������
������,�2r7�I��1�<t�H��P3^�p�����,�A4��������,�5(:,�6Wi{�,�7����,��8�!3,�MA�D�6 F,�OV_LD  KD��xO.�PARNUM�  ��C/%�S+CH� E
9'!8G)�3Y%UPD/���E�/P�_CMP_0��0@�0'7E�$�ER_CHK�%05H�&�/�+RS����bQ_MO�+?=5_�'?O�_RES_G6��:�I�o�?�?�? �?O�?O7O*O[ONO OrO�O�O�{4]��<�?�Oz5���O__ |3 #_B_G_|3V b_ �_�_|3� �_�_�_|3 � �_�_o|3Oo>o<Co|2V 1�:�k1�!�@c?�=2T?HR_INRc0i!�}�o5d�fMASS6�o Z�gMN�o�c�MON_QUEUE �:�"�j0��Ut4N� U1Nv�+DpENDFqd?`y�EXEo`u� BE�npPAsOPTIO�Mwm;DpPROGR�AM %$z%�Cp}o(/BrTASK�_I��~OCFG� �$��K�D�ATA��T���j12,ź�̏ޏ�� ���&�8�J�\�n���������ȟ{�INFO�͘��3t��!� 3�E�W�i�{������� ïկ�����/�A�@S�e�w�����Θ�a '��FJ�a K_N���T��˶ENB�g ڽw1��2��G�N�2�ڻ P(O�=���]�ϸ�@���v� ��u�uɡdƷ_E?DIT �T���|��G�WERFL�x��c)�RGADJ {Ҷ�A�  $Ձ?j00��a�Dqձ���5�?�D�ʨ�<u�j0�%e`������FӨ�2�R�V�	H;pl�G�b�_�>�pAod�t$��*�/� **:�j0�$�@킆5Y�T���^��q �߈b~�L��\�n�� ������������ ��4�F�t�j�|����� ��������bL BT�x���� :��$,�P b���/��� �/~/(/:/h/^/p/ �/�/�/�/�/�/V? ? ?@?6?H?�?l?~?�? �?�?.O�?�?OO O �ODOVO�OzO�O_�O �O�O�O�Or__._\_ R_d_�_�_�_�_�_�_�f	g�io�pWo�o{d �o�~o�ozo�B�PREF ��Rږp�p
�IOORITY�w[���MPDSP�q��pw�UT6����ODU[CT3���v��OG��_TG���8��ʯrTOENT� 1׶� (!AF_INE�p�,�7�!tcp|7�_�!udN�~��!icmv���ޯrXYK�ض���q)� ,�����p��&�	��R� 9�v�]�o�����П�������*��N�`�*�sK��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b��t����u�w�HANCE �R��:�Bwd��连�2s�9�Ks��PORT_WNUM�s�p����_CARTR�EP{p�Ω�SKS�TA�w d�LGmS)�ݶ��t���pUnothing�������{��TEMP ޾y���'e��_a_seiban�o\��o lߒ�}߶ߡ������� ��"���X�C�|�g� ������������� 	�B�-�f�Q���u��� ����������, <bM�q��� ����(LٟVERSIyp�w�} disa�bledWSAV�E ߾z	2600H768S	?�!ؿ�����/ 	5(�r)og+^/y�e{/�/�/�/�/"�*�,/? �p����_�p 1�Ћ�� ������Wh?z?�W*pURG�E��B�p}vgu,�W�F�0DO�vƲ�vW�%��4(�C�WRUP�_DELAY ��\κ5R_HOT %Nf�q׿GO�5�R_NORMAL�&H�r6O�OZGSEM�IjO�O�O(qQSKKIPF3��W3x= _98_J_\_]�_�_ {_�_�_�_�_�_�_	o /oAoSoowoeo�o�o �o�o�o�o�o+= aOq���� ����'��7�]��K�������)E�$R�A{���K/�zĀ~Á_PARAM�A�3��K @.�s@`�61�2C<�5�y��C�6$�=BÀBTIF�4`�RCVTMOUu��c��ÀDCR�F3��I ��+QB�s�D��ߚD�J:��ϗ9±"Z¹{�ޅ��_�1��J��_��k_ �;�Cd;���.<߈<�g��<F+<L�A��Ѱ��d�u�L� ������ϯ�����)�;�M�_���RDI�O_TYPE  �M=U�k�EFPO�S1 1�\�
 x4/�œS����0� )/T��x��uϮ�I� ��m��ϑ�ߵ����� �t�_ߘ�3߼�W��� {�����:���^��� ���/�A�{����� � ��$���H���E�~�� ��=���a������������D/h��S2 1�KԿX��T�x��3 1� ����nY�S4 1�'9K��/�'/�S5 1���/�/�/|�/:/S6 1�Q/�c/u/�/-??Q?�/S7 1��/�/
?D?��?�?�?d?S8 1�{?�?�?�?WOBO{O��?SMASK 1�L��O�D�GXN�O���F&�^��MOCTEZ�Ż��Q_ǁ��%]pA݂��PL_RANG!Q]�_QOWER �ŵ��P1VSM_DRYPRG %ź�%"O�_�UTART� �^�ZUME_PRO�_�_4o���_EXEC_EN�B  J�e�GS�PD`O`WhՅjbT3DBro�jRM�o�h�INGVERSI�ON Ź�#o�)I_AIRPURhP �O(�M�MT_�@T�P#_�ÀOBOT_ISOLC�NTVő'q�huNAME�l���o�JOB_ORD_NUM ?�X�#qH76�8  j1Zc@n�r
�rV�sw��r�?�r�?�r�pÀPC�_TIMEu�a�x�ÀS232>R1��� LTE�ACH PENDcANw�:GX��!O Maint�enance C�onsj2����"���No UseB�׏������1�8C�y�V�NPO�P@��YQ�cS�C7H_L`�%^ ��	ő��!UD�1:럒�R�@VA#IL�q@�Ӏ�J�Q�SPACE1 2�ż ��YRs�i�@Ct�YRԀ'{��?8�?��˯ ����"���7�2�c� u�����G���߯ѿ� ���(��u�AC�c� u�����Ͻ�߿���� ���(��=�_�qσ� ��C߹������߱�� $��9�[�m�ߑߣ� Q������߭��� ��� 	�W�i�{���M��� ����5���.S� e�w�����I����� ��*?as ��E����� /&//;/]o�� ����/2/�/?"? �/7?Y/k/}/�/�/O? �/�/�?�?�?O0OO~KA��*SYPp�M*�8.302�61 yB5/21�/2018 A� �WPfG|�H�_�TX`� !$C�OMME��$USAp �$ENABLED�Ԁ$INN`QpI�OR�B�@RY�E_�SIGN_�`�AP��AIT�C�BWRKz�BD<�_TYP�CRINDXS�@W��@%VFRI{�_G�RPԀ$UFR�AM�rSRTOOL�\VMYHOL�A�$LENGTH_�VTEBTIRST��T  $SE�CLP�XUFINV�_POS�@$�MARGI�A$�WAIT�`�ZX2l�\�VG2�GG1�AAI�@�S�Q	g�`_WR��BNO_USE_�DI�BuQ_REQ��BC�C]S$CUR_TCQP�R"a^f� �GP_STA�TUS�A @ ��A3`�BLk�H$�zc1�h�P@���@_��FX �@E_MLT_CT�C�H_�J�`CO�@O�L�E�CGQQ$W��@w�b#tDEA�DLOCKuDELAY_CNT�a�3qGt�a$wf �2 R1[1T$X<�2[2�{3[3$Zwy�q%Y�y�q%V0�@�c�@�b$V�`�R�V�UV3oh>b�@� � �d�0arMSKJ�LgWaZ�C`�NRK�PS_RATE�0$���S
`�Qv�TAC��PRD��$�e�S*��a4�A�0:�DG�A 0�P�f�lp bquS2�ppI�#`
`�P 
��S\`  ؾA�R_ENBQ ��$RUNN�ER_AXI�<`A�LPL�Q�RU�THI�CQ$FLIP�7��DTFEREN|��R�IF_CHS�U�IW��%V)�G1�����$PřA�Q�Pnݖ_JF�PR_P��	�RV_DA�TA�A  =$�ETIM���_$VALU$�	��OP_   ��A  2 ��SC*�	�� �$ITP_0!�SQ]PNPOU}�o��TOTL�o�DSP>��JOGLIb��P'E_PKpc�Of�i���PX]PTAS��$KEPT_MI�R��¤"`M�b�A	Pq�aE�@�y�q��g@١c�q�PG�BCRK6�x���L�I��  ?�SJ�q�P��ADEz�ܠBSO�Cz�MOTNv�D�UMMY16Ӂ�$SV�`DE_O�P��SFSPD_�OVR
���@L�D����OR��TP8�LE��F������OV��SF��F����bF�d�ƣ&c)�fQ~c�LCHDLY��RECOV���`���W�PM��gŢ�ROȲ�����_F�?� �@v�S �NVER\�@�`OFS�PC,�CSWDٱc�ձ���B,����TRG�š�`�E_FDO��MB�_CM}���B��BALQ�¢	�Q�̄VzaF�BUP�g��G
��AM���@`KՊ�fe�_M!�d�AMf�<Q��T$CA����uDF���HBKd��v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�Dd�9�1A��9�3A�^��ATIO�0���͠��US����WaAB��R+c�`tá`Dؼ�A��_AUXw�S�UBCPUP���S �`����3Եжc����3�FLA�B�HW�_Cwp"�Ns&�]sA�a��$UNIT�S�M�F�ATTR�Iz�Z�CYCL��CNECA���F�LTR_2_FI~��TARTUPJp0����A��LP����ޖ�_SCT*cF_�F�F_P���b�FS8��+�K�CHA/Q��p*�d�RSD��`Q����Q���_TH��PROr���հEM�PJ���G�T�c �Q�DI�@~y�RAILAC/��bMX�LOf�xS���ځ���拁���P�R#�S`app�C�� 	��FUsNC���RIN``QQP� ԱRA)]R ��AƠ��AgWAR֓��BLZa�WrAkg�ngD�AQ�B�rkLD@�र&q�M�K����TI���j���$�@RIA_SWV��AF��Pñ#���%%�p9r1��MO9IQ���DF_~P(��PD"LM-�FA��PHRDY�DORG�H; _QP�s%MULSE~Pz���**�� J��Jײ���FAN_ALMsLVG��!WRN�%�HARDP��UcO��� K2$SHADOW]�kp�a02��N� STOf�+�_^�w�AU{`R��eP_SBR�z5���:�F�� �3MPIN�F?�\�4��3R3EGV/1DG�+c1Vm �C�CFL(��?�DAiP���Z`Ɨ� �����Z�	 ��P(Q$�A$�Z�Q V�@�[�
7� ��EG��o����kAAR���㌵2p�axG��AXE��wROB��RED���W�QD�_�Mh�SY�A��AF��FS�GWRqI�P~F&�STR��(��E�˰EH�)��D�a\2kPB6P��=V���Dv�OTO�1)���ARYL�tR��v�3���FI&�ͣ$LINKb!\��Q%�_3S���E�N�QXYZ2�Z5�V'OFF���R�R�X%xPB��ds�G�cFI�03g�h������_J���'�ɲ�S&qR0LTV[6����aTBja�"�bCL���DU�F7�TUR� X��e�Qb�2XP�ЊgFL�@E���x@�`�U9Z8��^�� 1	)�K��	Mw��F9��劂����ORQj��G;W3���#�Ґd ���upz����1�tOVE�q_�M��ё?C�uEC�u KB�v'0�x-�wH��t ���& `��qڠ� B�ё�u�q�wh�ECh�L���ER��K	�!EP����AT�K�6e9e�W���AXs�'��v�/�R  ����!�� ��P ��`��`�3p�Yp�1�p�� �� � � (�� 8�� H�� X� � h�� x�� ������oDEBU�$`%3�I��·RAB�ȱ�ٱ�sV��� 
d�J、��@񘧕� ������Q���a���a ��3q��Yq+$�`%"<�.cLAB0b�u��'�GRO���b<��B_s��"Tҳ*`��0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθu�ݸ��PNT0����SERVE �Z@� $`EAV�!�PO����nP!��P@�$!Y@ w $>�TRQ�b�
=��BG�K�%"2�\��� _ � l��5�D6ERRVb(�I��V0`;���'TOQ:�7�L�@
�(R��e G�%�Q��q <�50F� ,��`�z�>�RA� �2 d!�����S�  M��px�U ����OCuG��  ��COU�NT6Q��FZN_wCFGF� 4#��6��TG4�_�=�����(���VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@H�EL�0��� 5b`B_BASN��RSR�6�C�SH����1�Ǌ�2���3��4��5��6ʭ�7��8��}�ROaO����P�PNLEAƭcAB)ë ��AC-Ku�INO�T��(B�$UR0� =�_P�U��!0��OU+�P�d�8j��� V��T�PFWD_KAR���� ��RE(ĉ P��P�>QUE�:RAO�p�`r0P1I� �x�j�P�f��6�QSCEM��0��� A��7STYL�SO j�DIX�&�����S!�_TMCMANR�Q��PENDIt�$KEYSWIT�CH���kHE��`BEATM83PE{@LE��>]���U��F��SpD_O_HOM# O�6@�EF�pPRaB(�A#PY�C� O�!���OV_M|b<0 �IOCM�dFQ�1�h�HKYA �D�Q�7��UF2��M����p�cFORC��3WAR�"�OM>|@  @S�#�o0U)SP�@1�2�&3&4E���T�O���L���8UN�LOv�D4K$ED�U1  �SY�HwDDNF� M��BLOB  p��SNPX_AS�� 0@�0��81�$SIZ�1$�VA{���MULTKIP-��# A� � $���� /4`�BS��0�C<���&FRIFBO�aS���3� NF�ODBUP߰�%@3�;9(��ҋ�Z@ x6��SI��TEs�r.�cSGL�1T�Rp�&�Н3B��@�0ST�MTq�3Pg@VByW�p�4SHOW�5n@�SV��_G��; 3p$PCJ�PЬ����FB�PHS�P AW�EP@VD|�0WC� ���A00��PB XG �XG XG$ XG5VI6�VI7VI8VI9VIAVIBVI�XG�YF�0BXGFVH��XbI1oIU1|I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1YU1Y2UI2bI2oI2|I2�I2�I�`�XP�I2p�X�I2�I2�IU2�I2�I2Y2Y��p�hbI3oI3|I3��I3�I3�I3�I3��I3�I3�I3�I3��I3�I3Y3Y4��i4bI4oI4|I4��I4�I4�I4�I4��I4�I4�I4�I4��I4�I4Y4Y5��i5bI5oI5|I5��I5�I5�I5�I5��I5�I5�I5�I5��I5�I5Y5Y6��i6bI6oI6|I6��I6�I6�I6�I6��I6�I6�I6�I6��I6�I6Y6Y7��i7bI7oI7|I7��I7�I7�I7�I7��I7�I7�I7�I7*�I7�I7Y7T�kVP� UD�y"Dՠ��
<A62��ut�R��CMD� ���M5�Rv�]��Q_h�R���e�����<�YSL���  � �%\2��+4�'���W�BVALAU��b��'���FH��ID_L���HIr��I���LE_���㴦�$0C�SA~C�! h �VE_BLCK���1%�D_CPU 5ɧ 5ɛ �����C��� ��R " � PWj��#0��LA�1SBћì����RUN_FLG �Ś����ĳ �����Ą����H���Х�"ށTBC2��# � @ B��e ��S�8=�FTDC����V���3d�Q�CTHF�����R�~L�ESERVE9��F��3�2�E��о��X -$��L�EN9��F��f�R1A��W"G�W_5�b�i1��д2�MO-�T%S60U�Ik�0�ܱ0F����[�DEk�21�LACEi0�CC8S#0�� _MA� j�8��z��TCV����z�T�������.Bi�'A�z�'AJh�#EMD5���J��@@i�V�
z���2Q �0&@o�lh��JK��VK9`��{���щ�J0�����JJ��JJ��A�AL���������42��5�ӕ N1����(���.�LD�_�1�* �CF�"% =`�GROU���1��AN4�C�#m R�EQUIR��E�BU�#��6�$Tk�2$���zя �#�& \�APP�R� C� 0�
$O�PEN�CLOSD�St��	i�
�.�&' �MfЩ�8��W"-_MG�7�CB@�A���BB{RK@NOLD@>�0RTMO_5ӆ$p1J��P��� �����������a6��1�@ )!|�#�(� ������'��+#PATH''@!6#@!�<#�� � '��1SCA����6IN��U�CJ�[1� C0@UM�(Y ��#�"�����*���*��� PAYL�OA~J2LؠR'_AN^�3L��9�1�)1AR_F2gLSHg2B4LO4��!F7�#T7�#ACRL_�%�0�'�$��9H��.�$HA�2�FLEX��J!�) P�2�D߫�����0��* :����z�FG]D����0z���%�F1]A�E �G4�F�X�j�|���BE����������� �(��X�T*�A���@@�XI�[�m�\At�T$g�QX<�=��2TX�� �emX�������������������+	�J>+ �-�K]o�|�٠AT�F�4�E�LFPѪs�J� *v� JEmCTR�!��ATN�vzHA_ND_VB.��1ܝ�$, $8`F24Av���SWu	#�-� $$M *0.�]W�lg��PZ����A��� 1��D��:AK��]AkAAz��LN�]Dk�DzPZ G��C�S�T_K�lK�N}DY��� A����0�� <7]A<7W1�'��d�@g`�P��������"
"J"�. M�2D%"��H����OASYMj%0�� Bj&-��-W1�/_� {8� �$�����/�/�/�/ 3J<�:9��/�89�D_VI��v����V_UNI�ӛ��cD1J����� ��W<��n5Ŵ�w=4�@�9��?�?<�uc�4��3�%�H���a/�j��0�DIz�uO���k�>S0 �`��I��A� �#���@ģ���@����IPl� 1 � -/�ME.Qp��49�ơT}�PT�;pG �+ Gt� ����'��T�0 $DUMMY1���$PS_�@RF��@  G b�'FLA@ YP(c|��$GLB_TP� ŗ���9 P�q���2 X� z!ST�9�� SBRM M�21_V�T$S/V_ER*0O�p�Ӧ��CL����AGPOl��f�GL~�EW>��3 4H �$Y
rZrW@�x�A1+��A���"	""�U&�4� 8`NZ�"�$�GI�p}$&� �-� �Y�>�5 L�H {��}$F�E^��NEAR(PN�CyF��%PTANC�B�	!JOG�@� �6.@$JOIN�Twa?pd�MSET.>�7  x�E��HQ�tpS{r��up>�8׼ �pU.Q?��� LOCK_FOxV06���BGLV�s�GLt�TEST_sXM� 3�EMP�����_�$U&@%�w`24� Y��5��2�d��3��C�E- ���� $KA�R�QM��TPDRqA)�����VECn@���IU��6��H=Ef�TOOL�C2�V�DRE IS3�ER6��@ACH� 7?Ox �Q��29Z�H I� � @$RAIL_�BOXEwa�R�OBO��?��HOWWAR�1�_�zROLMj��:q�w�jq� �@ O_=Fkp! d�l�>�9�� �R OB8B: �@�c�KOU�;�Һ�3ơ��r�q_�$PIP��N&`H�l�@���#@CORDED�d�p >f�fpO�� �< D ��OB⁴sd���Kӕи��qSYS�A�DR��f��TCH�t� = ,8`E�No��1Ak�_{��-$Cq,Be�VWVA~��> �  �&��PREV_R�T�$EDIT�r&VSHWRkqP�֑ &R:�v�D���JA�$�a$HECAD�6�� �z#�KE:�E�CPSP]D�&JMP�L~�2�0R*P��?��1�%&I��S�rC�pN�E; �q�wTICKğC��M�13�3HN��@ @� 1Gu��!_GPp6��0S3TY'"xLO��:��2l2?�A t 
�m G3%%$R!{�=:��S�`!$��w`����ճ���Pˠp6S�QU��E��u�TEsRC�0��TSUtB ����hw&`gw�Q)�pO����@�IZ��{��^�P�R�kюB1XPU����E_DO��, XuS�K~�AXI�@���UR�pGS�r � ^0�&��p_) ��ET�BPm��o���0Fo��0A|����Rԍ��a;�S=R�Cl>@P� �b_�yUr��Y��yU�� yS��yS���UЇ�U�� �U���U�]��Ul[��Y�bXk�]Cm������YRSC�� 7D h�DS~0��fQ�SP���eATހ��A]0,2N�AD�DRES<B} S�HIF{s��_2C�H���I��=q�+TVsrI��E"����a�Ce�
��
;�V8W�A��F \��qA��0l|\A@�rC��_B"R{zp�ҩq�T�XSCREE�Gzv��1TINA����t{����A�b?�H T1�ЂB��р��I��A��BE�y RRO������� B���v1UE4I �g��!p�S��RSM<]0�GUNEX(@~���j�S_S�ӆ��Á։񇣣�ACY�0�o 2H�pUE;��J�����@GMTJ��Lֱ�A��O	�/BBL_| W8��ЧK ��0s�OM���LE/r��� TO�!�s�RIGH��B�RD
�%qCKGR8л�TEX�@����WIDTH�� �Bh[�|�<��I_��}Hi� L 8K�B��_�!=r���R:�@_��Yґ��O6qJ�Mg0紐U��rh�Rm��LUMh��FpERVw �QP���`�N��&�/GEUR��FP)�M)� LP��(RE%@�a)ק�a�!��f ��5�6�7�8 Ǣ#B�É@���tP�f�W�S@M�U{SR&�O <�����U�Qs�FOC\)��PRI;Qm� �:���TRIP�Om�UN����Pv��0��f%��'���@��0 Q����AG �0T� �a>q�OS�%�RPo���8�R/�A�H�L4$����U¡�SU�g�p�¢5��OFF���T�}�O�� G1R�����S�GUN��6�B�_SUB?���,�SRTN�`TUg2���mCOR| D�RAU�rPE�TZ�#'�VC�C��	3V AC?36MFB1f$c�{PG �W (#�.�ASTEM����L�0PE��T3G��X �\ ��MOV1Ez�<���AN�� ����M���LIM_X��2��2��7�,������ı�
��VF@�`EӐ�~��04Y�F�IB�7���5S���_Rp� 2��� WİGp+@��}���P��3�Zx ���3���A�rݠCZ�DRID�����Vy08�90� D~e�MY_UBYd�@��6��@��!��X��P_S��3��mL�KBM,�$+07DEY(#EX`������UM_MU� X����ȀUS�� �z��G0`PACI�� �а@��:��:,�:����RE/�3qL�+���:[��TA�RG��P�r��R<�\ d`��A���$�	��AR��SWH2 ��-��@Oz��%qA7p�yREU�Uh�01�,�HK�2]g0�qP� N�� �EAM0GWORx���MRCV3�W^ ���O�0M��C�s	���|�REF_���x(�+T � ���������3_RCH4(a �P�І�hrj�NA�5��0�_ ��2����L@4��n�@@OU~7w�6���Z��a2[ư�RE�p�@;0\��c�a'2K�@SUL���]��C��0�^��� NT��L�3��@(6I�(6q�(3� L��@Q5��Q5I�]7q�}�)Tg`4D`�0.`0ПAP_HUC�5S]A��CMPz�F�6(�5�5�0_�aR��a��1I\!X�9|"GF}S��ad ��qM��0p�UF_x�0�B� �ʼ,RO��Q���'����UR�3GR�`.�3IDp���)�D�;��A��~�IEN��H{D���V@A J���S͓UWm�i=�����TYLO�*�5����b�t +�cPA�= �cCACH�vR��UvQ��Y��p�#CZF�I0sFR�XT����Vn+$HO��� �P!A3�XBf�(1 ���$�`VPy� ^bO_SZ313he6K3he12J�eh chG�6chWA�UMP�j���IMG9uPAD<�iiIMRE�$�b/_SIZ�$P�����0 ��ASYNBU=F��VRTD)u5t�qΓOLE_2DPJ�Qu5R��C��U���vPQuECCUlVEMV �U�r�W�VIRC�aIuVTPG���rv1s��5qFMPLAqa��v�V�0�cm� CKL�AS�	�Q�"��dC  �ѧ%ӑӠ@}���$�Q���Ue | �0!�rSr�T�#0! �r�iI��m�v6K�BG��VE�Z��PK= �v�Q�&�_�HO�0��f � �>֦3�@Sp�SL�OW>�RO��A�CCE���!� 9�V�R�#���p:���AD�����PAV�j�� uD����M_B"����^�JMPG ��g|:�#E$SSC�� x&�vPq��hݲvQ�S�`qVN��LEXc�i T`�sӂ��Q�FLD �DEsFI�3�02����:��VP2�VjO� �A��V�4>[`MV_PIs���t���A�@��FI��|�Z��Ȥ�����A0���A��~�GAߥ1 �LOO��1 JCB����Xc��^`�#PLCANE��R��1F�c �����pr�M� [`�噴��S����f�����Af��R�Aw�״t�U��pRKE��d�V�ANC�A���� �k���ϲϡ�R;_AA� l��2�� ��p�#Hć�m h�@��O K�$������kЍ0OU&A�"A��
p�pSK�TM�@FVIEM 2l ���P=���n <�<��dK�UMMYRK1P��`D倛�ACU��#AUކ�o $��TI}T�$PR�����OP���VS�HIF�r�p�`J�Qsԙ�fOxE-$� _R�`U�#�� ��s��q������G�"G�޵'�T�$�SsCO{D7�CNTQ  i�l�>a�-�a�;�a�H�a�V���1�+�2�u1��D���� � � SMO�Uq���a�JQ������a_�R[�r�n��*@LIQ�AA/`�XKVR��s�n�TL�ޡ�ZABC�tВt�c�
AZIeP��u���LVbc�Ln"�H�ZMPkCFx�v:�$��� ���DMY_L�N�������@y�w �Ђ(a�u� MCM��@CbcCART_��DPN� $J71D��=N�Gg0Sg0�BUXW|� ��UXEUL|ByX���	������x P	���m�YH�Db  y 80���0�EIGH�3n�?(�� H����$z a���|�����$B� �Kd'��_��L3�R�VS�F`���OVC�2'�$|�>P&���
q���5D�T�R�@ �VD��SP9HX��!{ ,� �*<�$R�B2 �2 ���C!��  �H�V+@b*c%g!)`+g"�`V*�,?8�?�V+�/ V.�/�/?�/�/V(7%3@/R/d/v/�/6?�/ �/�?�?�?O4OOION;4]?o?�?�?�?SO �?�?�O_�O0_Q_8_f_N;5zO�O�O�O�O p_�O_o8o�_MonoUo�oN;6�_�_�_�_ �_�oo%o4Uj�r�N;7�o�o�o �o�o� BQ�r�5� ��������N;8�� ���Ǐ=�_�n����R���ş��ڟN;G ;� џ�
������W�i� {�������ï�.��@�����A��dW� <�N�|�������Ŀֿ �ޯ���0�B�_� R�d�꿤϶������� ������*�L�^�� rτ�
������������&�8�J�l�~�; `ҟ @�з�@���ߩ��-��� �&�,���9�{��� ��a������������� ��A'Y�� �������a#1�
��N;�_MODE  ���S ��[�Y�B���
/\/�*	|/�/R4CWO�RK_AD�
 {9dT1R  ����� �/� _INOTVAL�+$���R_OPTION�6 �q@V_�DATA_GRPg 27���D��P�/~?�/�?�9��? �?�?�?OO;O)OKO MO_O�O�O�O�O�O�O _�O_7_%_[_I__ m_�_�_�_�_�_�_�_ !ooEo3oioWoyo�o �o�o�o�o�o�o /eS�w�� �����+��O� =�s�a�������͏�� �ߏ��9�'�I�o��]�����$SAF�_DO_PULS�� �~������CAN_TIM�����ΑR +��+Ƙ��5�;#U!P"�1!��� �?E�W�i�{� ����.�ïկ������'(~�T"2�F���dR�I�Y��2�o+@a얿�����)�u��� k0ϴ��_ ��  T�� � �2�D�)�T D��Q�zόϞ� ����������
��.� @�R�d�v߈ߚ�/V�������������R�;�o� �W�p��
�t��Diz$� �?0 � �T"1! ��������� ��������*�<�N� `�r������������� ��&8J\n ��������@"4FX ��� �������� /`4�=/O/a/s/�/ �/�/�/�/�/�!!/ �0޲k�ݵu�0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ ok$o 6oHoZolo~o�o�o�o �o1/�o�o 2D Vhz�/5?��� �����&�8�J� \�n���������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ���`Ò�ϯ� ���)�;�M�_�q� ��������˿ݿ� �����3� ����&2,��	12�345678v��h!B!��*2�Ch���0�� �����������!�3� 9ѻ�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�h�K߰����� ����
��.�@�R�d� v�������������� *<N`r� ������ &��J\n��� �����/"/4/ F/X/j/|/;�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�/ �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_�?L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o=_�o�o �o�o�o�o 2D Vhz�����h������u�o.��@�R���Cz  �B��   ����2&� � �_�
���  	�_�2�Տ�����_�p������ ďi�{�������ß՟ �����/�A�S�e� w���������N���� ��+�=�O�a�s��� ������Ϳ߿���'�9�K�_�������<v�_��$SCR�_GRP 1
�+� +�� t� ��� ���	 ���������� ������_������)��a����&�DE� DW8���l�&��G�CR-35�iA 901234567890��_M-20��8��?CR35 ��:�#
��������������:֦�Ӧ�G�D��&������	���]�o����:����H���>�� ���������&���ݯ:��j����g��,����B�t�����������A����  @��`��@� ( ?�=��Ht�P
���F@ F�` z�y������  �$H��G`s^p��B�� 7��/�0//-/ f/Q/�/u/�/�/�/8�@��P�� 7%?�����"?W?-2?<����]? H�1�?t���7�������?�-4A, �&E@�<�$@G�B-1 3OZOlO-:HA�H�O�O|O P�B(�B�O�O�_��EL_DEFAULT  ����`~SHOTSTR#]�JA7RMIPOWE?RFL  i�/U�YTWFDO$V� /URRVENT? 1����NU� L!DUM�_EIP_-8�j�!AF_INEx#P�_-4!FT�_�->�_;o!��`o ��*o�o!RP?C_MAIN�ojhq�vo�o�cVIS�o�ii��o!TP&pPU�Ydk�!
PMON_POROXYl�VeZ��2r��]f��!�RDM_SRV���Yg�O�!R���k��Xh>���!
��`M��\i���!RLSYNC��-98֏3�!R3OS�_-<�4"���!
CE4pMTC�OM���Vkn�˟!=	��CONS̟�W�l���!��WA'SRC��Vm�c�;!��USBd��XnR���Noӯ����� ��!��E��i�0����WRVICE_K�L ?%�[ (�%SVCPRG1��-:Ƶ2ܿ�˰3�	�˰4,�1�˰5T�Y�˰6|ρ�˰�7�ϩ�˰�����9����ȴf�!�˱ο I�˱��q�˱ϙ�˱ F���˱n���˱��� ˱��9�˱��a�˱� ���7߱��_���� �����)����Q� ���y��'���O� ���w������ ���˰��İd� c������ =(as^��� ���/�/9/$/ ]/H/�/l/�/�/�/�/ �/�/�/#??G?2?k? V?}?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O�O�O�O	_�O�-_��_DEV ��Y�MC:�5Xd�GTGR�P 2SVK ��b�x 	� 
 ,�P5_�_�R�_�_ �_�_�_�_3ooWo>o {o�oto�o�o�o�o�o �o/A�_e� ��������  �=�$�6�s�Z���~� ��͏���H�'�ޏ K�2�o���h�����ɟ ۟���#�5��Y� @�}�d�v���
�ׯ� Я���1��*�g�N� ��r��������̿	� ��?�&�c�u�̯�� PϽ��϶������)� �M�4�q�X�jߧߎ� �߲������%�|�� [���f������ �������3��W�i� P���t���������>� A(eL^ �������  =O6sZ��  ���/�'// K/]/D/�/h/�/�/�/ �/�/�/�/#?5??Y? �N?�?F?�?�?�?�? �?O�?1OCO*OgONO �O�O�O�O�O�O�O�O,_kT �"V		_R_�=_v_a_�_�_�_�[%���_�_�S��� a�Qeo)goIo7o mo[o�o�i�_�oi�o �o�o%'9o �o��o_���� ��!�w�n��G� ����ŏ���׏�O� 4�s���g���w����� �����'��K�՟?� -�c�Q�s��������� �#�����;�)�_� M�o���ׯ������� ݿ��7�%�[ϝ��� ��K�m�Gϵ������ ��3�u�Zߙ�#ߍ�{� �ߟ߱������M�2� q���e�S��w��� ����%�
�I���=�+� a�O���s�������� !���9']K ������q�m� �5#Y��� I�����/� 1/sX/�!/�/y/�/ �/�/�/�/	?K/0?o/ �/c?Q?�?u?�?�?�? ?�?O�?�?�?)O_O MO�OqO�O�?�OO�O _�O__%_[_I__ �O�_�Oo_�_�_�_�_ oo!oWo�_~o�_Go �o�o�o�o�o�o	_o �oV�o/�w�� ���7�[�O� �_���s�����͏� �3���'��K�9�[� ��o����̟����� �#��G�5�W�}��� ���m�ׯů���� �C���j�|�3�U�/� ��ӿ������]�B� ���u�cυχϙ��� ����5��Y���M�;� q�_߁߃ߕ������ 1߻�%��I�7�m�[� }�������	������ !��E�3�i������ Y���U������� A��h��1��� ����[@ 	sa����� �3/W�K/9/o/ ]/�/�/�/��/�/�/ �/�/?G?5?k?Y?�? �/�?�/?�?�?�?�? OCO1OgO�?�O�?WO �O�O�O�O�O�O	_?_ �Of_�O/_�_�_�_�_ �_�_�_G_m_>o}_o qo_o�o�o�o�o�oo Co�o7�oGm[ ���o��� �3�!�C�i�W���� ���}��Տ���/� �?�e�����ˏU��� ���џ���+�m�R� d��=��������߯ ͯ�E�*�i��]�K� m�o�������ۿ�� A�˿5�#�Y�G�i�k� }ϳ�����ϣ���� 1��U�C�e߻��ϲ� �ϋ�����	���-�� Q��x��A��=�� �������)�k�P��� ���q����������� C�(g���[I m���� ? �3!WE{i� �������// /S/A/w/��/�g/ �/�/�/�/�/+??O? �/v?�/??�?�?�?�? �?�?�?'Oi?NO�?O �OoO�O�O�O�O�O/O UO&_eO�OY_G_}_k_ �_�_�__�_+_�_o �_/oUoCoyogo�o�_ �oo�o�o�o	+ Q?u�o��oe� �����'�M�� t��=�����ˏ��� ݏ�U�:�L��%��� m�����ǟ���-�� Q�۟E�3�U�W�i��� ��ï��)����� A�/�Q�S�e���ݯ¿ ��������=�+� Mϣ�ɿ��ٿs��ϻ� ������9�{�`ߟ� )ߓ�%ߣ��߷����� �S�8�w��k�Y�� }�������+��O� ��C�1�g�U���y��� �����'���	? -cQ�����w �s�;)_ ���O���� �//7/y^/�'/ �//�/�/�/�/�/? Q/6?u/�/i?W?�?{? �?�?�??=?OM?�? AO/OeOSO�OwO�O�? �OO�O_�O_=_+_ a_O_�_�O�_�Ou_�_ �_o�_o9o'o]o�_ �o�_Mo�o�o�o�o�o �o5wo\�o%� }�����="� 4����U���y��� ��ӏ���9�Ï-�� =�?�Q���u����ҟ �����)��9�;� M���ş���s�ݯ˯ ��%��5������� ��[�����ٿǿ��� !�c�Hχ��{�ϋ� �ϟ�������;� �_� ��S�A�w�e߇߭ߛ� �����7���+��O� =�s�a�������� �����'��K�9�o� �����_���[����� ��#G��n��7 ������� aF�yg�� ����9/]� Q/?/u/c/�/�/�/� %/�/5/�/)??M?;? q?_?�?�/�?�/�?�? �?�?%OOIO7OmO�? �O�?]O�O�O�O�O�O !__E_�Ol_�O5_�_ �_�_�_�_�_�_o__ Do�_owoeo�o�o�o �o�o%o
�o�o�o =sa����o��!+q�$SERV�_MAIL  �+u!���OUTwPUT�$�}@�RV 2�v;  $� (�q�<}��SAVE7�	��TOP10 2>W� d 'ݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w�������0��ѿ�u��YP����FZN_CFG ;�u$�~�����GRP 2��D� ,B �  A[�+qD;�� B\��  B�4~�RB21ފ�HELL��u��j�k�2�����%RSR������ �
�C�.�g�Rߋ�v� ���߬�����	���-��?�Q��  �_�%Q���_����,p�������g�2,pd�����HK 1�� ��E�@�R�d����� �������������*<e`r���OMM ������FTOV_ENB��_���HOW_R�EG_UI�	�IMIOFWDL� ��^�)WAIT����$V1��^�NTIM����VA�_)_�UNIT����L]CTRYB���MB_HDD�N 2W�  2�:%0 �pQ/�qL/ ^/�/�/�/�/�/�/�/��"!ON_ALI_AS ?e�	f�he�A?S?e?w?�: /?�?�?�?�?�?OO &O8OJO�?nO�O�O�O �OaO�O�O�O_"_�O F_X_j_|_'_�_�_�_ �_�_�_oo0oBoTo �_xo�o�o�o�oko�o �o,�oPbt �1������ �(�:�L�^�	����� ����ʏu�� ��$� Ϗ5�Z�l�~���;��� Ɵ؟����� �2�D� V�h��������¯ԯ ���
��.�ٯR�d� v�����E���п��� ϱ�*�<�N�`�r�� �ϨϺ���w����� &�8���\�n߀ߒߤ� O�����������4� F�X�j�|�'����� �������0�B��� f�x�������Y����� ����>Pbt ������ (:L�p�� ��c�� //$/ �H/Z/l/~/)/�/�/ �/�/�/�/? ?2?D?�V?]3�$SMON�_DEFPRO ����1� *S�YSTEM*0�m6RECALL �?}9 ( ��}5xcopy �fra:\*.*� virt:\t�mpback�1=�>147.87.�149.40:15172 �1�>	O�O+L}J�2mdb�:schinde�l_5sem.t=p�5emp\HM�?�O�O�O }9�4s�:orderfil.dat�<tO�?�O_*_}0?F�?�O@�1�O_�_�_8C4�5��?�?�6t_�_o)o  �?�_�_�?o�o�o;O MO_OqO�o&�O�O T_�O��7_I_d m_�"��_HoZo�_ �����3oEoV�io{� ���o�o�o�o���� ��/ASv������ ��ڟ�������� =�Џ]�s����(����̯ޯ������9�
�xyzrate 11 J�\�n����4#�6���61߿� I��ϔϦ�9�K�]� o����$߷�ɟR�� �ϐߢ�5�G�b�k�}� � ﳯůؿ��ߌ� ��1�C�T�g�y�
�� ����������+���-� ?�Q�t����*�� ��������;��� [q�&���� ��������R�� /"/5G�k� �/�/��X�{/? ?1C�/g�/�?�? ���a?w?�?O-/ ?/�?c/�?O�O�O�/ P?]O�/�O_(_;?�O@�Oq?_�_�_��6ȿ�Z_l_~_o!o4�F�:1289]��_o�o��o7�tpdisc 0Io[a]ooo�o�$7�tpconn 0 �o�o�o��o���v�$SN�PX_ASG 2�����q�� P 0 �'%R[1�]@1.1��y?��s%�!��E�(� :�{�^�������Տ�� ʏ���A�$�e�H� Z���~���џ����؟ �+��5�a�D���h� z�����ů�ԯ��� 
�K�.�U���d����� ��ۿ������5�� *�k�N�uϡτ��Ϩ� �������1��U�8� Jߋ�nߕ��ߤ����� �����%�Q�4�u�X� j����������� ��;��E�q�T���x� ����������% [>e�t�� ����!E( :{^����� �/�/A/$/e/H/ Z/�/~/�/�/�/�/�/ �/+??5?a?D?�?h? z?�?�?�?�?�?O�? 
OKO.OUO�OdO�O�O �O�O�O�O_�O5__ *_k_N_u_�_�_�_�_ �_�_�_o1ooUo8o�Jo�ono�o�o�d�tPARAM �u��q �	���jP�d9p�h�t��pOFT_K�B_CFG  ��c�u�sOPIN_�SIM  �{�vn��p�pRV�QSTP_DSB�W~r"t�HtSR� Zy � �& SCHIN�DEL_5SEM��u�vTOP_�ON_ERR  �&�Dx8�PTN �Zuk��A4�RING_P�R�D��`VCNT_GP 2Zu:q�!px 	r���ɍ���׏��wVD>��RP 1�i p�y��K�]�o��� ������ɟ۟���� #�5�G�Y���}����� ��ůׯ�����F� C�U�g�y��������� ӿ��	��-�?�Q� c�uχϙϫ������� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�^�[�m��� �����������$�!� 3�E�W�i�{������� ��������/A Sew����� ��+=Ov s������� //</9/K/]/o/�/ �/�/�/�/�/?�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO)��PRG_COUN�T8v�k�GuKBENB��FEMpC:t}O_UPD 1�{T  
4Or�O �O�O__!_3_\_W_ i_{_�_�_�_�_�_�_ �_o4o/oAoSo|owo �o�o�o�o�o�o +TOas�� ������,�'� 9�K�t�o��������� ɏۏ����#�L�G� Y�k���������ܟן ���$��1�C�l�g� y���������ӯ���� 	��D�?�Q�c����� ����ԿϿ�����)�;�d�_�q�=L_I�NFO 1�E��@ �2@����������� �����_B+���!w'��2��mn�£n<LYSDEBUGU@ʶ@���d�If�SP�_PASSUEB�?x�LOG  *���C��*ؑ��  ��A��U�D1:\�ԘΥ�_MPC�ݵE&�8�A���V� �A�SAV !������ҶX���SVZ�T�EM_TIME �1"���@ 0*�Ќ��UX�X�����$T1SVGU�NS�@VE'�E���ASK_OPT�IONU@�E�A�A�+�_DI��qOG�B�C2_GRP 2�#�I�����@� � C���<Ko�CF�G %z��� ������`��	�. >dO�s�� �����*N 9r]����� ��/�8/#/\/n/ ��Z+�/Z/�/�/H/�/ ?�/'??K?]�k?=� @0s?�?�?�?�?�?�? O�?OO)O_OMO�O qO�O�O�O�O�O_�O %__I_7_m_[_}__ �_�_�X� �_�_oo /o�_SoAoco�owo�o �o�o�o�o�o= +MOa���� �����9�'�]� K���o���������ɏ ���#��_;�M�k�}� �������ß�ן� �1���U�C�y�g��� ������������	� ?�-�c�Q�s������� ���Ͽ����)� _�Mσ�9��ϭ����� ��m���#�I�7�m� ߑ�_ߵߣ������� ����!�W�E�{�i� ������������� �A�/�e�S�u�w��� ����������+= O��sa���� ���9'] Kmo����� ��#//3/Y/G/}/ k/�/�/�/�/�/�/�/ ??C?��[?m?�?�? �?-?�?�?�?	O�?-O ?OQOOuOcO�O�O�O �O�O�O�O__;_)_ __M_�_q_�_�_�_�_ �_o�_%oo5o7oIo omo�oY?�o�o�o�o �o3!CiW� ������� �-�/�A�w�e����� �����я���=� +�a�O���s������� ߟ͟��o�-�K�]� o�ퟓ�����ɯ����צ��$TBCS�G_GRP 2&�ץ� � �� 
 ?�  6�H�2�l�V� ��z���ƿ��������(�d��E+�?�	 HC{���>���G�����C�  A�.�e�q�C��>ǳ33��S�/]϶�Y���=Ȑ� C\  �Bȹ��B���>�����P���B�Y�z��L�H�0�$����J�\�n�����@�Ҿ��������߀=�Z�%�7����?�3�����	V�3.00.�	cwr35��	*�����
�������� �3��4�   {�CT�v�}��J2�)�������CFG +ץe'� *������qI���� .<
�<bM�q �������( L7p[�� ����/�6/!/ Z/E/W/�/{/�/�/�/ �/.�H��/??�/L? 7?\?�?m?�?�?�?�? �? OO$O�?HO3OlO WO|O�O����Oӯ�O �O�O!__E_3_i_W_ �_{_�_�_�_�_�_o �_/oo?oAoSo�owo �o�o�o�o�o�o+ O=s�E��� Y�����9�'� ]�K�m�������u�Ǐ ɏۏ���5�G�Y�k� %���}�����ßşן ���1��U�C�y�g� ������ӯ������ 	�+�-�?�u�c����� �����Ͽ���/� A�S�����qϓϕϧ� �������%�7�I�[� ��mߣߑ߳����� �߷��3�!�W�E�{� i����������� ��A�/�e�S�u��� ������������ +aO�s�� e�����'K 9o]���� ���#//G/5/k/ }/�/�/[/�/�/�/�/ �/??C?1?g?U?�? y?�?�?�?�?�?	O�? -OOQO?OaO�OuO�O �O�O�O�O�O___ M_�e_w_�_3_�_�_ �_�_�_oo7o%o[o moo�oOo�o�o�o�o �o!3�o�oiW �{������ �/��S�A�w�e��� ����я������� =�+�M�s�a������� ��ߟ�_	���_ן ]�K���o�������ۯ ɯ���#���Y�G� }�k�����ſ׿���� ����U�C�y�g� �ϋ��ϯ�������� 	�?�-�c�Q�s�u߇� �߫��������)�� 9�_�M����/���� i������%��I�7� m�[������������� ������EWi{ 5������� �A/eS�w �����/�+/ /O/=/_/a/s/�/�/ �/�/�/�/?'?��?? Q?c??�?�?�?�?�? �?�?O�?5OGOYOkO�)O�O}O�O�O�O�N s �@S V�_R�$TBJO�P_GRP 2,��E� / ?�V	-R4S�.;\��@|�u0{SPU >���UT @��@LR	 �C�� �Vf  C����ULQLQ>�33��U�R����U�Y?~�@=�ZC��P׌�ͥR��P � B��W$o/gC���@g�dDb�^���eeao�P�&ff�e=�7L3C/kaB o�o�P��P�efb-C�p��^g`�d�o��PL�Pt<�eVoC\  �Q@�'p}�`�  A�o�L`�_wC�BrD�S�^�]�_�S~�`<PB��P0�anaa`C�;�`L�w�aQoxp��x�p:��XB$4'tMP@�PCHS��n���=�P����trd<M�gE�2pb ����X�	��1�� )�W���c�������� ����󟭟7�Q�;�PI�w���;d�Vɡ��U	V3.00�RScr35QT�*�QT�A�� �E�'E�i��FV#F"w�qF>��FZ�� Fv�RF�~�MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
�D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt���ٵ=�_t��V �R�p�V9� ]ESTP�ARtp�HFP*SH�R\�ABLE 1%/;[%�SG��Q �W�G�G�GȨ WQG�	G�
G��GȖ�QG�G�8G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ߱���w�S]�CS !ڄ�� �����������&� 8�J�\�n��������� ���� ]\�`��	� �(�:�����
��.��@�w�NUM  ��EEQ�P�	P ۰ܰw�_CFG 0��)r-P�IMEBF_TT�b��CSo�,VER�ڳ-B,R 1=1;[ 8��R��@� �@&   �������/ /)/;/M/_/q/�/�/ �/�/�/?�/?J?%? 7?M?[?m?>�@�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_l_�Y�@cY�MI_CWHAN8 c c�DBGLV��:�cX�	`ETHER_AD ?f�\`��?�_uo�oQ��	`ROUTV!�	
!�d�o�lSN�MASKQhcba255.uߣ'�9ߣY�OOLOF/S_DIb��U;i�ORQCTRL �2		�Ϸ~T �����#�5�G� Y�k�}�������ŏ׏ �����.��R�V��PE_DETAI�/h|zPGL_CONFIG 8�	����/cel�l/$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c� u�����(���ϯ�� ����;�M�_�q��� ��$�6�˿ݿ��� %ϴ�I�[�m�ϑϣ� 2����������!߰� ��W�i�{ߍߟ߱�%}F�������/�A��C�i�H�Eߞ�� ��������?��.�@� R�d�v���������� ������*<N` r������ �&8J\n� �!�����/ �4/F/X/j/|/�// �/�/�/�/�/??�/ B?T?f?x?�?�?+?�? �?�?�?OO�?>OPO�bOtO�O�O�O����User Vi�ew ��}}12�34567890 �O�O�O_#_5_=T�P,��]_���I2�I:O �_�_�_�_�_�_X_j_�B3�_GoYoko}o�o�o o�op^46o�o�1CU�ovp^5 �o�����	�h*�p^6�c�u����� �����ޏp^7R�� )�;�M�_�q�Џ��p^8�˟ݟ���%����F�L� lCamera�J ��������ӯ���E~��!�3��OM�_�`q��������y  e� �Yz���	��-�?�Q� ��uχϙ�俽���������>��e�5i�� c�u߇ߙ߽߫�d��� ���P�)�;�M�_�q� ��*�<��i������� ��)���M�_�q��� ��������������<� û��=Oas�� >����*' 9K]f�Q��� ����/�%/7/ I/�m//�/�/�/�/ n<��^/?%?7?I? [?m?/�?�?�? ?�? �?�?O!O3O�/<׹� �?O�O�O�O�O�O�? �O_!_lOE_W_i_{_�_�_FOXG9+_�_�_ oo(o:o�OKopo�o )_�o�o�o�o�o 
��	g�0�oM_q ���No����o �%�7�I�[�m�& l�n��Ə؏����  ��D�V�h������� ��ԟ柍�g�ڻ}� 2�D�V�h�z���3��� ¯ԯ���
��.�@� R���3uF�鯞���¿ Կ������.�@ϋ� d�vψϚϬϾ�e�w� ��U�
��.�@�R�d� ψߚ߬��������� ��*���w���v� �������w���� �c�<�N�`�r����� =�w��-����� *<��`r�����������  ��1CUgy��������   -/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E_W_i_�  
���(  �%( 	 y_�_�_�_ �_�_�_o	o+o-o?o@uoco�o�o�o�Z* �Q&� J\n������o ���9�(�:�L� ^�p���������܏ � ��$�6�}�Z�l� ~�ŏ����Ɵ؟��� C�U�2�D�V���z��� ����¯ԯ���
�� c�@�R�d�v������ ��п�)���*�<� N�`ϧ����ϨϺ�� ������&�8��\� n߀��Ϥ߶������� ��E�"�4�F��j�|� ����������� �e�B�T�f�x����� ��������+�, >Pb������� ���(o� ^p������ � /G$/6/H/�l/ ~/�/�/�/�//�/�/ ?U/2?D?V?h?z?�?�/�`@ �2�?�?��?�3�7�P��!�frh:\tpg�l\robots�\m20ia\c�r35ia.xml�?;OMO_OqO�O�O�O�O�O�O�O �� �O_(_:_L_^_p_�_ �_�_�_�_�_�O�_o $o6oHoZolo~o�o�o �o�o�o�_�o 2 DVhz���� ��o�
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟�ݟ� �&�8�J�\�n����� ����ȯߟٯ���"� 4�F�X�j�|��������Ŀ־�8.1 ��?@88�?�ֻ�ֿ�3�5�G� iϓ�}ϟ��ϳ����� ���5��A�k�U�w���߿��$TPGL�_OUTPUT �;�!�! ��������,� >�P�b�t����� ��������(�:�L�@^�p�������������2345678901�������� �"��BTfx� �4�����
}$L^p�� ,>��� //$/ �2/Z/l/~/�/�/:/ �/�/�/�/? ?�/�/ V?h?z?�?�?�?H?�? �?�?
OO.O�?<OdO vO�O�O�ODOVO�O�O __*_<_�OJ_r_�_ �_�_�_R_�_�_oo &o8o�_�_no�o�o�o �o�o`o�o�o"4 F�oT|����\��}�����0�B�T�e�@������� ( 	 �� Џ������<�*� L�N�`���������ޟ ̟���8�&�\�J� ��n���������ȯ���"�������*�X� j�F�����|�¿Կ�� C���ϱ�3�E�#�i� {�忇ϱ�S������� ���/ߙ�S�e�߉� ��y߿���;����� ��=�O�-�s���ߩ� ��]��������'��� �]�o���������� ��E�����5G% W}������g� ��1�Ug	 w�{��=O	/ /�?/Q///u/�/� �/�/_/�/�/�/�/)? ;?�/_?q??�?�?�? �?�?G?�?O�?OIO [O9OO�O�?�O�OiO �O�O�O!_3_�O_i_ {__�_�_�_�_�_�R��$TPOFF_�LIM >�op:���mqbN_�SV`  l��jP_MON M<6�dopop�2l�aSTRTC�HK =6�f�� bVTCOMP�AT-h�afVWV_AR >Mm�h.1d �o �oop�`ba_DEFPROG %|j�%SCHIND?EL_5SE`N�if_DISPLA�Y`|n"rINST�_MSK  t|� ^zINUSE9R�odtLCK�|}{�QUICKMEN��dtSCRE�p�6��btps�cdt�q��b*�_�.�ST�jiRAC�E_CFG ?�Mi�d`	�d
�?�u�HNL 2E@|i����k r ͏ߏ���'�9�K�l]�w�ITKp2A��� �%$1234567890����  =<��П��  !���p��=��c��^��� �������.���R�� v�"�H�ί��Я��� ���*�ֿ���r�2� ������4�޿�ϰ��� &���J�\�n���@ߤ� d�v��ς������4� ��X��*��@��� ���ߨ�������T� ��x������l��� �����,�>�P����� ��FX��d����� �:�p"� �o�����F 6HZt~��N/ t/�/��// /2/�/ V/?(?:?�/F?�/�/ �/j?�??�?�?R?�? v?�?QO�?lO�?�O�O O�O*O|O_`O _�O 0_V_h_�Ot_�O__ �_8_�_
oo�_@o�_ �_�_Lodo�_�o�o4o �oXojo3�oN�or���o��s�S��B���z�  h��z ��C�:y
 P�v�]�����UD1:\������qR_GRP �1C��� 	 @Cp���$� �H�6�l�Z��|������f���˟���ڕ?�  
���<�*� `�N���r�������ޯ ̯��&��J�8�Z����	�u�����sS�CB 2D� �����(�:�L��^�pς��|V_CONFIG E����@����ϖ�OUT?PUT F�������6�H�Z� l�~ߐߢߴ������� �����#�6�H�Z�l� ~������������ ��2�D�V�h�z��� ������������
� .@Rdv��� ����)< N`r����� ��//%8/J/\/ n/�/�/�/�/�/�/�/ �/?!/4?F?X?j?|? �?�?�?�?�?�?�?O O/?BOTOfOxO�O�O �O�O�O�O�O__+O >_P_b_t_�_�_�_�_ �_�_�_oo'_:oLo ^opo�o�o�o�o�o�o �o $����!�b t������� ��(�:�-o^�p��� ������ʏ܏� �� $�6�G�Z�l�~����� ��Ɵ؟���� �2� D�U�h�z�������¯ ԯ���
��.�@�Q� d�v���������п� ����*�<�M�`�r� �ϖϨϺ�������� �&�8�J�[�n߀ߒ� �߶����������"� 4�F�W�j�|���� ����������0�B� S�f�x����������� ����,>Pa� t��������(:L/x���k}gV� K���//&/8/ J/\/n/�/�/�/W�/ �/�/�/?"?4?F?X? j?|?�?�?�?�/�?�? �?OO0OBOTOfOxO �O�O�O�?�O�O�O_ _,_>_P_b_t_�_�_ �_�O�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����o� ��� �2�D�V�h� z��������ԏ��� 
��.�@�R�d�v��� ������Ϗ����� *�<�N�`�r������� ��˟ޯ���&�8� J�\�n���������Ż��$TX_SCR�EEN 1G�g�}�ipnl/��gen.htmſ�*��<�N�`ϽPa�nel setupd�}�dϥϷ����������ω�6�H� Z�l�~ߐ�ߴ�+��� ����� �2�߻�h� z������9�g�]� 
��.�@�R�d���� �����������}� ��<N`r�� ;1��&8 �\��������QȾUALRM_MSG ?��� �Ȫ-/?/ p/c/�/�/�/�/�/�/��/??6?)?Z?%S�EV  -��6"ECFG �I��  �ȥ@�  A�1 �  B�Ȥ
  [?ϣ��?OO%O7O IO[OmOO�O�O�G�1�GRP 2J�;; 0Ȧ	 �?�O� I_BBL_N�OTE K�:T��lϢ��ѡ�0RDEF�PRO %+ (%N?u_Ѡc_�_�_ �_�_�_�_o�_o>o�)oboMo�o\INU?SER  R]�O��oI_MENHI�ST 1L�9  �( _P���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1�oCUgy�)
13/��� ��p|o"�4�F�X�j� |������ď֏��� ���0�B�T�f�x�� �����ҟ������ ,�>�P�b�t������ ��ί����9Rq ��B�T�f�x������� ��ҿ����ϩ�>� P�b�tφϘ�'�9��� ������(߷�L�^� p߂ߔߦ�5�������  ��$����Z�l�~� ����C��������  �2��/�h�z����� ����������
. @��dv���� �_�*<N �r�����[ �//&/8/J/\/� �/�/�/�/�/�/i/�/ ?"?4?F?X?C�U��? �?�?�?�?�?�/OO 0OBOTOfO�?�O�O�O �O�O�O�O�O_,_>_ P_b_t__�_�_�_�_ �_�_�_o(o:oLo^o po�oo�o�o�o�o�o  �o$6HZl~ i?{?������ 2�D�V�h�z���� -�ԏ���
���� @�R�d�v�����)��� П���������N� `�r�������7�̯ޯ ���&���J�\�n�����������$U�I_PANEDA�TA 1N����ڱ  �	�}/fr�h/cgtp/w�idedev.stm���%�7�I�Y�)priρ�@�}�ϩϻ�������� )�)��M�4�q� ��jߧߎ�����������%�7��[�7���q}�ϕ��� ������B����%�I� [�m������
����� ������!E,i {b������l� ݰܳ7�<N `r����-�� �//&/8/�\/n/ U/�/y/�/�/�/�/�/ ?�/4?F?-?j?Q?�? �?%�?�?�?OO 0O�?TO�xO�O�O�O �O�O�OKO_�O,__ P_b_I_�_m_�_�_�_ �_�_oo�_:o�?�? po�o�o�o�o�oo�o  sO$6HZl~ �o�������  �2��V�=�z���s� ����ԏGoYo�.� @�R�d�v�ɏ���� П������<�N� 5�r�Y�������̯�� �ׯ�&��J�1�n� ������ȿڿ��� �c�4ϧ�X�j�|ώ� �ϲ���+�������� 0�B�)�f�Mߊߜ߃� �ߧ��������� P�b�t�������� ��S���(�:�L�^� ���i�����������  ��6ZlS`�w�'�9�}��@�"4FX)� }��l����� /j'//K/2/D/�/ h/�/�/�/�/�/�/�/�#?5??Y?��C�=���$UI_POST�YPE  C��� 	 �e?�?�2QUICK�MEN  �;��?�?�0RESTO�RE 1OC��  ��L?��6OCC1O��m aO�O�O�O�O�OuO�O __,_>_�Ob_t_�_ �_�_UO�_�_�_M_o (o:oLo^oo�o�o�o �o�o�oo $6 H�_Ugy�o�� ���� �2�D�V� h��������ԏ ����w�)�R�d�v� ����=���П���� ��*�<�N�`�r��� �����ޯ���&� ɯJ�\�n�������G��ȿڿ�����7SC�RE�0?�=�u1sc+@uU2K�3K�4K�5Kĕ6K�7K�8K��2U�SER-�2�D�ksTMì�3��4��5�ĕ6��7��8���0N�DO_CFG �P�;� ��0PDA�TE ����None�2��_INFO 1QC�@��10%�[��� Iߊ�m߮��ߣ����� �����>�P�3�t���i���<-�OFFS_ET T�=�� ��$@������1�^� U�g������������ ����$-ZQcu���?�
�����UFRAME  �����*�RTO?L_ABRT	(��!ENB*GR�P 1UI�1Cz  A��~��@~���������0UJ�9MSK  M@�;-N%8�%��/��2VCCM��V��ͣ#RG�#Y�9����/����D�BeH�p71C����3711?�C0�$MRf2_�*S��괰	���~XC56 *�?�6�Y��1$�5����A@3C��. 	��8�?��OO KOx1FOsO�5�51ⴰ_O�O�� B����A2�DWO �O7O_�O8_#_\_G_ �_k_}_�__�_�_�_��_"o�OFoXo�%TCC�#`mI1�i���u��� GFS�»2aZ; �| 2�345678901�o�b�����o@��!5a�4BwB�`�56 311:�o=L�Br5v1�1~1�2 ��}/��o�a��# �GYk}�p�� �����ُ�1�C� U�6�H���5�~���ߏ����	���4�dSEGLEC)M!v1b3��VIRTSYN�C�� ���%�SIONTMOU�������F��#b�U��U�(�u FR:\�H�\�A\�� ��� MC��L�OG��   U�D1��EX����'� B@ �����̡m��̡  �OBCL�1�H�� �  =	 �1- n6 � -������[�,xS�A�`=��͗���ˢ��TRA�IN⯞b�a1l�
�0d�$j�T2cZ; (aE2ϖ�i�� ;�)�_�M�g�qσϕ� ���������	��F�STAT dmB~2@�zߌ�*j$i�\���_GE�#eZ;7�`0�
� 0}2��HOMIN� �fU��U�� ~�����БC�g��X���JMPERR� 2gZ;
   ��*jl�V�7������ ��������
��2�@��q�d�v�B�_ߠREr� hWޠ$LEX�ԹiZ;�a1-e��V�MPHASE  �5��c&��!OF�F/�F�P2n�jJ�0�㜳E1�@��0ϒE1!1?s#33�����ak/�@kxk䜣!W�m[�䦲�[����o3;� [ i{���� /�O�?/M/_/q/ ��/��//�/'/9/ �/=?7?I?s?�/�?�/ �/�?�??Om?O%O 3OEO�?�?�O�?�O�O �?�O�O�O__gO\_ �OE_�O�_�O�O/_�_ �_�_oQ_Fou_�_|o �o�_�oo�o�o�o�o ;oMo?qof-�oI �����7� [P��������� ˏ��!�3�(�:�i��[�ŏg�}������TD_FILTEW��n�� �ֲ:���@���+�=�O�a� s���������֯� ����0�B�T�f�x����SHIFTME�NU 1o[�<��%��ֿ����ڿ� ���I� �2��V�h� ���Ϟϰ�������3��
�	LIVE/�SNAP'�vs�fliv��E�����ION * U<b�h�menu~߃������ߣ���p����	����E�.ォ50�s�P�@� �Z�AɠB8z�z�!�}��x�~�P��� ���MERb���<�0���kMO��q���z��WAITDINE�ND������O9K1�OUT���SD��TIM����o�G���#����C���b������RELEASE������TM�������_�ACT[�����_DATA r�%L����xRD�ISb�E�$X�VR�s���$Z�ABC_GRP �1t�Q�,#�r0�2���ZIP�u'�&����[�MPCF_G 1	v�Q�0�/� �w�ɤ� 	|�Z/  85�`�/�/H/�/l$?��+ �/�/�/?�/�/???|r?�?  �D0 �?�?�?�?�?�;����x�]hYLI�ND֑y� ���� ,(  * VOgM.�SO�OwO�O�M i?�O�O^PO1_ �OU_<_N_�_�O�_�_ �__�_�_x_-ooQo�8o�_�o�oY&#2z� ���oC� e?a?>N|�oq��햋qA�$DSPH�ERE 2{6M� �_�;o���!�io |W�i��_��,��Ï ���Ώ@��/�v��� e�؏��p�����������ZZ�� � N