��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ���!C�OUPLED�� $!PP_� C�ES0s!_81s!J�!PC> �! �� $SOFT��T_IDk2TO�TAL_EQs �$�0�0NO�2U SPI_INDE]��5Xk2SCREE�N_(4_2SIG�E0_?q;�0PK�_FI� 	$�THKYGPAN�E�4 � DUMMY1dDDd!OEU4LA R�!R��	 � $TI=T�!$I��N ��Dd�Dd �Dc@�D5��F6�F7�F8�F9�G0�G�GJA�E�GbA�E�G1�G1�G �F��G2�B!SBN_�CF>"
 8F CNV_J� ; �"�!�_CMNT�$�FLAGS]�C�HEC�8 � EL�LSETUP �� $HO30I�O�0� %�SMA�CRO�RREPR�X� D+�0��R{��T UTOBAC�KU�0 }�)DEVIC�CTI*0�� �0�#��`B�S$INT�ERVALO#IS�P_UNI�O`_�DO>f7uiFR_F�0AIN�1��x�1c�C_WAkd�a�jOFF_O0N.�DEL�hL� ?a8A�a1b?9a�`FC?��P�1E��#�sATB�d��MyO� �cE D �[M�c��^qRE�V�BILrw!X�I� QrR  �� OD�P�q/$NO^PM�Wp�t�r/"�w� ��u�qJ1X�0D`S� p E RD�_E�pCq$FS�SBn&$CHKBoD_SE^eAG �G�"$SLOT!_��2=�� V�d�%���3 a_ED�Im   � )�"��PS�`(4�%$EP�1�1$�OP�0�2�a�p_�OK�UST1P_�C� ��d��U �PLACI4!�Q�4�<( raCOMM� ,0$D����0�`���EOWBn�IGALL;OW� (K�":(2�0VARa��@h�2ao�L�0OUy�� ,Kvay��PS�`�0M_O]�����CCFS_U	T~p0 "�1�3�#��ؗ`X"�}R0 { 4F IMCM�`O#S�`��upi �	_�p�B}�a����M/ h�pIMPEE_F�N���N���@O��r�D_(�~�n�Dy�F� d�CC_�r0  aT� '��'�DI�Pn0"��p�P줇$I������Fn�t X� GRP0���M=qNFLIx�7��0UIRE���$g"� SWITC�H5�AX_N�PS~s"CF_LIM�� � �0EED��!��qP�t�`�PJ_dVЦMOD�Eh�.Z`�PӺ�ELBOF� ���� ��p� ���3���� �FB/��0�>�G�� �� WARNM�`/��qP���n�NST� CORz-0bFLTRh�/TRAT�PT1�� $ACC1a��N |��r$ORI�lo"V�RT�P_S�� CHG�0I���rT2��1�I��T�m���� x� i#�Q��HDERBJ; CQ�2L�U3L�4L�5L�6L�Q7L� N�9s!�h@{CO`S <F �+�=�O��#92��LL�ECy�"MULTI�b�"N��1�!�Ѻ�0T�� �S�TY�"�R`�=l�)�2`����)�`T  �|� �&$��۱m�0�P�̱�UTO���E��EXT����Á8B���"2� (�
��![0������<�8b+�� "D"�� �ŽQ��<煰kc!(�9�#���1��ÂM8�ԽP��" '�3�$ L� E���P�<��`A�$JOB�n�T���l�TRIG3�% dK��������<���\��+�Y�p�_yM��& t�p3FLܐBNG AgTBA� ���M��
 �!��p� �q��0�aP[`��O�'[����0tna*���"J���_R���CDJ���IdJk�D�%C��`�Z���0���Pq_�P��@ ( @F �RO.��&�t�IT�c�NOM�
�����S���`T)w@����Z�P�d���R�A�0��2b"����
s$T����MD3��T��`U31���p(�5!HGb�T1�*E�7�c�KAb�WAb��cA4#YNT���PODBGD�� *(��PUt@X��W����AX��a��eTAI^cBUF�"0>!+ � 7n�[PIW�*5 P�7EM�8M�9
0�6F�7�SIMQS@>K;EE�3PATn�^��a" 2`#�"�L64wFIX!, ��ֈ!d��D�2Bus=CC9I�:FPCH�P:BAD�aHCEhAOGhAD]HW�_�0>�0_h@ �f�Ak���F�q\'M�`#�""EE3�- l�p3G��@FSOES]FgHBSU�IBS9W|C��. ` ���MARG쀳��F�ACLp�SLEW�xQe�ӿ��M�C�/�\pSM_JBM����QYC	g��e#�0 �n��CHN-�MP�G$G� Jg�_� <#��1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�fJR���rSEG�FR�PIO� S�TRT��N��cP!V5���!41�r�Ӏ
r>İ�b�B�O�2` +�[��� ,qE`�,q`y�Ԣ}t8��yaSIZ%����t�vT�s� �z�y,qRSINF}Oбc����k��`��`�`Lp�ĸ T`7�CRCf�ԣCC/�9��`a�ua8h�ub�MIN��uaPDs�#�G�D�YC��C�����e�q0��� ��EV�q�F�_
�eF��N3�s�ahƔ�Xa+p,5!�#=1�!VSCA?� �A��s1�"!3 ��`F/k��_�U��g���]��C�� a�s���R>�4� �����N����5a�R�HA;NC��$LG��P�6f1$+@NDP�t�AR5@N^��a�q���c��ME�18���}0f��RAө�AZ �𨵰�%O��FCT K��s`"�S�PFADIJ�OJ�ʠ� ʠ���<���Ր��qGI�p�BMP�dp�p�Dba��AES�@�	�K�W_��BAS��� �G�5  zM�I�T�CSX[@�@�!62�	$X����T9�{sC��N��`�~P_HEIG9Hs1;�WID�0�VT ACϰ�1�A�Pl�<���EXP�g���|��CU�0M�MENU��7�T[IT,AE�%)��a2��a��8 P,� a�ED�E.`��wPDT��REM.���AUTH_KEGY  ������ ��b�O	Ѫ�}1ERR9LH� �9 \� �q�-�OR�DB�_IDx�@l �PUN_O��>Y�$SYS0��4�g�-�I�E�EVx�#q'�PXWO��z �: $SK7!�f2.aDBTd�TR�L��; �'AC��`��ĠIND9DIJ.D��_��f1�Ԭf���PL�A�RWAj���SD�A��!�+r|��UMMY9d�F�10dѕ����J�<��}1PR�; 
3�POS��J�g= �$VS$�q�PL~�>��H�SܠK�?����CJ��@����ENE�@TƷ�A���S_�RE�COR��BH �5 O�@=$LA�>$~�r2�R��`��qU�`�_Du��0R	O�@V�T[�Q�U��������! }У�PA�US���dETURYN��MRU� v CRp�EWM�b��AGNAL:s2$�LA�!?$=PX�@$P�y #A �Ax�C0 #ܠDO�`X�k�W�v��q�GO_AWAYƁ�MO�ae���$��DCSS_CCwSCB C �'N��CERI��гJ`u�QAP�}�\�@�GAG� R�0��`��{`��{`O�F�q�5��#M5A��X��H�ш�LL�D� �$���sU�D)E%!`|���OVR10W��,�OR|�'�$E�SC_$`�eDSB#IOQ��l ��B.�VIB&� �c,������f�=pSSW����f!VL��PL|���ARMLO
���`����d7%SC� �bALspH�MPCh �Ch �#h �#
h 5�UU���C�'��C�'�#�$'�d�#C \4�$�pH��Ou��!Y��!�SB���` k$4�C�P3Wұ46�$VOLT37$$`�*�^1���$`O1*�$o��0R�QY��2b4�0DH_THE����0S�<�4�7ALPH�4�`����7�@ �0�qb7
�rR�5�88� ×@���"��Fn�	MӁVHBPFUAF�LQ"D�s�`�THR��i2dB�����G
(��PVP�����������1�J2�B�E�C�E�CPSu�Y@��F b3���H�(V�H:U�G��
X0��FkQw�[�N�a�'B���C INH=BcFILT��� $��W�2�T1�[ @��$���H YАAF�sDO��Y�R p� fg�Q�+�c5h`�Q�iSh�QPL��x�Wqi�QTMOU�# c�i�Q\��X�gmb��Hvi�h�bAi�fI�aCHIG��ca	xO��hܰ��W�"vAN-uX!��	#AV�H!Pa8$P�ד#p�RE_:�A�a��B�qN0�X�MCN�0��f1[1�qVE�p��Z2;&f�I�QO�u�r�x�wGldDN{G|d��aF>!�9��a9M:�U�FWA�:�Ml���X�Lu��$!����!l�ZO����0%�O�lF�s�13�DI�W�@��Q����_��!CURVAL԰0rCR41ͰZ�C <�r�H�v���<�`U�<�(�f�CH�QR3��S���t���Xp�VS!_�`�ד�F��ژ����%҈NS�TCY_ E 	L����1�t�1��U���24�2B�NI O�7������DEVIn|� F��$5�wRBTxSPIB�P���BYX����yT��HNDG��G H tn����L��Q�C���5�:@Lo0 H���閻�FBP�{tFE@{�5�t��T��I��DO���uPMCS��v>�f>�t�"HO�TSW�`s��҈E;LE��J T���e �2��25�� O� ���HA7�E��344�0 � 8���A�K �� MDL� 2J~PE��	A��s��tːÈ�s�JÆG!�rD"�ó�����\�TIO��W�	��5�@�SLAV�L  \0INPڐ���`�%ن_CFd�M�� $��ENU��OG��b�ϑ]զPƟ0`ҕ�]�ID�MA�Sa��\�WR0�#��"]�VE�$a�SKI�STs��sk$��2u���J��������	��Q���_SV>h�EXCLUMqJ2NM!ONL��D�Y���|�PE ղI_V>�APPLYZP���HID-@Y�r�_Mz�2��VRFY�0���r�1�cIOC_�f�� 1������O̥�u�LS���R$�DUMMY3�!����S� L_TP�/Bv�"���AӞ�ّ �N ���RTy_u�� (鵹G&r[�O D��Pw_BA�`�3&x�!F ��_5����H������ �� �P $�KwARG�I��� q�2O ���SGNZ�Q q�~P/�/PIGNs�l�$�^ sQ>ANNUN�@�T`<�U/�ߴ�LAzp�]	Z�d~�����DEFwPI�@ �R @�F?I�T�	$TOTA@%��d���!��EM�NIY�S�+���E�A[�
D7AYS\�ADx�@���	� �EFF/_AXI?�TI��0�zCOJA �ADJ_RTRQ��Up��<P�1D D�r5̀Ll�T�p ? ]P�"p��mtpd��V 0w�G���������SK�SU�� ��CTRL_�CA�� W�T�RANS�6PIDLE_PW���!�4�A�V��V_�l��V �DIAG�S���X� /$�2�_SE�#TAC ���t!�!0z*@��RR��vPA���p ; SW�!�!�  ���ol�U��oOH̅�PP� ��IR�r��BRK'#��"A_Ak���x 2x�9@ϐZs2��%l�W�pxt*�x%RQDW�%3MSx�t5AX�'�"���LIFECAL,���10��N�1{" �5Z�3{"dp5�ZU`^}�MOTN°Y$@���FLA�cZOV�C@p�5HE	��SUPPOQ�ݑAq� aLj (C�1_X6�*IEYRJZRJWRJ�0�TH�!UC��6�XZ_�AR�p��Y2�HCiOQ��Sf6AN�кw$�ICTE��Y `��CACH�E�C9�M�PL{AN��UFFIQ@�Ф0<�1	��u6
�F�MSW�E�Z 8�KEYIYM�p��TM~�S�wQq�wQ#����OC�VIE� �[ �A�BGL��/�}�?M����D?��D\p�mذST��!�R � �T� �T� �T	��PEMAIf�ҁо�_FAUL�]$�Rц�1�U������TRE�^O< $Rc�uS�v% IT��BUFW�}�W��N_� SU	B~d��C|��Sb�q�bSAV�e�bu �B ��� �gX�^P�d�u+p�$�_~`�e�p%yGOTT����sP��aM��OtT�LwAX ě ��X~`9#�c_G:�3
�YN_1�E_�D��1 �2UM���T�F���H@ g�`�� 0p��Gb-sC_R�AIK���r�t��RoQ�u7h�qDS�Pq��rP��A�IM@�c6�\����s2�U�h@�A�sM*`IP��d�s�!D��6�TH�@�n�)�OT�!6�HS{DI3�ABSC���@ Vy��� �{_D�CONVI�AG���@3�~`F�!pd��psq��SC8Z"���sMERk��qcFB��k��pET����aeRFU:@DUdr`����x�CD,�P��@p;cHR�A!���bp�ՔՔ+PUSԕC���C��p�QғSp�cH *�LX�:cd� Rqa�| ����W��U� �U��U�	�U�OQU�7R�8R�9R��0T��^�1k�1x�1��1���1��1��1��1Jƪ2Ԫ2^�k�2x�U2��2��2��2��U2��2ƪ3Ԫ3^�	3k�x�3���o���U3��3��3ƪ4Ԣ��AEXTk!0�d <� 7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr�¸��䂴2REM� F�j��BOVM��A��TROV�DTl�`-�MX<�IN�8�0,�W!INDKЗ�
w�׀�p$DG@~q36��P�5�!D��6�RIV���2�BG�EAR�IO�%K�¾DN�p��J�82���PB@�CZ_MCM��@�1��@U��1�f� ,②a? ����PI�!?I�E��Q���am��©g� _0Pfqg R�I9ej�k!UP2_� h � �cTD �p���! a���i�:w�C�ri T�P�b��`�) OG��%p���p��IFI�!`�pm�>��	�PT�"�EP�FMR2��j ��Ɛ+"�� ��\��������$�B`�x%��_ԡ�ޭ_����� M������D�GCLF�%DGDMY%LDa��5�6H�ߺ4��M���Sk���� T�FS#p�Tl P���e�|qP�p$EX_����1M2��2� 3��5��G ���m� ��Ѝ�SW�eO>e6DEBUG����%GR���pU�#B�KU_�O1'� �@PO�I5�l5MS��OOfswSM��E�bi��0��0_E n ��p `�TERM�o�J`�ORI�+�p�?�SM_����b�q�GN.��TA�r����UP�Rs�s -�1�2n$�>' o$SEG,*> �ELTO��$U�SE�pNFIA�U"4�e1���#$p$UFR���0ؐO!�0̫���OT�'�TA�ƀU�#NST�P�AT��P�"PTH	J����E�P rF�V"ART�``%B`�ab�U!REL:�aSH�FT��V!�!�(_SEH+@M$���� ���@N8r����OVR�q��rSHI%0��UzN� �aAYLO����qIl����!�@��@ERV]��1�?: �¦'�2��%��5��%�RCq��EASY1M�q�EV!WJi'���}�E���!I�2��U�@D��q�%Ba��
5P�o��0�p6OR�MLY� `GR��t2b 5n� � ��%�a�U�u Ԭ")���T�OCO!S�1PO�P ��`�pC��������Oѥ`REPR�3��aO�P�b�"e�PR�%WU.X1��eo$PWR��IMIU��2R_	S�$VIS���#(AUD��LE��Bv" v��$�H���P_ADDR
��H�G�"�Q�Q�Q�БR~pDp1�w H� SZ�a��e�ex�e��SE��r���HS��MNvx ���%Ŕ��OL���p<P��-��ACROlP_!QND_C��ג�1�T� �ROUPT��B_$�VpQ�A1Q�v� �c_��i���i��hx�`�i���i��v�ACk�IOU��D�gfsu<^d�y $|�P�_D��VB`bPR�M_�bi�HTT�P_אHaz (��OBJEr��P��[$��LE�#�s>`{ � ��u��AB_x�T~�S|�@�DBGLV���KRL�YHITC�OU�BGY LO: a�TEM��e�0>�+P'�,PSS|�P��JQUERY_F;LA�b�HW��\!�a|`u@�PU�b�PIO��"�]�ӂ�/dԁ=dԁ�� �IWOLN��}����CXa$SLZ�$INPUT_�$IP#�P��'���SLvpa~��!�\�`W�C-�Bi�IO�p�F_ASv���$L ��w �F1G�U�B0m!���0�HY��ڑ����UOPs� `������@[�ʔ[�і"�[PP�S�IP�<�іI�2���P�_MEMB��i`� X��IP�P�b{�C_N�`����R0�����bSP��p�$FOCUSBG�;� �UJ�Ƃ �  � o7JOG܄'�DIS[�J7��cx�J8�7� I�m!�)�7_LAB�!�@�A��APHMIb�Q�]�D� �J7J\���� _K�EYt� �K^ՀLMONa����$XR��ɀ��WATCH_��3��&�EL��}Sy~���&s� �Ю!V�g� �CTR3򲓥��;LG�D� �R���I�
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�G� �I�F�%SO���q �ƀ����v��ƴ��K�S ����w�k�N����E��\���D'�*�U�s5��@L>�n4�DAUZ�EA�p�Հ�Dp�f�GH�BD��OGBOO���� C���PITp���� ��REC��OSCRN����D_p<�aMARGf�`���:���T�L���S��s��W�Ԣ�Iԭ�J{GMO�MNCH�c���FN��R�Kx�PRGv�UF��p0��FWD��HL��STP��V��+������RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28��2��Gh�0PO���������M8�Ģ��EX.��TUIv�I��(�4�@�t�x�J0J�~�P��J0��N�a�#ANA��O"�0�VAIA��dCLE�AR�6DCS_H�I"�/c�O�O&�SI��S��IGN_�vpq�uᛀ�T�d� DEV-�L1LA �°BUW`Ո�x0T<$U�EM��Ł����0�A�R��x0�σ\�a�@OS1�2��3���@�� `� �ࠜh�AN%-���.-�IDX�DP�2MRaO��Գ!�ST���Rq�Y{b! �$E&C+��p�.&A&d���a� L ��ȟ%Pݘ��T\Q�U�E�`�Ua��_ � �@(��`������# �MB_PN�@ R`r��R�w�TR�IN��P��BAS8S�a	6IRQ6d�{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?��?RIAt,1ID`�D�� d1��RQQp�rpDSTB
`� 1�F�HAXD2��|�G�LEXCES?R��ёBMhPa�͠@�BD4��B�q`�`�F_A�J�C[�Ot�H� K��� \��d�bTf$� ��LI�q��SREQUIRE��#MO�\�a�XDESBU��,1L� M�� �p���P�c��AA,1N��
Q�q�0/�&���-cDC��B�sIN�a?�RSM��Gh� N#B��N�iP�ST9� � 4n��LOC�RI��v�EX�fANG���A,1ODAQ䵗ƞ@$��9�ZMF �����f��"��%u�#ЖVSUP�' ��FX�@IGGo�� �rq�"��1��#B��$���p%#by���rx���vbPDAT	AK�pE;����R���M��*� t�`MD�qI��)�v� �tĀA�wH�`��tDIyA��sANSW�P�th���uD��)�b�ԣ(@$`� PC�U_�V6�ʠ�d�PL�Or�$`�R���B����B�p�����,1R�R2�E�  ���V�A/A d$OCALI�@��G~��2��!V��<$R�SW0^D"���ABC�hD_J2�SE�Q�@�q_J3:M�
G�1SP�,��@PG�n�3m�u�3p
�@��JkC���2'A�O)IMk@{BCS�KP^:ܔ9�wܔJy�{BQܜ������`_AZ.B��?�E�L��YAOCMP0�c|A)��RT�j�ƚ�1�ﰈ��@1�茨����Z��SMG0��pԕ� ER!���aINҠACk�p����b�n _������{A%P4�/R��DIU��C�DH�@
�#a�qc$V�Fc�$x�$���`@���b���̂�E�H ��$BELP����!A/CCEL���kA>°IRC_R�p P��T!�$P)S�@B2L+0����W3�ط9� ٶPACTH��.�γ.�3���p�A_��_�e�-Br�`C���_MG"�$DD��ٰ��$FW�@�p����γ칲��DE��PPA�BN�ROTSPEEu��O0���DEF>Q��+0$OUSE_��JPQP�C��JY����-A 6qYN�@A�L�̐��L�MOU�NG̭�|�OL�y�INCU��a�¢ĻB��ӑ�AENCS���q�B������D�IN�I`�����pzC�VE��<���23_U ��b^�LOWL���:�O0��0�Di�B�P�Ҡ� ��PRC����M3OS� gTMOpp�@�-GPERCH  M�OVӤ ����� !3�yD!e�]�6�<�$� ʓA����LIʓ�dWɗ��:p3�.�I�T3RKӥ�AY���� ?Q^���m�b��`p�CQ�� MOM�B?R �0u��D���y�0�̂��DUҐZ�S_�BCKLSH_C ����o�n��TӀ����
c��CLAL�J��A��/PKCH�KO0�Su�RTY�� �q��M�1�q_�
#c�_UMCP�	C����SCL���LMTj�_L�0X����E�� �� � ��m�h���6��PC����H� �P��2�CN@�"XT����CN_��N^C�kCSF����V6�����ϡj���nCAT�SHs�����ָ1����֙���������P�A���_P���_ P0� e���O1u�$x�JG� P{#�OG|���TORQU(� p�a�~����Ry������"_W��^�����4Pt�
5z�
5I;I ;Iz�F�`�!��_8�1��VC��0�D�B�2�1�>	P�?�B�5JR�K�<�2�6i�DBL�_SM�Q&BMD`_sDLt�&BGRV4`
Dt�
Dz��1H_��8�31�8JCOSEKr�EHLN�0hK�5oDt� jI��jI<1�J�LZ1�51Zc@y��1MYqA�H�QBTHWMYTHE{T09�NK23z��/Rn�r@CB4VCBn�CqPASfaYR<40gQt�gQ4VSBt��RN?UGTS���Cq���a��P#���Z�C$DUu ��R䂥э2��Vӑ��Q�r�f$N	E�+pIs@�|� �	$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b��F�c�j�FR�VrhV�ghd��lV�jV�kV��kV�kV�kV�kV�iHrh�f�r�m!�x��kH�kH�kH�kH��kH�iOclOrhOT��nO�jO�kO�kUO�kO�kO�kO�F�F.bTQ���E��egS�PBALANCEl��RLE�PH_'USP衅F��F��FPFULC�3���3��E��1�l�UT�O_p �%T1T2t���2NW������ǡ��5�`�擳�T��OU���� INSsEG��R�REV���R���DIFH��1ٟ��F�1�;�OB��;C��2� �b~�4LCHWAR���i�ABW!��$MECH]Q�@k�q��AXk�P��IgU�i�� 
���!����7ROB��CR��ͥ�O�C��_s"T� � x $�WEIGHh�9��$cc�� Ih�.�I9F ќ�LAGK�8qSK��K�BIL?�cOD��U��STŰ�P�; �����
�����
�Ы�L���  2�`�"�DEKBU.�L&�n��POMMY9��NA#�δ9�$D&����$��� Q _)�DO_�A��� <	���~��LђBX�P�N��+�_�7�L�t�OH  �/� %��T�����T�����TICYK/�C�T1��%�Ä����N��c�Ã�R� L�S���S�����P�ROMPh�E� $IR� X�~ 8���!�MAI�0��4j���_9����tt�l�R�0COD��sFU`�+�ID_" �=�����G_SU;FF<0 3�O����DO��ِ�� R��Ǔن�S����!{�������	�H)�_F�I��9��ORDfX� ����36h��X�����GR9�\S��ZDTD��|v�ŧ4 *�L_NA4���K��DEF_I[�K��� g��_���i��Ɠ������IS`i �萈�����e����4�0i�Dg�����D� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{ԓ� {ԡ�{����}��v� �Ա��g������^� ��K�Փ����!w�N�P'���^���,`b�W\�[R�?7�sTEFĨ �OULOMB_u��0�VISPI�TY�A�!OY�A�_FRId��(�SI���R�����R�3���W�W���0��0_,�EAS%��!�& "����4p�G;� h� ��7ƵCOEFF_Om���m��/�G!%�S.�߲CaA5����u�GR`� � � $hR� �X]�TME��$R�s�Z�/,)�ER��T;�:䗰�  �]�LL��S�_3SV�($~��q��@���� "�SETU��MEA���Z�x0�u������� � � �� ȰID�"���!*��&"P���*�F�'��A��)3��#����"�5;`*��RE�C���!�t�SKy_��� P	�?1_USER��,���4���D�0��VEL@,2�0���2�5S�I��|��MTN�CFG>}1�  ���=Oy�NORE��3�l�2�0SI���� ��\�UX-�ܑP�DE�A $K�EY_����$gJOG<EנSVIA`�WC�� 1DSWy�x��
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��|�����z�� �@_ERR���! ��S L�-���@���s0BB$BUF�-@X17ࡐMORn�� H	�CU�A 3�z�1Q�
��3���O$��FV��2p0��bG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų7�=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	�����B�t�#}1G� @�@;���OE�RI#A��
N��X��s�f�7���PL}1��,RTv�m�ATUS>RBTRC_T(qR��B �����$ �Ʊ8��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���UP(4����PX��؆�q�3�w� �PG��5� $S�UB������t�J?MPWAITO��s��LOyCFt�!D=��CVF	ь�y���R�`�0��CC_CT�R�Q�	�IGNR�_PLt�DBTB2m�P��z�BW)���2�0U@���IG�a��=Iy�TNLN��Z�R]aK� N��`B�0��PE�s���r��f�S�PD}1� L	�A`�`gఠ�S��UN��{���]�R!�`BDL�Y�2���6�PH_�PK�E��2RETRIEt��2�b���;FI�B� �����8� 2��0DB�GLV�LOGS�IZ$C�KTؑUdy#u�D7�_�_T1@�EM�@C\1aA��ℽR��D�FCHEsCKK�1P�P�0ʳ���@&�(bLE,c�" PA9�T���PJ�C߰PN�����ARh�0���Ӯ�P�O�BORMATTnaF�f1h���2�S��UXy`	��L|B��4�  rE�ITCH3�8PL�)�AL_ � �$��XPB�q� C�,2D�!��+2�J3�D��� T�pPD�CKyp��oC� _AgLPH���BEWQo���� ��I�wp� � �b@PA�YLOA��m�_1�t�2t���J3AR���؀դ֏�laTI�A4��5��6,2MOMCP�����������0BϐAD�����\���PUBk`R�Ԁ;���;���tQ��z4�` I$PI\D s�oӓ1yՕ�w�2�w�UZ��I��I��I�〛�p����n���y��e`�9S)bT�SPEED� G��(�Е�� /���Е�`/�e�>���M��ЕSAMP��6V��/���ЕMO�@ 2@�A��QP�� �C��n����������� LRf`kb�ІE9h�EIN09��7S.�В9
yPy�GA�MM%S���D$GGET)bP�cD]Ԛ�2
�IB�q�IN�G$HI(0;A��$LREXPA8)LWVM8z�)��g���C5�C�HKKp]�0�I_��h`eT��n�q���eT,���� ��$�� 1��iPI� RCH_D`�313\��30LE�1��1\�o(Y�7 �t�M�SWFL �M��SCRc�7�@�&��%�n�f�SV���P�B``�'�!�B�sS_�SAV&0ct5B3NO]�C\�C2^�0� mߗ�uٍa��u���u:@e;��1���8��D�P ���������)� �b9��e�GE�3���V�=��Ml�� � �YL��QNQSRlbfqXG�P �RR#dCQp� �S:AW70�B�B[�CdgR:AMxP�KCL�H����W�r�(1n�g�M�!o�� �F�P@}t$WP�u�P r�� P5�R<�RC�R�� %�6�`��� ��qsr %X��OD�qZ�Ug��ڐ>D� ��OM#w�J?\?n?�?�?0��9�b"���f�]�_��� |��X0 ��bf��qf��q`�ڏgdzf��Eڐ� 5C�Fb�"ɐ���FdPnB��PM�QU��� � 8L�QCsOU!5�QTHI�sHOQBpHYSY�3ES��qUE�`�"��O���  �P��@\�UN���Crf�O�� P���Vu��!����OGR)AƁcB2�O�tVu�ITe �q:pINF�O�����{�qcB�v��OI�r� (�@SLEQS��q��p�vgqS���� =4L�ENABDRZ�PTIONt�����Q���)�GCF�ЎG�$J�q^r�� R���U�g���OS_ED����ѓ �F��PK���E'NU߇وA�UT$1܅COPY������n�00MNx���PRUT8R� �Nx�OU���$G[rf�@bRGAkDJ���*�X_:@�բ$�����P��W��P��} ��)�}�[EX�YCDR��/RGNS.��F@r��LGO�#�NYQ__FREQR�W� 0�#�h�TsLAe#�p���ӄ �CRE� �s�IF��sNA���%a�_Ge#S�TATUI`e#MAIL�����q t��������ELEM��� �/0<�FEASI?�B��n�ڢ@�vA�]� � I�p���Y!q]�t#A�AIBM���E�p<�VΡY�BASR�Z��S�qUZ��0$q�~��RMS_TR;� qb ���SY�	�ǡ��X$���>C�Q`	�? 2� _�T M������̲�@ �Ap��)ǅ�i$DOU�s2]$Nj���PR+@3�=��rGRID�qM�oBARS �TY@�N�OTO�p��� �Hp_}�!����d�O|�P/�� � �p�`POR�s��}��SRV��)����DI&0T����� #�T	�#�4!�5!�6!�%7!�8��F�2���Ep$VALU�t��%��ֱ��/���� ;�.1�q�����(_�AN�#�ғ��Rɀ(���TOTA�L��S��PW�I|l��REGEN�1�cX��ks(��a����`TR��R��_S� ��1ଃV��������Z�E��p�q��Vr����V_H��DA8�S����S_Y,1�R�4�S� AR�P2�� ^�IG_SE�	s����å_Zp��C�_�Ƃ�ENHAN�C�a� T �;�������INT��.��@FPsİ_OVRsP�`p�`��Lv��o��7�}��Z�N@�SLG�AA�~��25�	��D��S,�BĤDE�U������TE�P����# !Y��
�J��$2�IL_MC�x r#_��`TQ�`��q��Ԍ'�BV�C�P_h� 0�M�	V1�
�V1�2�2�3*�3�4�4�
�!����� � m�A�2IN~VIBP��T�1�2�2�3�3�4�4�A@-¸C2���p� MgC_Fp+0�0�L	11d���M50Id�%"E� S`�R/��@KEEP_H/NADD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0��#i��#REM�"@�$��½%�!�(U}��e�$HPWD  �`#SBMSK*|)G�qU2:�P~	�COLLAB� ��!K5�B�� ��g��pITI1{9p#>D7� ,�@FLAP���$SYN �<M��`C6���UP_�DLYAA�ErDE�LA�0ᐢY�`A�D�Q� �QSK;IP=E� ���Xp�OfPNTv�A�0P_Xp�rG�p�RU@,G ��:I+�:IB1:IG�9J T�9Ja�9Jn�9J{�9J�9<��RA=s� X���4�%1�QB>� NFLIC�s�@�J�U�H�LwNO_aH�0�"?��RITu�]�@_PA�pG�QO� ��^�U���W��LV�d�NGRLT�0_q��O�  " 8��OS��T_JvA V�	�APPR_WE�IGH�sJ4CH�?pvTOR��vT��LCOO��]�+�tVJ�Є��ғA�Q�U�S�XO�B'�'�v �J�2P���7�X�T �<a43DP=`Ԡ\"<a8�q\!�RDC��LW� �рR��R�`� �RV��jr�b��RGE��*��cN�F�LG�a�Z���SP9C�s�UM_<`^2TH2NH��P.a� 1� m`E�F11��� l�Q �!#� <�p3AT � g�S��Vr�p�tMq��Lr���HOMQEwr�t2'r�-@?Qcu��w3'r�������w4'r�'�9�K�]�o����w5'r뤏��ȏPڏ����w6'r�!�@3�E�W�i�{��w7'r힟��ԟ����w8'r��-�?�Q�c��u��uS$0�q�p �� sF��`)a�"`P�����`/���-�IO[M�I֠��q�POWE�� ���0Za�0p�� ��5��$DSB� GNAL���0C�pm�S2323�� �~`��� / I3CEQP��PEp���5PIT����OPB�x0��FLOW�@T�RvP��!U���CU:�M��UXT�A��>w�ERFAC�� mU��ȳCH��'� tQ  _��>�f�Q$����OM���A�`T�P#UP%D7 A�ct�T��U�EX@�ȟ�U EFqA: X"�1RSPT�N����T ��PPaA�0o񩩕`EXP��IOS���)ԭ�_`���%��C�WR�A���ѩD�ag֕`ԦF�RIENDsaC2U�F7P����TOOLΫ�MYH C2LE�NGTH_VTE��I��Ӆ$S�E����UFINV�_���RGI��{QITI5B��X�v��-�G2-�G1@7�w�SG�X��_��UQQD=#���AS�Äd~C�`��q�� ��$$C/�S�`������S0S0 }��VERSI� ������5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����S0����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT��C��  ��DI�N�O�A�Dq�EXE��HPV_��AT�Qz
��LARM�RECOV ��RgLMDG �*�5�OLM?_IF *�%�d�O�_�_�_�_j�_�'o9oKo]onm, 
��odb��o�o�o0�o^��$� z, �A   2D{�P�PINFO u[ �Vw��������`����� ��*��&�`�J���n�����DQ���� 
��.�@�R�d�v���𚟬���a
PPLI7CAT��?�P���`Ha�ndlingTo�ol 
� 
V�8.30P/40�Cpɔ_LI
8�83��ɕ$ME�
F0G�4�-
?
398�ɘ��%�z�
7�DC3�ɜ
�No+neɘVr���ɞ_@6d� ~Vq_ACTIVU���C죴�MOD�P���C�I��HGA�PON���O�UP�1*�� Ai�m����Қ_��6��1*�  �@��������Q����Կ�@�
���=�� ���5��Hʵl�K�HTTHKY_��/�M� SϹ���������%� 7ߑ�[�m�ߝߣߵ� ���������!�3�� W�i�{�������� ������/���S�e� w��������������� +�Oas� ������ '�K]o��� �����/#/}/ G/Y/k/�/�/�/�/�/ �/�/�/??y?C?U? g?�?�?�?�?�?�?�? �?	OOuO?OQOcO�O �O�O�O�O�O�O�O_ _q_;_M___}_�_�_��_�_�_�_kŭ�TO�p��
�DO_CL�EAN9��pcNM  !{衮o�o��o�o�o��DSP�DRYRwo��HI��m@�or��� ������&�8�J���MAXݐWdak�H�h�XWd�d��>�PLUGGW�Xg\d��PRC)pB�`E�kaS�Oǂ�2DtSEGF0�K � �+��o�or�����p�����%�LAPO b�x�� �2�D�V�h� z�������¯ԯ�+�TOTAL����+�_USENUO�\�� e�A�k­�RGD�ISPMMC.�2��C6�z�@@Dr\��OMpo�:�X�_S�TRING 1	~(�
�M!��S�
��_ITwEM1Ƕ  n� �����+�=�O�a� sυϗϩϻ����������'�9�I/�O SIGNAL���Tryou�t Modeȵ�Inpy�Simu�lateḏO�ut��OVE�RRLp = 10�0˲In cy�cl�̱Pro?g Abor��̱�u�Status�ʳ	Heartb�eatƷMH �Faul	��Aler�L�:�L�^�p����������� ScûSaտ��-�?� Q�c�u����������� ����);M_q��WOR.�û� �����+ =Oas��������//'.PO����M �6/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�?8�?�?H"DEVP.�0 d/�?O*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8_J_\_n_PALT	��Q�o_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o8�o�_GRIm�û 9q�_as��� ������'�9� K�]�o�������'�R	�݁Q����)� ;�M�_�q��������� ˟ݟ���%�7�I�ˏPREG�^���� [�����ͯ߯��� '�9�K�]�o�������෿ɿۿ�O��$A�RG_� D ?	����0���  	]$O�	[D�]D���O�e�#�SBN_�CONFIG �
0˃���}�C�II_SAVE � O�����#�T�CELLSETU�P 0�%  ?OME_IOO�O�%MOV_H������REP��J��UTOBACK�����FRwA:\o� Q�,o���'`��o����� ��  f�o�����*�!�3�`��Ԉ��f���� ������o�{��&�8� J�\�n���������� ��������"4FX j|�������끁  ��_�i�_\ATBCK�CTL.TMP �6.VD GIF? .TP D_8q��NLQ���.f�INI�P�Օ��c�MESSAG�����8��ODEC_D����z��O�0��c�PAUSM!!��0� (783�U/g+(Od/�/ x/�/�/�/�/�/�/? ??P?>?t?1�0$: ?TSK  @-��<T�f�UPDT���d�0
&XWZD�_ENB����6S�TA�0��5"�XI�S��UNT 2�0Ž� � 	 ���z���eng��-뷛�S��o�U@��H�����zF�Oo�}Cw�gJ�^����.�O��O�O�O/_2FMET�߀2CMPTAA���@�$A�-�@���@����@���]5���5�(d5���P5�r�5F*5�338]�SCRDCFG }1�6��	��Ź�_�_oo (o:oLo��o�Q���_ �o�o�o�o�o�o]o �o>Pbt���o9�i�GR<@M/��s/NA�/�	�i��v_ED�1��Y� 
 �%{-5EDT-��'�GETDATAU�o�9��?�j�H�o�f�\��A�^�  ���2�0&�!�E���:IB����~�ŏ׏m����3 ��&۔��D��ߟJ� ����9�ǟ�4��� ϯ�(����]�o�����5N������(��w��)�;�ѿ_��6 ϊ�gϮ�(�CϮ���ϝ�+��7��V�3� z�(��z�����i���B�8��&���~�]����F�ߟ�5����9~������]����`Y�k�����CR� !ߖ���W�q���#�5����Y��p$�NO_D�EL��rGE_U�NUSE��tIG�ALLOW 1���(*S�YSTEM*S�	$SERV_G�R�V� : REGƟ$�\� NU�M�
��PMU|B ULAYNP�\PMPA�L�CYC10�#6 $\UL�SU�8:!��Lr�BOXOR=I�CUR_���PMCNV��10L�T4�DLI�0��	�� ��BN/`/r/�/�/�/�/�/���pLAL_?OUT �;����qWD_ABOR�=f�q;0ITR_�RTN�7�o	;0NgONS�0�6 
H�CCFS_UTI�L #<�5CC�_@6A 2#; h ?�?�?O#O6]�CE_OPTIO�c8qF@RI'A_Ic f5Y@�25�0F�Q�=2qz&}�A_LIM��2.� ��P��]B��KX�P
��P�2O�Q��B�r�qF�PQ5T1�)TR�H�_:JF_�PARAMGP 1�<g^&S�_��_�_�_�VC�  +C�d�`�o!o�`�`�`�`�Cd��Tii:a:e>e�Ba�GgC�`� D_� D	�`�w�?��2HE ON�FI� E?�aG_Pv�1#; � ��o1CUg|y�aKPAUS�s1�yC ,�� �������	� C�-�g�Q�w�������Ы�я���rO�A��O�H�LLECT�_�B�IPV6�ENp. QF�3�NDE>�� �G�71�234567890��sB�TR����%'
 H�/%)�� �����W���0�B��� f�x���㯮���ү+� ����s�>�P�b��� �������ο��Kπ�(�:ϓ�^�|��B!�F� �I|�IOG #��<U%e6`�'�9�K���TR�P2$��(9X�t�Yކ�`%�̓ڥH��_�MOR�3&�=�>�@XB��a� �A�$��H�6�l�~���~S��'�=�r_A? �a�a`��@K��RʭdP��)F�haÃ-�_�'�9�%
@�k��G� ��%Z�^%��`�@c.��PDB��+���cpmidbg��X	�`:��0!�0�"QU��p��N�  ��@3�@4b/���]ܭ@�v5w<�^�,`@`�wg�$V� �@wf�l�q��ud1�:��:J��DEFg *ۈ��)��c�buf.tx�t����_L64FIX ,�� ����l/[Y/�/}/�/ �/�/�/
?�/.?@?? d?v?U?�?�?�?�?�?��?,/>#_E -���<2ODOVOhOzO��O6&IM��.o�YU>���d�
�I�MC��2/����dXU�C��20�M�QT|:Uw�Cz  B��i�A���A����Au�gB3��*CG�B<��=w�i�B.��B����B��5B��$�D�%B���ezVC�q��C�v�D����D-lE\D�n �k��B9"6��22o�D|�KU ���� �� -����
�xObi�Dv ebv`D��`/��`v`s]E�D D��` E4�F�*� Ec��F�C��u[F���E���fE��fF�ކ3FY�F��Pr �X��@�3�3 ;��>L̩��Aw�n,a@��@e�5Y���a���`�A��w�=�`<#����
��?�ozJRS�MOFST (X�,bIT1��D @3��
д����a���;��bw?����<�M�NT�EST�1O�CR�@�4��>VCv A�w�Ia+a�aORI`mCTPB�U�C�`�4���r��:d�T���qI?�5��q�T_�PROG 	��
�%$/ˏ�t��NUSER  �U�������KEY_?TBL  �����#a��	
��� !"#$%&'�()*+,-./���:;<=>?@�ABC�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~��������������������������������������������������������������������������������͓���������������������������������耇���������������������9�����LCK�
�<���STAT/��s�_AUTO_DO�+ ��[�INDT_'ENBP���Rpqn��`�T2����STO�r`���XC�� 2�6���8
SO�NY XC-56t�"b����@��F( А�HR50w���>�P�y7b�t�Aff����ֿ� Ŀ���� C�U�0�yϋ�fϯ��π���������-ߜ�T{RL��LETEͦ� ��T_SCR�EEN ��Okcs���U��MMENU 17�� <ܹ��� w���������K� "�4��X�j���� ��������5���k� B�T�z����������� ����.g>P �t����� �Q(:�^p ����/��;/ /$/J/�/Z/l/�/�/ �/�/�/�/�/7?? ? m?D?V?�?z?�?�?�? �?�?!O�?
OWO.O@O�fO�OvO�O�O(y��REG 8�y�����`�M�ߎ�_MA�NUAL�k�DB;CO��RIGY�9��DBG_ERRL&��9�ۉq��_��_�_ ^QNUMSLI�pϡ�pd
��
^QPXWORK 1:���_5oGo�Yoko}oӍDBTB�_N� ;������ADB_�AWAYfS�qG�CP 
�=�p�f_CAL�pR��bbRY��[�
�WX_�P 1<
{y�n�,�%oc��P��h_M��IS�O��k@L��sONT�IMX��
����vy
��2sMOT�NEND�1tRECORD 1B��� ���sG�O�]�K��{�b������ ��V�Ǐ�]����6� H�Z���������#� ؟������2���V� şz��������ԯC� ��g��.�@�R���v� 寚�	���п���c� χ�#ϫ�`�rτϖ� Ϻ�)ϳ�M���&� 8ߧ�\�G�Uߒ�߶� ����I������4�� �p7�n���ߤ�� ��������"���F� 1���|��������[� ����i���BTf����bTOLER7ENC�dB�'r�`�L��^PCSS_�CCSCB 3C$>y�`IP�t}�~ �<�_`r� K�����/�{��5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O`�O�O_�~�LL� D��&qET�c�a� C[C�p�PZP^r_ A� %p� �sp��QGPt[	 A�p�Q�_��[? �_�[oU��p�P�pSB� V�c�(a�PWoio{h+�o�X�o�o�Y��[	r�hLW���N:p����}6ڿ��c��aD�@VB��|��G���+��K� �otGhXGr�So�����eB   =��eͶa>�tYB�� ��pC�p�q�aA"�H �S�Q-��q���ud��v�����AfP ` 0���D^P��pk@�a
�QXT�HQ����a aW>� �a9P��b�e:�L�@^�h�Hc�́PQ�R FQ�PU�z�֟�o\ ^��-�?��c�u���,�zCz�ů�b�2�Щ�RE����D��v����S ̡0��]�0�.��@���EQ�p��F�X�ѿ�Uҁп�VSȺNSTCY 1E�
�]�ڿ��K�]� oρϓϥϷ������� ���#�5�G�Y�k�}���ߒ��DEVIC�E 1F5�  MZ�۶a��	� ��?�6�c���	{䰟����_HNDGD �G5�VP���R�LS 2H�ݠ��/�A��S�e�w����� ZPA?RAM I�Fg�He�RBT 2-K��8р<��WPVpC�C��,`¢PQ�Z�z��%{�C*  �2�jMT`LU,`"nPB,  s��M� }�gT�g���
B��!�bc y�[2Dchz ����/��/�gT#I%D��C��` b!�R��A���A,��Bd�ךA��P��_C4kP�!2�C��$Ɓ�]ߚffA�À�W�B�� �| ���/�/�T (��54a 5�}%/7/d?/M? _?q?�?�?�?�?�?O �?OO%O7OIO�OmO O�O�O�O�O�O�O�O J_!_3_�_�_3�_�_ �_�_�_o�_(ooLo ^oЁ=?k_IoS_�o�o �o�o�o�o�o# 5G�k}��� ����H��1�~� U�g�y�ƏAo�Տ� ��2�D�/�h�S���go ����ԟ����ϟ�� �R�)�;���_�q��� �������ݯ�<�� %�7�I�[�m������� ��}�&��J�5�n� YϒϤϏ��ϣ�ѿ� �����F��/�Aߎ� e�w��ߛ߭������� ��B��+�x�O�a�� ����������,��� %�b�M���q������� ��������L# 5�Yk}���  ��61C Ug������ ��	//h/���/w/ �/�/�/�/�/
?�/.? @?I/[/1/_?q?�? �?�?�?�?�?�?OO %OrOIO[O�OO�O�O �O�O�O&_�O_\_3_ E_W_�_?�_�_�_�_ �_"ooFo1ojoE?s_ �_�om_�o�o�o�o�o 0f=Oa� �������� �b�9�K���o���Ώ ��[o��(��L�7��I���m������$D�CSS_SLAV�E L����ё��__4D  љ�◿CFG Mѕ��������_FRA:\ĐL-��%04d.CSVn��  }�� ���[A i�CHq�z�������|�����  �����Ρޯ̩ˡ�Ґ-��*����_�CRC_OUT �N������_�FSI ?њ ����k�}� ������ſ׿ ���� �H�C�U�gϐϋϝ� ���������� ��-� ?�h�c�u߇߽߰߫� ��������@�;�M� _����������� ����%�7�`�[�m� ��������������� 83EW�{� ����� /XSew��� ����/0/+/=/ O/x/s/�/�/�/�/�/ �/???'?P?K?]? o?�?�?�?�?�?�?�? �?(O#O5OGOpOkO}O �O�O�O�O�O _�O_ _H_C_U_g_�_�_�_ �_�_�_�_�_ oo-o ?ohocouo�o�o�o�o �o�o�o@;M _������� ���%�7�`�[�m� �������Ǐ����� �8�3�E�W���{��� ��ȟß՟���� /�X�S�e�w������� �������0�+�=� O�x�s���������Ϳ ߿���'�P�K�]� oϘϓϥϷ������� ��(�#�5�G�p�k�}� �߸߳����� ���� �H�C�U�g���� ���������� ��-� ?�h�c�u��������� ������@;M _������� �%7`[m ������� /8/3/E/W/�/{/�/ �/�/�/�/�/??? /?X?S?e?w?�?�?�? �?�?�?�?O0O+O=O OOxOsO�O�O�O�O�C��$DCS_C_�FSO ?�����A P �O�O_?_ :_L_^_�_�_�_�_�_ �_�_�_oo$o6o_o Zolo~o�o�o�o�o�o �o�o72DV z������� 
��.�W�R�d�v��� ����������/� *�<�N�w�r������� ��̟ޟ���&�O� J�\�n���������߯ گ���'�"�4�F�o� j�|�������Ŀֿ�������G�B�T��OC/_RPI�N_j� �����ς��O����1�XZ�U��NSL��@&� h߱���������"�� /�A�j�e�w���� ����������B�=� O�a������������� ����'9b] o������� �:5GY�} ������// /1/Z/U/g/y/�/�/ �/�/�/�/�/	?2?-? ??Q?z?u?��ߤ߆? �?�?�?OO@O;OMO _O�O�O�O�O�O�O�O �O__%_7_`_[_m_ _�_�_�_�_�_�_�_ o8o3oEoWo�o{o�o �o�o�o�o�o /XSew��� �����0�+�=� O�x�s���������͏ ߏ���'�P�K�]��o����� �PRE_?CHK P۪��A ��,8��2��� 	 18�9�K���+�q� ��a�������ݯ�ͯ �%��I�[�9���� o���ǿ��׿���)� 3�E��i�{�Yϟϱ� ������������-� S�1�c߉�g�y߿��� �����!�+�=���a� s�Q�������� ������K�]�;��� ��q������������� #5�Ak{� ����� CU3y�i�� ����/-/G/ c/u/S/�/�/�/�/�/ �/??�/;?M?+?q? �?a?�?�?�?�?�?�? �?%O?/Q/[OmOO�O �O�O�O�O�O�O_�O 3_E_#_U_{_Y_�_�_ �_�_�_�_�_o/oo SoeoGO�o�o=o�o�o �o�o�o=- s�c����� ��'��K�]�woi� ��5���ɏ������� �5�G�%�k�}�[��� ����ן�ǟ���� C�U�o�A�����{��� ӯ����	��-�?�� c�u�S�������Ͽ� ������'�M�+�=� �ϕ�w�����m���� ��%�7��[�m�K�}� �߁߳��߷����!� ��E�W�5�{��ϱ� ��e�������	�/�� ?�e�C�U��������� ������=O- s����]�� ��'9]oM �������/ �5/G/%/k/}/[/�/ �/��/�/�/�/?1? ?U?g?E?�?�?{?�? �?�?�?	O�?O?OO OOuOSOeO�O�O�/�O �O�O_)__M___=_ �_�_s_�_�_�_�_o �_�_7oIo'omoo]o �o�o�O�o�o�o! �o1W5g�k} ������/�A� �e�w�U�������я ��o����	�O�a� ?�����u���͟��� ��'�9��]�o�M� ��������ۯ��ǯ� #�ůG�Y�7�}���m� ��ſ�����ٿ�1� �A�g�E�wϝ�{ύ� ������	�߽�?�Q� /�u߇�e߽߫ߛ��� �����)���_�q� O���������� ���7�I���Y��]� ��������������! 3WiG��} ����%�A �1w�g��� ���/+/	/O/a/ ?/�/�/u/�/�/�/�/ ?�/9?K?�/o?�? _?�?�?�?�?�?�?O #OOGOYO7OiO�OmO �O�O�O�O�O_�O1_ C_%?g_y__�_�_�_ �_�_�_�_o�_+oQo /oAo�o�owo�o�o�o �o�o);U__q ������� �%��I�[�9���� o���Ǐ�����ۏ!� 3�M?�i��Y����� ��՟�ş����A� S�1�w���g�����������ӯ�+�=��$�DCS_SGN �QK�c��7m�� 13-F�EB-19 13?:48   O�l��4-JANt�08�:3|����� N.DѤ����������h�x,rWf*σ�^M���  O�VERSI�ON [�V3.5.13��EFLOGIC �1RK��?  	���P��?�P�N�!�PROG_ENB  ���6Ù�o�ULSE�  TŇ�!�_�ACCLIM�����Ö��WR�STJNT��c��K�EMOx̘���� ���INIT �S.�G�Z���OPT?_SL ?	,���
 	R57Y5��Y�74^�6_ح7_�50��1��2�_�@ȭ��<�TO C Hݷ���VЗDEX��dc�����PATH A[�A\�g�y���HCP_CLNT�ID ?��6� �@ȸ����IA�G_GRP 2X�K� ,`���� �9�$��]�H�����12�345678908����S�� |��������!��  ��H���;�dC�S���6����� .�Rv�f ��H��//� </N/�"/p/�/t/�/ �/V/h/�/?&??J? \?�/l?B?�?�?�?�? �?v?O�?4OFO$OjO |OOE��Oy��O�O _�O2_��_T_y_d_t�_,
�B^ 4�_ �_~_`Oo�O&oLo^o I��Tjo�o.o�o�o�o �o �O'�_K6H �l������ �#��G�2�k�V����B]�?�  �7����O�L���޷��LS.��/K�Q;ƁDrx�@��PC����� �Ƈ����(��L�B\�ډ�4  79���$��>���:������ߟʟܟ���C�T_CONFIG� Y��Ӛ��egU���ST�BF_TTS��
@��b����Û�u�O��MAU��|��MS�W_CF6�Z�� � �OCVIE�W��[ɭ��� ���-�?�Q�c�u�G� 	�����¿Կ����� �.�@�R�d�v�Ϛ� �Ͼ�������ߕ�*� <�N�`�r߄�ߨߺ� ��������&�8�J� \�n���!������ �������4�F�X�j�X|����RC£\�e��!*�B^�������C2g{�SBL�_FAULT �]��ި�GPMS�Kk��*�TDIAOG ^:�աI���UD1: �67890123C45�G�BSP� -?Qcu��� ����//)/;/(M/tJ��
@q�|�/$�TRECP��

��/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO�i/{/xO�/UMP_?OPTIONk��F�ATR¢l��	�E�PMEj��OY_T�EMP  Èϓ3B�J�P�AP�DUNI��m�Q���YN_BRK �_ɩ�EMGDI_STA"U�aQ�SUNC_S1`ɫ C�FO�_�_�^
�^dpOoo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �E�����y�Q� �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d��z��� ����˟����%� 7�I�[�m�������� ǯٯ����!�3�E� W�i���������ÿݟ �����/�A�S�e� wωϛϭϿ������� ��+�=�O�a�{�i� �ߩ߻�տ������ '�9�K�]�o���� �����������#�5� G�Y�s߅ߏ�����i� ������1CU gy������ �	-?Qk�}� ��������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?u?�?�?�? ��?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_m? w_�_�_�_�?�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9Ke_W��� �_�_����#�5� G�Y�k�}�������ŏ ׏�����1�C�] oy��������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;���g�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� _�i�{ߍߟ߹����� ������/�A�S�e� w����������� ��+�=�W�E�s��� ���ߧ������� '9K]o��� �����#5 O�a�k}�E��� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-?GYc?u? �?�?��?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_Q?[_m__�_�?�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/I_Se w��_����� ��+�=�O�a�s��� ������͏ߏ��� '�A3�]�o����� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����9�K�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� ߑ�C�M�_�q߃ߝ� �߹���������%� 7�I�[�m����� ���������!�;�E� W�i�{��ߟ������� ����/ASe w������� 3�!Oas�� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?+= G?Y?k?!?��?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	_#?5??_Q_c_u_ �?�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o-_ 7I[m�_��� �����!�3�E� W�i�{�������ÏՏ ����%/�A�S�e� q�������џ��� ��+�=�O�a�s��� ������ͯ߯��� �9�K�]�w������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� �������'�1�C�U� g߁��ߝ߯������� ��	��-�?�Q�c�u� �����������m� �)�;�M�_�y߃��� ����������% 7I[m��� �����!3E Wq�{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ �/+?=?O?i_?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O�O�O�O�O? �$�ENETMODE� 1aj5_�  00�54_F[PRRO�R_PROG �%#Z%6�_�YdUTABLE  #[�t?�_�_�_gdRSEV_NUM 2R  �-Q�)`dQ_AUTO_?ENB  PU+S�aT_NO>a b�#[EQ(b  *U��`��`��`��`�4`+�`�o�o�oZdH�IS%c1+PSk_A�LM 1c#[ e�4�l0+�o�;M_q���o_\b``  #[a�FR�zPTCP_V_ER !#Z!�_��$EXTLOGo_REQ�f�Qi�,�SIZ5�'�ST�KR�oe�)�T�OL  1Dz��b�A '�_B�WD�p��Hf��D�_�DI�� dj5�SdDT1KRņST�EPя�P��OP�_DOt�QFAC�TORY_TUN��gd<�DR_GR�P 1e#YNad �	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ�ԟ��� 1��U�@�y�d�v������ӯ����LW
 �J}8*�,��t�ۯ�j�U���y�B��  B୰���$�  A@��s�@U�UUӾ�������Eﻀ E�`F@ F�5U/�,���L���M���Jk�Lzp��JP��Fg�f��?�  s��9��Y9}�9���8j
�6��6�;���A���O ���� � I ������[�FEATURE �fj5��JQ�Handlin�gTool � �"
PEn�glish Di�ctionary��def.4�D St�ard��  
! h�Analog �I/OI�  !�
IX�gle S/hiftI�d�X��uto Soft�ware Upd�ate  rt �sѓ�matic �Backup�3�\st��gr�ound Edi�t��fd
Camera`��Fd�e��CnrROndIm���3��Common calib UI��_ Ethe�n���"�Monitor��LOAD8�tr~�Reliaby��O�ENS�Data Acquis>���m.fdp�ia�gnos��]�i�D�ocument �VieweJ��8�70p�ual �Check Saofety*� cy�� �hanced Us��Fr�����C �xt. DI�O :�fi�� m�8���end��ErrI�L��S������s  t Pa��r[�� ���J9�44FCTN_ Menu��ve��M� J9l�TP �InT�fac{� � 744��G��p� Mask Ex�c��g�� R85��T��Proxy� Sv��  15� J�igh-S�pe��Ski
� �R738Г��m�munic��on�s�S R7��uqrr�T�d�022���aю�connecwt 2� J5���Incr��str�u,Қ�2 R�KAREL Cmod. L��ua���R860hRunw-Ti��EnvL��oa��KU�el u+��s��S/W����7�Licensye���rodu� �ogBook(S�ystem)�A�D pMAC�ROs,��/Of�fs��2�NDs�M�H�� ����M�MRC�?��ORD�E� echSto�p��t? � 84�fMi$�|� 13dx��]е�׏����Modz�witc�hI�VP��?��.� sv��2Op�tm�8�2��fi�l��I ��2g �4 !+ulti�-T�����;�PCM funY�Po|���4$�b&/Regi� r �Pri��FK+7����g Num Se-lW  F�#��� Adju���6�0.��%|� fe<���&tatu�!$�6���%��  9 �J6RDM �Robot)�sc�ove2� 561N��RemU�n@�� 8 (S�F3Se�rvo�ҩ�)�SNPX b<�I�\dcs�0}��Libr1��H� �5� f�0��[58��So� tr��ssag4%G 91��p ��&0����p/I��  (�ig TMILIBx(MӋ�Firm�����gd7���s�Ac�c����0�XATX��Heln��*LR�"1��Spac��Arquz�imu�laH��� Q���Tou�Pa��I���T��c��&��ev�. f.sv?USB po��"��iP�a��  r�"1Unexcep�t��`0i$/����H[59� VC&�r��[6���P{��RcJ�PRIN�V�; d� T@�TSP C�SUI�� r�[X�C��#Web P9l6�%d -c�1R�@4d�����I�R66?0FV�L�!FV�GridK1play C�lh@���і5RiR�R.@���R-35iA���Ascii���"�η� 51f�cUp9l� � (T�����S��@rityA?voidM �`���CE��rk�C�ol%�@�GuF� 5P��j}P����
 B�zL�t� 120C C� o�І!J��P�Бy��� o=q�b �@DCS b ./��c��O��q��`�;� ���qckpaboE4�DH@�OT�~��main N��r�1.�H��an.�t�A> aB!FRLM����!i ���MI 7Dev�  (�1�G h8j��spiJP@��� �@��Ae1/�r����!hP� M-A2� i��߂^0i��p6�PC��  �iA/'�Pass�wo�qT�ROS� 4����qeda�SN��Cli�����G6x Ar�� 47��!���5s�DER\��Tsup>RtОI�7 (M�a�T2�DV�
�3D Tri-���&��_�8;�
�A�@Def�?����Ba: d7eRe p 4t0���e�+�V�st6�4MB DRAM��h86΢FR�O֫0�Arc� v#isI�ԙ�n��7|� ), �b�He�al�wJ�\h��C'ell`��p� �sh[��� Kqw�c�� - �v���pX	VCv�tyy�s�"^Ѐ6�ut� �v�m���xs ���TD_0��J�m�` �2��a[�>R ts=i�MAILYk��/F2�h��ࠛ 9�0 H��F02]�q2�P5'���T1C��5�����FC��U�F�9�GigEH�S�t8�0/A� if�!2v��boF�dri=c� �OLF�S�����" H5k�OgPT ��49f88���cro6���@��l�ApA�Sy�n.(RSS) �1L�\1y�rH�L� �(2x5�5�d�pCV�x9����est�$S�Р��> \pϐSS�F�e$�tex�D �o���A�	� BP����a�(R00�Qi#rt��:���2)�D���1�e�VKb@l �Bui, n��WACPLf��0��Va��kT�XCGM��D��L8����[CRG&a&�YBU��YKfL�p�pf��k�\sm�ZCTAf�@�О�Bf2�и��V#�s���� r���CB���
Pf���WE��!��
���T�p��DT�&4 Y�V�`���EH����
�61�Z��
�R=2�
�E 	(Np��F�V�PK�B����#��Gf1`?GD���H�р?I�e ����LD�L��N��7\s@���`����M��dela�<,��2�M�� "L[P��`?��_P�%�����S��-F��TSO�W�J5�7��VGF�|�V;P2֥ 5\b�`0�&�cV:���T;T�� �<�ce,?V{PD��$
T;YF��DI)�<I�'a\so<��a-�6J�c6s6�4L�M�V9R�h���Tri�� ���5�` �f�@��������P
� ����`��IOmg PH�[l�6�I/A  VP�S��U�Ow��!%S|�Skastdpn)���t�� SWIMEkST�BFe�00��-Q� �_�PB�_�RGued�_�T�!�_��S ��_bH573�o2c2��-oNbJ5�N�Iojb)�Cdo�cx E��o�_�lp��o�TdP �o�c�B�or�2.r�ٱ(Jsp�EfrSE�o�f1�}�r3 R�GoeELS��sL ����s�����B	�0�S\ $�F�ryz�ftl�o~�g�o����������?�����P   �n�&�"�l ��T �@<�^��Y��e�uy8Z���alib���Γ��ɟ3���埿�\v ��e\c�6�Z�qf�T�v�R VW�r��8S��UJ91��0��i�ů[c91+o�wy8���847� :��A4�j��Q��t6�<m���vrc.����0HR���ot�0ݿN��  ��8ޯf�460�>eS0L�97���U�ЄϦ�60.� g�н�+���'�ܠ�Ϻ�8co��D	M߱U"�����ߕp�i�߲T! ��n	a;�� ���u%��ⅰI��loR�d��1a59gϱŭ�&��95�ϔ�R����1��?��o�#��1A��/���vt{�UWe0ǟ���ￇ73[���97�ρ�C W���62K�=fR���8���������d����2 �ڔ����@�@y" "http������t7 �� v 3R7��78�����4�� ��TTPT��#	��ePCV�4/v߀�j�Q�Fa�7��$N�0�/2�rI�O�)/;/M/6.sv�3�64i�oS�l? torah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4c.K?�g'�)�s24g?�� (B�O�d�\iOA5sb�?U_�?vi�/i��/��/Wn��`�o%�F o�4l�$of��oXF� I)xo�cmp\�7��mp���duC`��lh����o(A�_Bt� �o]6P��m�I?0�w�@���naO��	4*O0wi�%P�?"�bsg?�]7�YE$M���8woVJ�/ե311?o��DMs�BC��7J�\���r(�52�XFa AP��ڟ<�v�`/şaqqs����/Of���1�9�VR`K���ph�քH5+��=�IN/¤SkiW�/�IF��_�%��fs�I�O�l����"<𜿚$�`�����\jԿz5bO�vr�ouς�3(�ΤH (DϮ��?sG��|� �F�Ou�������D)O��*�3P$�FӅ�@k��ϻ���럴� �P�L��ʿ��pbox��ߦebo���Sh$ �>�R.�0wT{����fx6��P��D`��3��#_I\m;YEe�OԆM�hxW��=Ete,���dct\���O$kR���d���Xm*���ro30��D�l�j9��Vx'�  FC����|@�ք f?6K�ARE0�_�~ (1Kh��.cf����WpoO�_K�up���a���H/j#- 3Eqd/�84���$qu�o��/ o2o?DVo<�7C�)�s�NJ�Ԇ�|?�3l\sy`�?�40�?Τwio��u]?�w58�?,F�a$OJ�
?Ԇ"io��!�V��u&A��P�R�ߩ5, s��v1�\  Hg552B�Q21p�0R78P5�10.R0  n�el J61�4Ҡ/WA�TUP��d8P54�5*�H8R6��9_VCAM�q97P�CRImP\1tPUI�F�C8Q28  i�ngsQy0��4P P6�3P @P PSCH~��DOCVڀD �PCSU���08Q�0=PqpVEIcOCr��� P54Pwupd�PR69aP܄��PSET�pt\!hPQ`Qt�8P7`Q�!?MASK��(P?PRXY���R�7B#POCO  /\pppb36���@PR�Q��b1Pd60Q^$cJ539.eHsb~��vLCH-`~(�OPLGqK\bPQ0]`��P(`GHCR��4`S�awund�PMCSIPR`e0aPle5=Ps�p(`DSW� �  qPb`0`�aPa��(`PRQ``Tq�RE`(Poa601P�<cPCM�PHcR0@q\j23b�V�`pE`�S`UPvisP�`E` c�`UPcPR9S	a�bJ69E`s�FRDmPsRMC�N:eH931PHcS�NBARa�rHLB��USM�qc�Pg5�2�fHTCIP0cT�MIL�e"P�`eJ� �PA�PdSTPT�X6p967PTEL��p��P�`�`
Q8P8$Q48>a"PPX�8Pc95�P`[�95qq�bUEC-`F
�PUFRmPfahQCvmP90ZQVCO�`�@PVIP%�53�7sQSUIzVSX��P�SWEBIP�SH�TTIPthrQ6�2aP�!tPG���cI�G؁�`c�PGSξeIRC%��cH7�6�P�e Q�Q|�Ror��R51P s:PL�P,t53=P8u8=P
y�C�Q6]`�b�P�I��q52]`sJ5�6E`s���PDsCLt�qPt5�\rd�q375UP cR8���u95P sR55]`,s � P8s��P�`CP�P�P�SJ77P0\o�6��cRPP�cR6�ap�`�QtaT�379P`�64�Pd387]`�d90P0c ��=P,���5�9ta�T91P� ��1P(Sܒ��Qpai�P06�=P- C�PF�T`	���!aLP PTS�p.L�CAB%�I Б�IQ` ;�H�UPPa[intPMS�Pa�иD�IP|�STY%�t7\patPTO�b8�P�PLSR76�`�5�Q��WaNN�Pa�ic�qNNE`�OsRS�`�cR681Pwint'�FCB�P"(�6x�-W`M�r���!(`OBQ`pluug�`L�aot �`GOPI-���PSP�Z�PPG�Q7�`7�3ΒPRQadv�RL��(Sp�P�S��n�@�E`��� �PTS-��q W��P�`apw�`8��P`cFVR�Plc�V3D%�l�PBV�I�SAPL�Pcy�c+PAPV1�pa�_�CCGIP - uU��L�Prog+PGCCR�`�ԁB�Pi �PԁK=�"L�PH��p��(h�<�P���h�̱�@g�Bـ
�TX�%���CTC��ptp��2��P927"0ҝPs2�Qb��;TC-�rmt;�	`�#1ΒTC9`HcC[TE�Perj�EIPp.p/�E�P�c�ЮI�use��Fـverv�F%���TG�Pp� CP��%�d -h��H-�Tra�PCT�I�p��TL� TRS���p�@נ��IP�PTh�M%�lex�sQTMQ`ver, �p�SC:���F��P�v\e�PF�IPSV�"+�H�$cj�ـtr��aCTW-���CPVsGF-��SVP2mPOv\fx���pc�bؚ�e��bVP4�fx�_m��-��SVPD�-��SVPF�P_m�o�`V� cV��t�\��LmPove4���-�sVPR�\t|�tPV�Qe5.W`V6�*u"��P}�o`�М�`��CVK��N�I�IP��CV����IP=N9�Gene���D���D�R�D����  ��f谔�pos.^��inal��n�D�DeR���`��d�P��omB���on,����R�D�R��\��T�Xf��D$b��omp��� "N��P��m����! ��=C-qf����=FXU�����g F��(��Dt II��r�D���u�� "����Cx_ui X�������f2��h	Crl02��D,r9ui�Ԣ>� it2c�0�co��e"���Խا(.)� ����� ���� IQnQ �{I[ ��_= �wo��,bD�� ��|GG�� �����{4 �e� �vʷ� ��&�� 2��Z u{z������ ��TW&q~q� 5�׷&�o�? ;0��  ��2� �y�� ���W&��� ?�3� {A��e�/> ��\�3&T���� 77߸ ��{�� ���� �ֵ��&��8� �l1��S��) ���d *�J� F's� ~��� 6:0ݙ ��,��s�{�- Q�v� ���� �,սT �ZBLx6�ۯ�6 ��6����Par ��s�>�E��j�6dsq��F  ���������Dhel�����ti-S�� �Ob��Dbcf�O���V��t OFT��P< A�_�V�ZI��D���V\�qWS��= d7tle�Ean�(b{zd��titv�JZ�z�Ez XWO� H6�6���5 �H�6H691�E4܀TofkstF� Y�682�4�`�f8�04�E91�g�`3<0oBkmon_�E��xeݱ�� qlm��W0 J�fh��B�__  ZDTfL0��f(P7�Eckl`KV� �6|��D85��ّ�m\b����xo܊k�ktq��g2`.g���yLbkLV�ts��IF�bk������Id I/�f��GR� �han�L��Vy��%���%ere�����io��� ac�- A��n�h���cuA2Cl�_�^ir��)�dg��	.�@�& G��R630���p v��p�&H�f��un���R57v�OJa�vG�`Y��owc��-ASF��O��7���SM������
af��rafLa�vl�\F c�w a���?VXpoV� �30��NT "L�FFM��=����yPh	a�G-�w�� �m2.�,�t��̹π6ԯ��sdF_�MC'V����D����fslm�is�c.  �H5522��21�&dc.pR7�8����0�708J614V�ip ATUtu�@�OL�545Ҵ�INTL�6�t8 ?(VCA����sseCRI���ȑ��UI���rt�\rL�28g��N�RE��.f,�63�!��,�SCH�d =Ek�DOCV���p���C,�<�L�0Q�i;sp��EIO��xEF,�54����9���2\sl,�SETp���lр�lt2��J7�ՌMA�SK��̀PR�XY҇��7���O[CO��J6l�3�<l�� (SVl�A��H�L�@Օ��539fRsv���#1���LCH���OPL]Gf�outl�0���D��HCR
sv�g��S@�h��CSa�!�{�50��D�l�q5!�lQ��DSW��aS����̀��OP����7��PR���L<�ұ�(Sgd���gPCM���R0 �\s��5P՝���0����n�q� AJ�1��N�q�2��PRS�a���69�� (A?uFRD�Խ���RMCN���9�3A�ɐCSN�BA�F9� HLB��� M��4���h��2A�95z�HTC�aԈ�TMIL6�j�95,��857.v,PA1�ito��oTPTXҴ JK�'TEL��piL��i XpL�80�I)��p.�!��P;�J95�ԏs "N���H�U{EC��7\cs��FR��<Q��C��5;7\{VCOa�,����IP1jH��S;UI�	CSX1�A�WEBa��HsTTa�8�R62���m`��GP%�IG� %tutKIPG�Sj�| RC1_m�e�H76��7�P�ws_+�?x�R;51�\iw�N�L��H�53!��wL�98!�h�R66��H����Ԡ���@;J56��1���N0��9�ej��L���R5`%��A|�5q�r�`,�8 5��{165!��@�"�5��H84!�29���0��PJ���n; B[�J77!ԨӃR6�5h3n���y36P��3R6��-`;о pԨ@��exeK�J87��#J90�!�stu+�~@!�۵�k90�koAp�B����@!�p�@|BA�g*�n@!��Q��#06!�@[�F�FaPb�6��́,�TS�w NC[�CAB$iiͰl1I��R7��p@q�y�CMS1�rog+QM�� �� sTY$x�CTOa�nv\+��1�(�,�6�con�~0�Ի15��JNN�%ep:��P��9ORS%tx���8A�815[�FCBaUnZQ�P!�p�p{��CMOB���"G��OL��x�O�PI�$\lr[�S�Š�T	D7�U��CP�RQR9RL���S��V�~`���K�ETS�$1��0���3\�Ԩ�FVR1�LZQ�V3D$ ���BV�a�SAPL1�CL�N[�PV��	rCC1Gaԙ��CL�3�CCRA�n "Wr!B�H�CSKQ�n\0�p��)�0CTPn�ЌQe��p.!$bCt�aT0U��pCTC�yЋRC�1�1 (�s��trsl,�r��
TX��;TCaerrm�r��MC"�s��#CT]E��nrr�REa��XPj�^��rmcH�^�a"�P�QF!$����$p "�rG,1�tTG$c8��Q�H�$SCTI�!� s��CTLqdACCK�Rp)��rLa�R82��M��YPk�.���OF��.���e��{�CN���^�1�"M�^�a�С�Q`US���!$��M�QW�$m�VGF�$R M�H��P2�� H5�� ΐq��ΐ�$(M-H[�VP�uoY���h�$)��D��hg���VPF��"MHG�̑`e!�+�V/vpcm�N��ՙ�N��$��VPRqd)��CV�x�V� "�X�,�1��($TIa�t\mh:��K��etpK��A%Y�VP%ɠ�!PN����GeneB�rip����8��extt���Y�m�"�(��HB� ��)��x��������Ȣ�res.�yA�ɠn����*���p�@M�_�N��6L���Ș�yAvL�Xr�Ȉ2��"R;�Ƚ\rax��	P�� h86���Gu+ʸ�Ͽ�Se0Lɨm�9�69�P����r�Ȩ2�ɹ1��n2��h� �0L�XR}�R�I{�e� L�x���c �Ș���N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1��/�k�@���A���ruk�ʘ L�scop��H�}�ts{������s��9��j7965��Sc��h���5 J9�{�
t�PL�J	een���t I[
x�comr��Fh�L�4 J���fo��DIF�+�6�Q����rat�i|��p��1�0�
R	8l߾�M�����PB��8� �j�mK�@X�HZ����N��oڠ��3�q��v�i���80�~�l� Sl�yQ��tpk�xb�j�.�@�R� d������,/n(�8�A8�0���
:�O8��<�Q}�CO���PT.��O (��.�Xp�|�~H���?�v� �wv��8�228�pm���722�j7�^�@ƙ���c�f�=Yvr���vcu���O�O�O�O�_#_5_7�3Y_��w3v4{_�_w�ʈ��ust_�_�cus�_�Z��oo,o>opPo�io��nge���(pLy747�jWe�lʨHM47ZKE�q {���[m�MFH�?�(wsK�8J��n���o��fh9l;��wmf���?� :�}(4	<g 9J{��II)̏މ9w��X�774kﭏ&/7ntˏ݊e+���3se�/�aw��8ͤɐ��EX \�!+: X�p��~�00��nh��,:Mo+�xO��1 �"K�O��\a��# 0��.8���{h�L?��j+�mon�:��tL�/�st�?-�w�: ���)�;��(=h��;
d Pۻ�{: 7 ��� �J0֛�re�����STD�!treLANG���81�\tqd����<���rch.��x����htwv��WWָ� R79��"Lo�51 (�I�W�h�Ո�4֧aww� �v�y �623c�h a?�cti�֘!�$X�iؠ�t �Ձn,�։����j<��"AJP@�3�p�vr{�H�6��!���- SeT� Ex3�) G�J934��{LoW�4 (S������� <���91 ��8!4�j9�所+�d��y�
��	�btN�ite{�R ��I@ Ո�����P��������	 ����Z�vol ��X ��9�<�I�p����ld*���F�86!4{��?��K�	��k扐�֘1�wmsk��M�q�Xa�Ae����p���0RBT�1ks.?OPTN�qf��U$ RTCam T��y��U��y�� U��UlU6L�T@�1Tx����SFq��Ue�6T��USP; W�b DT�qT2h�T�!/&+��8TX�U\j6&��U U�Usfd�O&�&ȁT���662DPN�abi��%�Q�%62V� �$���%�� �#(�(6{To6e St�%���#5y�$�)5(To�%tT0�%5�W6�T���%�#�#orc���#I���#���%c�ct�6ؑ?�4\W6965"p6}"�#\j536���4�"��?kruO O,Im ?Np�C �?t�0<O�;�e �%���?�
;gcJ7 "AV<�?�;avsf�O__&_8WtpD_V_0GT�F|_:UcK6�_�_9r�O�3e\s�O2^�y`O:�migxGvNgW! m�%��!�%T�$E A{6�po6̀�#37N�)5R5�_2E���$0���$Ada�Vd���V�?;Tpz7�_�e7DDTF9���#8�`�%��4~y�ted Z@0�A}�@�}�04N�}�0}���}�dc& }����u 6�v��v1�u1\b�u$2}�<��}� R83�u�"x}��"}�valg���Nrh�&�8�J��Y�o�ue��� j7q0�v=1��MIG�uerfa��{q����E�N�ء��EYE�ce A���� �pV�e�A!���2Յ�Q �%��u1�e�i�@��@H�e����J0� '��b��T��E In��B�  W�|��5�37g����(MI�t�Ԇr��ݟ�Cam���nеv!g�U -�v J߆8⹖0F���P�y�ac���28���Rɏ jo��2�� djd�8r}�� og\k�0��gܕ�wmf�Fro/� Eq'�4"}��3 J8��oni[��ᅩ}Ĵ��C o� ��ʛ��m@�R�e��{n�Д�V��o������  �����裆"P�OS\����ͯ mcenϖ�⑥OMo��43��� �(Coc� An[�t���"Fe�a\�vp��.��ocflx$�le��`8�hr�tr�NT�w CF+�x E/�at	qi�M�ӓxc�֌p�f�lx����Z�c�x��
0 h��h8f��mo��=� H����)� (�vSER�,���g�0߆0\�r�vX�= ��I � - �ti��H���VC�828�5ص�L"�RC��n �G/���w�P�y�\v�vm "o�lϚ��x`��=e�ߠ-�R-3?������vM [��AX/2�)�S�r�xl�v#�0��h8�߷=� RAX�AТ����9�H�E/�Rצ����h߶"R�Xk��F�˦85ή�2L/�xB88�5_�q�Ro�0iA��5\rO�9�K��v����8���.�gn "�v��88��8s�i ?�9 �����/�$�y O�MS"����&�9R H784&�`�745�	pp��p��ycr0C�Rc�hP0� j�-�a�%?o��6D950R7tsrl��ctlO��APC���j�ui�"�L���  ����K^棆!�A��qH���&-^7����� ��616C�q�794h����� M�ƔI��99���(��$F�EAT_ADD �?	���Q~%P  	�H ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n���������TDEMO �fY   WM_��� �����//%/ R/I/[/�//�/�/�/ �/�/�/�/?!?N?E? W?�?{?�?�?�?�?�? �?�?OOJOAOSO�O wO�O�O�O�O�O�O�O __F_=_O_|_s_�_ �_�_�_�_�_�_oo Bo9oKoxooo�o�o�o �o�o�o�o>5 Gtk}���� ����:�1�C�p� g�y�������܏ӏ� ��	�6�-�?�l�c�u� ������؟ϟ���� 2�)�;�h�_�q����� ��ԯ˯ݯ���.�%� 7�d�[�m�������п ǿٿ���*�!�3�`� W�iϖύϟ������� ����&��/�\�S�e� �߉ߛ��߿������� "��+�X�O�a��� ������������� '�T�K�]��������� ��������#P GY�}���� ��LCU �y������ /	//H/?/Q/~/u/ �/�/�/�/�/�/?? ?D?;?M?z?q?�?�? �?�?�?�?
OOO@O 7OIOvOmOO�O�O�O �O�O_�O_<_3_E_ r_i_{_�_�_�_�_�_ o�_o8o/oAonoeo wo�o�o�o�o�o�o�o 4+=jas� �������0� '�9�f�]�o������� ��ɏ�����,�#�5� b�Y�k���������ş ����(��1�^�U� g������������� ��$��-�Z�Q�c��� ����������� � �)�V�M�_όσϕ� �Ϲ���������%� R�I�[߈�ߑ߫ߵ� ��������!�N�E� W��{�������� �����J�A�S��� w������������� F=O|s� ����� B9Kxo��� ���/�/>/5/ G/t/k/}/�/�/�/�/ �/?�/?:?1?C?p? g?y?�?�?�?�?�? O �?	O6O-O?OlOcOuO �O�O�O�O�O�O�O_ 2_)_;_h___q_�_�_ �_�_�_�_�_o.o%o 7odo[omo�o�o�o�o �o�o�o�o*!3` Wi������ ��&��/�\�S�e� ������������� "��+�X�O�a�{��� �������ߟ��� '�T�K�]�w������� ���ۯ���#�P� G�Y�s�}�������� ׿����L�C�U� o�yϦϝϯ������� �	��H�?�Q�k�u� �ߙ߫��������� �D�;�M�g�q��� ��������
���@� 7�I�c�m��������� ������<3E _i������ �8/A[e �������� /4/+/=/W/a/�/�/ �/�/�/�/�/�/?0? '?9?S?]?�?�?�?�? �?�?�?�?�?,O#O5O OOYO�O}O�O�O�O�O �O�O�O(__1_K_U_ �_y_�_�_�_�_�_�_ �_$oo-oGoQo~ouo �o�o�o�o�o�o�o  )CMzq�� �������%� ?�I�v�m����������ُ���;�  2�Q�c�u��� ������ϟ���� )�;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����� ��1CUg y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����'>9  :> Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{��������/=C6Yk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A���$FEAT_D�EMOIN  VE��q��>�Y�_INDEXf�u���Y�ILECOM�P g������t�T���S�ETUP2 h������  �N ܑ��_AP2�BCK 1i��  �)B���%�C�>���1�n� E����)���M�˯�� �����<�N�ݯr�� ����7�̿[��ϑ� &ϵ�J�ٿWπ�Ϥ� 3�����i��ύ�"�4� ��X���|ߎ�߲�A� ��e�����0��T� f��ߊ�����O��� s�����>���b��� o���'���K������� ��:L��p��� �5�Y�}�$ �H�l~�1 ��g�� /2/� V/�z/	/�/�/?/�/ c/�/
?�/.?�/R?d? �/�??�?�?M?�?q?@O�?O<O���P�� 2�*.V1RCO�O�0*�O�O`�3�O�O�5w@PC�O|_�0FR6:�O"=^�Oa_�KT���_ �_&U�_�\h�R_�_�6�*.FzOo�1	�(SoEl�_io�[STM �b�o�^+P�o��m�0iPen�dant Panel�o�[H�o �g��oYor�ZGIF |��e�Oa��ZJPG �*��e���z��JJS�����0�@���X�%
Ja�vaScriptُ�CSʏ1��f��ۏ %Casc�ading St�yle Shee�ts]��0
ARGNAME.DT��
�<�`\��^���Д�៍�АDISP*ן���`$�d��V��e��CLLB.cZI��=�/`:\���\�����Col�labo鯕�	P�ANEL1[�C�%��`,�l��o�o�2 a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V���zό��!ߘ�TPEINS�.XML(�@�:\�<����Custo�m Toolba�r}��PASSW�ORD���>FR�S:\��� %�Password Config� �?J���C��"O��3� ����i����"�4��� X���|�����A��� e�����0��Tf �����O�s ��>�b�[ �'�K���/ �:/L/�p/��/#/ 5/�/Y/�/}/�/$?�/ H?�/l?~??�?1?�? �?g?�?�? O�?�?VO �?zO	OsO�O?O�OcO �O
_�O._�OR_d_�O �__�_;_M_�_q_o �_�_<o�_`o�_�o�o %o�oIo�o�oo�o 8�o�on�o�!� �W�{�"��F� �j�|����/�ďS� e���������T�� x������=�ҟa��� ���,���P�ߟ񟆯 ���9����o���� (�:�ɯ^�����#� ��G�ܿk�}�ϡ�6� ſ/�l�����ϴ��� U���y�� ߯�D��� h���	ߞ�-���Q߻���߇��,��$FI�LE_DGBCK� 1i������ (� �)
SUMM?ARY.DG,���OMD:`�����Diag Su�mmary���
CONSLOG���y����$���Co�nsole lo�g%���	TPACCN��%g������TP Acco�untinF����FR6:IPKD?MP.ZIP�����
��)����Exc?eption-�����MEMCHEC�K�����8�M�emory Da�ta��LN�=)�RIPE����0�%� �Packet L�E���$Sn�S�TAT*#�� %LSta�tus�i	FTAP�/�/�:��mment TB�D=/� >)ETHERNE��/o�/�/��Et�hernU<�fi�guraL��'!DCSVRF1//)/�B?�0 verify allE?��M(5DIFF:? ?2?�?F\8diff�?}7o0CHGD1�?�?�?�LO �?sO~3&��
I2BO)O;O�O� bO�O�OGD3p�O�O�OT_ �O�{_
VUPDAT�ES.�P�_��FORS:\�_�]���Updates �List�_��PS�RBWLD.CM�o���Ro�_9�P�S_ROBOWEyL^/�/:GIG��o>_�o�Gig�E ��nosti�cW�N�>�)}�aHADOW�o�o�ob�Sha�dow Chan�ge��8+"rNOTI?=O���Notif�ic�"��O�A=�PMIO�o���h��f/��o�^U�*�UI3�E�W��&{�UI������B� ��f��_�������O� ��������>�P�ߟ t������9�ί]�� ���(���L�ۯp��� ���5�ʿܿk� Ϗ� $�6�ſZ��~��w� ��C���g���ߝ�2� ��V�h��ό�߰��� Q���u�
���@��� d��߈��)��M��� ������<�N���r� ���%�����[���� &��J��n� �3��i��" �X�|�� A�e�/�0/� T/f/��//�/=/�/��/�$�$FILE�_�PPR�P���� �����(MDONLY� 1i5�  
 �z/Q?�/u?�/ �?�?t/�?^?�?O�? )O�?MO_O�?�OO�O �OHO�OlO_�O_7_ �O[_�O_�_ _�_D_ �_�_z_o�_3oEo�_ io�_�oo�o�oRo�o vo�oA�oew �*��`�����&�O��*VIS�BCK,81;3*�.VDV����F�R:\o�ION\�DATA\��/���Vision� VD file ̏��&�<�J�4�n� �����3�ȟW���� ��"���F�՟�|�� ����m�֯e������ 0���T��x������ =�ҿa�s�ϗ�,�>� ��b���ϗϼ�K� ��o��ߥ�:���^�����ϔ��*MR2_�GRP 1j;��C4  B�}�	 71�������E�� E�  �F@ F�5U�������L����M��Jk��Lzp�JP���Fg�f�?� � S����9�Y�9}�9���8j
�6���6�;��A� � ���BH��B���B���$�������������@UUU#�����Y�D�}� h����������������
C��_CFG� k;T �M���]�NO {:
F0�� � \�RM_CHKTYP  0��}�000��O=M_MIN	x�g��50X� �SSBdl5:0��bx�Y����%TP_DEF'_OW0x�9��IRCOM���$GENOVRD�_DO*62�T[HR* d%d�o_ENB� �/RAVC��mK�� ��՚�/3�/���/�/�� ��M!OUW s���}��ؾ��8��g�;?�/7?Y?[? 7 C��0����(7l�?�<B�?B�����2��*9�N SMT�T#t[)��X�4�$�HOSTCd1u�x���?�� kMCx��;zO�x�  27.0z�@1�O  e�O �O	__-_;Z�O^_p_��_�_�LN_HS	anonymous�_ �_�_oo1o yO��FhFk�O�_�o�O�o �o�o�oJ_'9K ]�o�_���� �4o�XojoG�~�o ^�������ŏ��� ��1�T���y��� ��������,�>�@� -�t�Q�c�u������� ��ϯ���(�^�� M�_�q�����ܟ� � ݿ��H�%�7�I�[� ��ϑϣϵ����l� 2��!�3�E�Wߞ��� ¿Կ����
������ �/�v�S�e�w��� �����������+� r߄ߖ�s�����߻� ���������'9K ]�������� �4�F�X�j�l>�� }������ //1/T��y/�/��/�/�/.D\AENT� 1v
; P!\J/?  ��/ 3?"?W??{?>?�?b? �?�?�?�?�?O�?AO OeO(O�OLO^O�O�O �O�O_�O+_�O _a_ $_�_H_�_l_�_�_�_ o�_'o�_Koooo2o {oVo�o�o�o�o�o �o5�oY.�R�v��zQUICC0���3��tA14��"����t2���`�r�ӏ!ROU�TERԏ��#�!?PCJOG$����!192.168.0.10�~�sCAMPRTt�P�!d�1m������RT폟�����$N�AME !�*!�ROBO���S_CFG 1u�)� �A�uto-star�tedFTP&��=?/֯s�� ��0�B��f�x��� ������S������ ,���������ϼ�ޯ ���������ʿ'�9� K�]�oߒ�ߥ߷��� ������(:~� k�Ϗ�������� ����1�C�f���y� �����������,�>� R�?��cu�� `�����(� $M_q������  /H%/7/I/ [/m/4�/�/�/�/�/ �~/?!?3?E?W?i? ����?�/�?/�? OO/O�/�?eOwO�O �O�?�ORO�O�O__ +_r?�?�?�?�O|_�? �_�_�_�_o�O'o9o Ko]ooo�_o�o�o�o �o�o�oF_X_j_~o k�_������o ���1�TU��y����������U�)�_ERR w3�я��PDUSIZ  �g�^�p���>~�WRD ?r��Cq�  guestb�Q�c��u�������"�SCD�MNGRP 2x�r�����Cqg�\�b�K� 	�P01.00 �8(q   ��5p�5pz�5pB�  �{ ���H���L���L��L������O8�����l�����Ua4� x��Ȥ�x���8���\���)j�`�;�������d�.�@�R�ɛ__GROUېy�����	ӑ���QUPD  ?u�����İTYg�����TTP_A�UTH 1z��� <!iPen'dan��-�l����!KAREL�:*-�6�H�KC�]�m��U�VISION SET�� �ϴ�g�G�U������ R�0��H�Bߏ�f�x���ߜ߮���CTRL� {����g�
�S�FFF9E�3��AtFRS:DEFAULT;��FANUC �Web Server;�)����9�K� �ܭ���������߄�WR_CONFI�G |ߛ �;��IDL_CP�U_PCZ�g�B��Dpy� BH_�M�INj�)�}�GNR_IO��g���a��NPT_SIM_�D_�����STA�L_SCRN�� ����TPMODN�TOL������RT�Y��y���� �EN�O���Ѳ]�OLN/K 1}��M���������eM�ASTE��ɾeSLAVE ~��|c�O_CFG�ٱBUO�O@C�YCLEn>T�_?ASG 1ߗ+�
 ����/ /+/=/O/a/s/�/�/p�/�/��NUM���
@IPCH��^RTRY_CNZ���@��������� @kI��+E�z?E�a�P_�MEMBERS �2�ߙ� $���2���ݰ7�?�9a��SDT_ISOL�C  ����$�J23_DSM�+�3JOBPRO�CN��JOG��1�+�d8��?��+�O�/?
�LQ�O__/_@�OS_e_w_�_`�O� Hm@��E#?&BPO�SREQO��KANJI_���a[�?MON ����b�yN_goyo�o�o�oH�Y�`3�<� ��e�_ִ��_L���"?�`EYLOGGI�NLE��������$LANGUA�GE ��<�T� {q�LGa2��	�b���g�xP��W  ��g��'��b���>��MC:\RSCH�\00\<�XpN_DISP �+�G�J��O�O߃LOClp�Dz���As�OGBOOK ������󑧱����X�����Ϗ�����a�*��	 p�����!�m��!����=p_BUFF 1-�p��2F幟����՟D� Co�llaborativǖ���F�=�O� a�s�������֯ͯ߯����B�9�K���D�CS �z� =���'�f��?ɿۿ����H@{�IO 1�� ~?9ü��9�I�[�mρϑϣ� �����������!�3� E�Y�i�{ߍߡ߱���h�����E��TMNd�_B�T�f�x��� ������������,� >�P�b�t�������L�N�SEVD0��TYPN1�$6���QRS"0&��><2FL 1�"�J0��������GTP:pO}F�NGNAM1D��mr�tUPS�G�I"5�aO5�_L�OADN@G %��%TI�pZU�ZAUN#�(MA?XUALRM�'��8�(��_PR"4F0�d��1�B_PN�P� V 2�C�	MDR077�1ߕ�BL"80{63%�@ �_#�?�ߒ|/�C���z�6��/���/Po@Pw 2��+ �ɖ�	T 	t  ��/�%W?B?{? �k?�?g?�?�?�?O �?*OONO`OCO�OoO �O�O�O�O�O_�O&_ 8__\_G_�_�_u_�_ �_�_�_�_o�_4oo XojoMo�oyo�o�o�o �o�o�o0B%f Q�u����� ���>�)�b�M��� ��{��������Տ� �:�%�^�p�S��������D_LDXD�ISApB�ME�MO_APjE {?C
 �, �(�:�L�^�p�������� 1�C ����4��������4��X���C_MS�TR ���w�S_CD 1���L� ƿH��տ���2�� /�h�Sό�wϰϛ��� ����
���.��R�=� v�aߚ߅ߗ��߻��� ����<�'�L�r�]� ������������ ��8�#�\�G���k��� ������������" F1jUg��� ����B- fQ�u���h��MKCFG �����/�#LTARMU_��7"0��0N/V$� MET�PUᐒ3����N}D� ADCOLp%�� {.CMNT�/ 9�%� ����.�E#>!�/4�%POS�CF�'�.PRP�M�/9ST� 1�޿� 4@��<#�
1�5�?�7{? �?�?�?�?�?�?)OO O_OAOSO�OwO�O�O�O�O_�A�!SIN�G_CHK  ~�/$MODAQ,#����.;UDEV� 	��	MC}:o\HSIZE�����;UTASK �%��%$123456789 �_��U9WTRIG 1���l3%%��9o��`"ocoFo5#�VYP�Q�Ne��:SEM_I�NF 1�3'� `)AT&FV0E0po��m)�aE0V1�&A3&B1&D�2&S0&C1S�0=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o '��K������ �я:�L�3�p�#�5� ��Y�k�}������$� [�H���~�9����� Ưد��������ӟ� V�	�z�������c�Կ ����
��.���d� �)�;��Ͼ�q���� ���˿<���`�G߄� ��IϺ�m�ϑϣ�� ��8�J��n�!ߒ�M��������h_NIT�OR� G ?�[ �  	EXESC1�/�25�35�E45�55��P7�75�85�9�0�Қ� 4��@��L��X�� d��p��|����T���2��2��2��U2��2��2��2��U2��223���3��3@�;QR_G�RP_SV 1��k (�A�z��4�~�K��������K:z3�j]�Q_D��^��PL_NAME� !3%,�!�Default� Persona�lity (from FD) ��RR2� 1�L6(L?�,0	l d��� �����//(/ :/L/^/p/�/�/�/�/�/�/�/ZX2u?0? B?T?f?x?�?�?�?�?\R<?�?�?O O2O DOVOhOzO�O�O�OZZ�`\R�?�N
�O_\TP�O:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHo_)_~o �o�o�o�o�o�o�o  2DVhz�[o mo����
��.� @�R�d�v����������Џ� Ef � Fb� F7�<��   ��!��d��@�R�6�t� �����l���ʝ����� ݘ��� �"�@�F�d���� "������ݐA�  HϩU[�$n�B�E ��� � @D� M �?�� �?�@<��A@�;f��F�H� ;�	l,�	O |��j�s�^d�>��� ���� K(��Kd$�2K ��J7w��KYJ˷�ϜJ�	�ܿ�� �@I���_f��@�z��f�|��γ�N�������	Xl��������S�Ľ�����I ����~5���  �����A?oi#�;����� ���l� �Ϫ�-���PܛG�G�Ѳ��@�n�@a   ?�  ��ܟ�*�͵	'� �� H�I� ��  �Рn�:��Èl�È=��9̈́�в@�ߚ� �����/������̷NP�  '�,���-�@
�@W���?=�@A����B�  C�j�a�Be�Ci��#��Bи�E F� ,ee��^^ȹBР��P�����̠�����ADz ՟�n�3��C�i�@��R�R�Y����  ��@� ���  <���?�ff������n� ɠ#ѱ@y9G
(���I�(�@uP~����t�t����>����;�Cd;���.<߈<��g�<F+<AL�������,�d�|,�̠?fff?���?&&��@���@x��@�N��@���@T� H�ِ�!-�ȹ�| ��
`������ �//</'/`/r/]/�/��eF���/�/ �/�/m?��/J?�(�E��G�#�� FY�T?�?P?�?�? �?�?�?O�?/OO?O eOk��O�IQOG�? �O1?�OmO_0_B_T_"������A_�_@	_�_�_�_ o��A��aAn0 bФ/o C�_pUo�_�Op��؃o��o�o�o���W������oC�E�  q�H�d��؜a@q���e�F�BµWB�]�NB2�(A���@�u\?��D�������b��0�|�uR�Ｃ�
x~������Bu*�C��$�)`��$ ���GC�#���rA�U����1��eG�D�I�m�H�� I:��I�6[F����C�I��J��:\IT�H
~QF�y���p�*J�/ �I8Y�I��KFjʻCe�o�� s�����Џ���ߏ� *��N�9�r�]����� �������۟���8� #�\�G�����}����� گů���"���X� C�|�g�����Ŀ��� ����	�B�-�f�Q� ��uχ��ϫ������ ��,��P�b�M߆�q� �ߕ��߹�������(� �L�7�p�[����������s($���33:����$���3���d�,�4���@�R�wa����l�~�wa���ex����wa4 �{�� ����(L:ue%P�P~�A�O�������	����G2W} h������/����O�O7/m/[(d =�s/U/�/�/�/�/�/ ?�/1??U?C?y?�=  2 Ef9g�Fb��77�9fBX)aa)`C9A`�&`w`@-o�?w`e�O)O�?MO�Ow`�?�?�O�O�O�O9c?�0�A7h�t4w`w`!:w`xn
 �O9_ K_]_o_�_�_�_�_�_��_�_�_o#ozzQ ���h��G����$MR_CABL�E 2�h ��a�T� @�@�0�Ae��a�a�a�%�`��0�`C�`�a�O8�tB�nׇd��`�aE�4�E�#�o�f-�#��0��0�D�O��By`���Š��bED4E�c,��o�go8  ���C�0�7�d4
vے��0 �b��XE'�Z&�l�`y`r
qC�p�bHE�
v�#g�5D�Ү(�qz�lҠ`��0�q��p�b0�
v�%�c���b=%	E;h��u/o�c-��4 tH�\�?�9�K�]�o� ԏϏ��
�ɏۏ@���?��e o<�\����������������*,�** \cO�M �ii���3Jq { %�% 234567O8901i�{� f�H����������1�����
��`��not sent� 5���;��TESTFECSALGR  e�q�iG�1d.�š
:�� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.x�ml��ֿqY��DEFAULT�-�i4\bGRP 2�M�  =��a�7��E  �%Fo�rce�sor check  ��
�b�z��p����h5-��ϻ���������%!1st cl�eaning o�f cont. �v�ilatio!n��}�Rߗ+��[��ߔߦ߸���mwech�cal`������0��h5k�@�R�d�v��|��(�rolle_������/����(�:�L��Bas�ic quarterly�������,�����������#M��:C@"GpP�a�b`i4�������#C���M"��{Pbt�|��Suppq�?grease���?/&/8/J/�\/��C+ ge��./ batn�y`/��/h5	/�/�/�/?� ?_�ѷen'�v��/�/��/��?�?0�?�?�?�G=?O��qp"CrB1O��0 �/`OrO�O�O�O�t$,��Lf��C-ݐ�A�O:�OO$_6_H_Z_�l_�t*cabl,�Oݒ��S<ݐ�Q�_:�
_�_�_oo�0oo)(Ӂ/�_�_����_�o�o�o�o�o��O@hau1�l�2r xݐ<qC:��op������_ReplaW�fU��2�:�._4�F�X�j�|�ݐ$%���ߟ ����#���
��.�@� ��d���ŏ׏����П ����U�*�y����� r���������	�q�� ?�߯c�8�J�\�n��� ϯ�����ڿ)���� "�4�Fϕ�jϹ�˿�� ����������[�0� ϑ�fߵϊߜ߮��� ��!���E�W�,�{�P� b�t����߼��� ��A��(�:�L�^��� ������������  $s�H������q �����9] o�Vhz��� U�#�G/./@/ R/d/��/�/��// �/�/??*?y/N?�/ �/�?�/�?�?�?�?�? ??Oc?u?JO�?nO�O��O�O�O+J1B	 H �O�O__6M2_@OBE :_p_>_P_�_�_�_�_ �_ o�_�_oHoo(o Zo�o^opo�o�o�o�o��o �o :z ̾bA?�  @!Q _���Fwp�� �H* �** @q>v�p2T��f�x�:�������ҏ��eO^C7�Տ#�5� G�	�k�}���ُ��� c�����W��C�U� g���ß)�����ӯ� ��	��-�w�����9� ������m�Ͽ��=��O�E!Q�$MR�_HIST 2��>uN�� 
 \�
B$ 2345678901^�f�#�
�]�9O���φ� ��O�)�;����q� �ߕ�L�^߬����ߦ� ���7�I� �m�$�� ��Z���~������!� ��E�W��{�2������h�����:�SKCF�MAP  >uKQ��r5�!P�����ONREL7  .�3����EXCFENB�8
��QFNC�XJJOGOVL�IM8dNá ��K�EY8��_�PAN7����R�UN����SFSPDTYPx<C��SIGN8J�T1MOT�G���_CE_GRP7 1�>uV� �@�����/Ⱥ ��/�/U//y/ 0/n/�/f/�/�/�/	? �/???�/c??\?�? P?�?�?�?�?�?O)O�OMO,���QZ_E�DIT5 )TC�OM_CFG 1����[�O�O�O }
�ASI �yB3�
__+[_�O_��>O�_bHT__ARC_U.���	T_MN_MO�DE5�	UA�P_CPL�_gN�OCHECK ?��� ��  o.o@oRodovo�o�o �o�o�o�o�o*�!NO_WAITc_L4~GiNT�A����EUwT_E�RRs2���3��@ƱJ�����>_�)��|MO�s��}x�:Ov���8�?������ l��rP�ARAM�r�����j���5�5�G� = ��d�v�~� X������������֟0�0����b�t������SUM_RSPACE�����Aѯ�ۤ�$ODRDS�P�S7cOFFS?ET_CARt@�_��DIS��PE?N_FILE:�7��AF�PTION�_IO��q�M_�PRG %��%�$*����M�WOR�K �yf ���춍��� ������	 �������gT��R�G_DSBL  ���C�{u��R�IENTTO7 f�C� A ��UT_SIM_D�y���V�LCT ��}{B �<٭��_PEX�P=�n�RAT�W dc���UP ���`���e�w�]߬�ߩ��$�2r��L6(L?�>��	l d���� ��&�8�J�\�n�� ������������� "�4�F�X���2�߈� ������������*�<w�Tfx� ������J`[ˣG���Tz��Pg�� ����/"/4/F/ X/j/|/�/�/�/�� �/�/??0?B?T?f? x?�?�?�?�?�?�?�? �/�/,O>OPObOtO�O �O�O�O�O�O�O__`(_:_��O��y_�]2ӆ��_�^�_�_ �W^]^]��/ooSog�Hgrohozo�o�o �o�o�oF`�#|`�A�  9y�����OK�1�k������<o�EA�nq? @D�  �q��4��nq?��C��s�q|1� ;�	l���	 |�Q�s��r�q>��u ��sF`H<zH~��H3k7GL��zHpG��99l7�k_B�T�F`SC4��k�H���t���-�Ae���k������s��� � �ሏ����EeBVT���dZ=����ڏ ���q-�Fk�y�{jFbU�= n@}6�  ����z�Fo��Be	'�� � ��I� �  �:p܋=���ڟ웆�@���B�,�D��B���g�AgN����  '|���g���B��p�BӀC�׏����@  #��Bu�&�ee^�^^މB:p 2���>�m�6p�Z�=Dz?o}�܏�������׿������Ǒ��� ~f�  � �M�z��*�?�ff�_8�J�ܿ 3pϑ�ñ8= �ϵʖq.·�	(= ��P���'��s��tL�>��/�;�C�d;��.<���<�g�<F+<L ��^oiΚr�d@��r6p?fff�?�?&�п�@���@x��@��N�@���@T싶�Z���ћtމ �u�߈w	�x��ti�>� )�b�M��q����� ��������:�%�^��������W���S�E��  G�=F�� Fk��������� 1U@yd�� ����q��	�� {�A��h����D�a��ird��A{�/w/J/5/n/	�A�A���":t�/ C�^/�/Z/ ލ?����/�/1??���Wҵ���g��pE�! ~1�?04�0
1ή1@IӀ��B���WB]�NB2��(A��@��u\?��������������b�0�|�uR����
�>��ؽ��B�u*C��$��)`�? ����GC#����rAU�����1�eG���I��mH�� I�:�I�6[Fߍ��C4OI���J�:\IT��H
~QF��y�Ol@�*J��/ I8Y�I���KFjʻC ��-?�O�O__>_)_ b_M_�_�_�_�_�_�_ �_o�_(oo%o^oIo �omo�o�o�o�o�o  �o$H3lW� {������� 2��V�h�S���w��� ��ԏ�������.�� R�=�v�a�������П ����ߟ��<�'�`� K�]���������ޯɯ���&�8�#�\��3(�J���3:a���9���J�3��c4�����������������ڿ�n�����e��n�4 �{2�2�r�`ϖτ�(�Ϩ��%PR�P���!�h�!�K�6�o�Z�����u�|ߵ� �����������3�� W�B�{�f�4���������d�A����!�� 1�3�E�{�i��������������  2 �Ef�7Fb�7���6B�!�!� C9� �� n�@�/`r@������#x�@�+=�3?, TV�8v�n�n���n��.
  D�����// %/7/I/[/m//�/�:� ��ֻ�G����$PARAM�_MENU ?�2�� � DEFP�ULSE�+	W�AITTMOUT��+RCV? �SHELL_W�RK.$CUR_oSTYL� 4<�OPTJJ?PTB�_?Y2C/?R_DECSN 0�Ű<�?�? �?�?�?OO?O:OLO�^O�O�O�O�O�O�!S�SREL_ID � .����EUS�E_PROG �%�*%�O0_�CCC�R0�B��#CW_H�OST !�*!HT�_=ZT��O_�S�h_zQ�S�_<[_TGIME
2�FXU� ?GDEBUG�@�+��CGINP_FLgMSKo5iTRDo�5gPGAb` %l��tkCHCo4hTY+PE�,� �O�O �o#0Bkfx �������� �C�>�P�b������� ��ӏΏ�����(��:�c�^�p�����7eW�ORD ?	�+
? 	RSc`n�/PNS��C4�sJOv1��TE�P�COL�է�2�Z�gLP 3��n���OjTRACEC�TL 1�2���! �� ��Қ�q�DT� Q�2�Ǡ��D � :����Ԡ�Ԡ��}�ׯ���;�4��4� �4���;�u:�q:�T��;�8�	8�
8�U8�8�8�8�Q8��@:�8�8����� ���ٱ
޴���ؿ�$� 6���
�l�~�@�R�d� �ϰ���������
�� V�h�zߌߞ߰����� ����
�,�>�P�*�<�v��*� +8�+ (��)��*���� ������)�;�M�_� q��������������� %,�>�P�b�t� �����������С� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 @ubt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀�V�߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�?�?�?�?�1�$PG�TRACELEN�  �1  �_��0��6�_UP �����A@�1�@�1_CFG M�E�3�1
@�<D�0<DZO<C��0uO$BDEFSP/D �/L�1�0���0H_CON?FIG �E�3W �0�0d�DM��2 �1�APpD�sA�A�0��0IN~'@TRL �/M�OA8pEQPE�E��G�A<D�A�ILID(C�/M	~bTGRP 1ýI� l�1B�  �����1A��33FC� F�8� E�� @eN	�A�AsA�Y�Y�A�@� 	RO�Hg��_ ´8cokB ;`baBo,o>oxobo�o��1>о�?B�/�o�o~�o =?%<��
C @yd��"�������  Dz@�I�@A0�q� ��� ����ˏ���ڏ��� 7�"�4�m�X���|����Ú)ґ
V7.10beta1HF @�����Aq��Q m �?� �BܠPz�p �C��&�?B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@��8�f������ҡ�R9�ܣ�Rљ���1��i�������t<B!CeQKNOW_M  lE7FbT�SV ĽJ �BoC_�b�t�������@������1�]aSM�S]ŽK ���	NB~�0���Ŀ�K���-�bb ��A�RP����0��Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1�K
 4MU�iǨj� K�]�oߠߓ� �߷�������2��#� h�G�Y��}�����@��
������,�27�9I��1�<t�H���P3^�p�����,�4 ��������,�5(:,�6Wi{��,�7����,�8��!3,�MAD��6 F,�OVL/D  KD�xO�.�PARNUM � �MC/%�SCH� E
9'!G)�3Y%UPD/��E|�/P�_CMP_���0@�0'7E�$E_R_CHK�%5H�&�/�+RS���bQG_MO�+?=5_'?~O�_RES_G6��:�I�o�?�?�?�? O�?O7O*O[ONOO�rO�O�O�{4]��< �?�Oz5���O__|3  #_B_G_|3V b_�_ �_|3� �_�_�_|3�  �_�_o|3Oo>oCo|2V 1�:�k1!��@c?�=2THR_INRc0i!}�zo5d�fMASS�o� Z�gMN�o�cM�ON_QUEUE� �:�"�j0��*O�N� U1Nv�+�DpENDFqd?`yEcXEo`u� BEnp|PAsOPTIOMw�m;DpPROGRAoM %$z%Cp�}o(/BrTASK_�I��~OCFG ��$��K�DAkTA��T���j12/ď֏���� ��+�=�O�a������𩟻�͟��INFO
�͘��3t��!�3� E�W�i�{�������ï կ�����/�A�S��e�w�����Θ� �'��FJ�a K_N�q�T��˶ENBg Hڽw1��2��GN��2�ڻ P(�O�=���]ϸ��@���v� ��u�uɡdƷ_EDIT �T�����>G�WERFL�x�c�)�RGADJ �Ҷ�A�  $�?@j00��a�Dqձӆ5�?�����<u�)%e���Ș��FӨ�2�R��	�H;pl�G�b_�>��pAod�t$��*�/� **�:�j0�$�@�5 Y�T���^��q�߈b ~�L��\�n���� �����������4� F�t�j�|��������� ����bLBT �x����:� �$,�Pb� ��/����/ ~/(/:/h/^/p/�/�/ �/�/�/�/V? ??@? 6?H?�?l?~?�?�?�? .O�?�?OO O�ODO VO�OzO�O_�O�O�O �O�Or__._\_R_d_��_�_�_�_�_�_�f	 g�io�pWo�o{d�o��~o�ozoB�P?REF �Rږp��p
�IORI�TY�w[���MP�DSP�q��pwUT�6����ODUCT�3�����OG��_TG��8�����rTOENT 1�׶� (!AF_INE�p,�7�?!tcp7�_��!udN���!icmv��ޯrkXYK�ض���q�)� ,�����p��&�	��R�9�v� ]�o�����П����� �*��N�`�*�sK���9}�ߢ���Ư �,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE� �R��:�wd��连�2s�9Ks���PORT_NUUM�s�p����_CARTREP�{p�Ω�SKSTAv�w d�LGS)��ݶ��tӁpU�nothing��������{��TEMP ޾y��'e���_a_seiban�o\��olߒ� }߶ߡ���������"� ��X�C�|�g��� ����������	�B� -�f�Q���u������� ������,<b M�q��������(L�VE�RSIyp�w} �disabl�edWSAVE �߾z	260_0H768S?��!ؿ����/ !	5(�r)og+^/yÁe{/�/�/�/�/�*��,/? �p���_��p 1�Ћ�? �����Wh?xz?�W*pURGE��aB�p}vgu,�WF�0#DO�vƲ�vW%��4�(�C�WRUP_DELAY �\���5R_HOT �%Nf�q׿GO�5R_?NORMAL&H�rx6O�OZGSEMIjO��O�O(qQSKIPF3��W3x=_9 8_J_\_]�_�_{_�_ �_�_�_�_�_	o/oAo Soowoeo�o�o�o�o �o�o�o+=a Oq������ ��'��7�]�K���x����)E�$RA{����K/�zĀÁ_�PARAM�A3���K @.�@`\�61�2C<��y�M�C�6$�BÀ�BTIF�4`�RC_VTMOUu�cŻ�ÀDCRF3��I �+Q;�/�CC�SeD��#�1=h��-0�t]�/��ޅ�����1��0��_��k_����Cd;��.<�߈<�g�<?F+<L���Ѱ��d�u�L������� ϯ����)�;�M��_���RDIO_T?YPE  M=U��k�EFPOS1 ;1�\�
 x4/�����+�$/<�� $υ�pϩ�D���h��� ���'������o�
� ��.ߤ�Rߌ������ ��5���Y���i��*� <�v���r������� ��U�@�y����8��� \�����������?��xc����2 1�KԿX�T�x��3 1�����nY�S4 1�'9K�/�|'/�S5 1����/�/�/�/:/S6 1�Q/c/u/�/�-??Q?�/S7 1��/�/
?D?�?�?�?>d?S8 1�{?�?��?�?WOBO{O�?SM?ASK 1L�8�O�D�GXNO���Fx&�^��MOTEZ�hŻ��Q_ǁ�%]�pA݂��PL_RA�NG!Q]�_QOWE/R �ŵ�P1V�SM_DRYPR/G %ź%"O�_��UTART ���^�ZUME_PR�O�_�_4o��_EX�EC_ENB  yJ�e�GSPD`pO`WhՅjbTDBro�jRM�o�hING�VERSION �Ź#o�)I_AIRPURhP� �O(�MMT_ҡ@T�P#_ÀOB�OT_ISOLC��NTV@A'qhuN�AME�l��o�JO�B_ORD_NU�M ?�X#q�H768  �j1Zc@�r
��rV�s���r�?�r?��r�pÀPC_TI�MEu�a�xÀS2�32>R1�� �LTEACH PENDANw��:GX�!O �Maintena�nce Cons�j2����"��?No UseB�׏ ������1�C�y�V��NPO�P@�YQ��cS�CH_Lf`�%^ �	ő~��!UD1:�z��R�@VAIL�q�@�Ӏ�J�QSPA�CE1 2�ż ��YRs�i�@Ct��YRԀ'{��8�?��˯���� "���7�2�c�u����� G���߯ѿ򿵿�(� �u�AC�c�u����� Ͻ�߿���ϵ��(� �=�_�qσϕ�C߹� �����߱��$��9� [�m�ߑߣ�Q����� �߭��� ���	�W�i� {���M�������5� ��.S�e�w��� ��I������� *?as��E �����/&// ;/]o����� �/2/�/?"?�/7?Y/ k/}/�/�/O?�/�/�?��?�?O0OOKA�o�*SYPpM*��8.30261 �yB5/21/2018 A �WP�fG|�H�_TX`�� !$COMM�E�$US�Ap $EN�ABLEDԀ$sINN`QpIOR�B��@RY�E_SIG�N_�`�AP�AIT\�C�BWRK�BD<��_TYP�CRIN�DXS�@W�@%VF{RI{�_GRPԀ$UFRAM�r�SRTOOL\VMY�HOL�A$LE�NGTH_VTE�BTIRST�T ? $SECLP�X�UFINV_PO�S�@$MAR�GI�A$WAI�T�`�ZX2�\�VG-2�GG1�AI�@�S��Q	g�`_WR�BNO_USE_DI�B^uQ_REQ�BC�C�]S$CUR_T�CQP�R"a^f �G�P_STATUS>�A @ �A3`X�BLk�H$zc1�h��P@���@_�F�X �@E_MLoT_CT�CH_�J6�`CO�@OL�E�C�GQQ$W�@w��b#tDEADLO�CKuDELAY_CNT�a3qGt�a�$wf 2 �R1[1$X<�2*[2�{3[3$Zwy �q%Y�y�q%V�@�c�@��b$V�`�RV�UV�3oh>b�@ � q�d�0arMSKJ��LgWaZ�C`NRK�P�S_RATE�0�$���S
`�Q�TAC���PRD���e�SD*��a4�A�0�DG�A� 0�P�flp bquS2ppI�#`\
`�P 
�S\`�  �A�R_�ENBQ ��$RUNNER_SAXI�<`ALPL�Q��RU�THICQ�$FLIP7��DT�FEREN��R�IOF_CHSU�IW��%V)�G1����$P�řA�Q�Pݖ_J�F�PR_P�	�RV_DATA�A�  $�E�TIM���$VA�LU$�	�OP_ �  �A�  2 �S�C*�	� �$ITP_!�SQ]P�NPOU}�o�TOT�L�o�DSP��JO�GLIb��PE_P�Kpc�Of�i��PX�]PTAS�$KE?PT_MIR��¤2"`M�b�APq�aE�@�y�q�g@١c�vq�PG�BRK6��x���L�I��  �?�SJ�q�P�ADE�z�ܠBSOCz�M�OTNv�DUMM�Y16Ӂ$SV��`DE_OP��S�FSPD_OVR4
���@LD�����OR��TP8�LEb��F������OV��CSF��F����bF��d�ƣ&c)�fQc�LC�HDLY��REC�OV���`��W�PM��gŢ�RO�������_F�?� @v�S� �NVER�@�`O�FS�PC,�CSWD�ٱc�ձ���B����T�RG�š�`E_F�DO��MB_CM4}���B��BLQ�¢�	�Q�̄Vza�BUP��g��G
��AM����@`KՊ�e�_M�!�d�AMf�Q��T�$CA����DF����HBKd�v���I�OU��I'R��PA����������p���~��DVC_DB�S�!�x�Q�!�s�d�9�1�A��9�3A��AT�IO�0��͠��U0S����WaAB��R�+c�`tá`DؾA��_�AUXw�SUBCPUP���S�`�����3Եжc���3�FLyA�B�HW_Cwp�"�Ns&�]sAa��_$UNITS�M�>F�ATTRIz�Z�ެ�CYCL�CNE�CA���FLTR�_2_FI��TARTUPJp����Aƴ�LP������_S�CT*cF_F�F_P���b�FS��+�K�CHA/Q��*�d�RSD��Q�����Q���_TH�PRO8r���հEMPJ���rG�T� ��Q�DI�@y�RAOILAC/�bMX�CLOf�xS��ځ����拁���PR#�S�`app�C� {	��FUNC���RIN`QQP� �ԱRA)]R ���AƠ��AWAR�֓��BLZaWrA0kg�ngDAQ�B�rkLD�र&q��M�K���TI����j��$�@R�IA_SW��AF
��Pñ#��%%�p89r1��MOIQ���gDF_~P(�PD"�LM-�FA�PHR�DY�DORG�H�; _QP�s%MULCSE~Pz���*�� �J��Jײ��FAN_ALMLVG���!WRN�%HARDP��UcO�� K�2$SHADOW�]�kp�a02��� ST�Of�+�_^�w�AU�{`R��eP_SBR�z5���:F�� ��3MPINF?�p\�4��3REGV&/1DG�+cVm �C��CFL(��?�D�AiP���Z`�� �8����Z�	 �P(Q�$�A$Z�Q �V�@�[�
� ���EG��o���kAAR���㌵2�axG���AXE��ROB.��RED��W�QD�_�Mh�SYA��AF�:�FS�GWRI�P~F&�STR����E�˰EEH�)��D�a\2BkPB6P��=V��DvЗOTO�1)���ARYL�tR�v�3����FI&�ͣ$LI�NKb!\��Q�_�3S���E��QXY�Z2�Z5�VOFF����R�R�XxPB��ds�G�cFI�03g�������_J��'�ɲ�S�&qR0LTV[6���aT�Bja�"�bC���D�U�F7�TURB� X��e�Q�2XP�ЊgFL�E���x@��`�U9Z8���� +1	)�K��Mw��F�9��劂����OR!Qj��G;W3��� #�Ґd ���uz����1N�tOVE�q_�M�� ё?C�uEC�uKB�v'0 �x-�wH��t��� & `��qڠ�B�ё�u��q�wh�ECh����E)R��K	�EP�$���AT�K�6e9`e�W���AXs� '��v�/�R ��� �!�� ��P��`�@�`�3p�Yp�1�p �� �� �� (��  8�� H�� X�� h�� �x�� ������DEBU�$%3�I��·RAB���ٱ�s9V��� 
d�J� ����@񘧕������ �Q���a���a��3q���Yq+$�`%"<�cLA�B0b�u�'�GR�O���b<��B_ s��"Tҳ*`�0A�u�p�uq�p1}�ANDGp��������U��p1��  �ѷ0�Qθuݸ��P�NT0���SERsVE �Z@ $`�EAV�!�PO ����nP!�P@�$!�Y@  $.>�TRQ�b
=��B2G�K�%"2\��~� _  l���5�D6ERRVb(�I��V0`;���TOQ:�7�L�@
�R��e %G�%�Q�� <�50�F� ,�`�z��>�RA� 2� d!�����S�  M��pxU �����OCuG�  }��COUNT6Q���FZN_CFG�F� 4#��6��T G4�_�=�����Î�^VC ���M ��"��$6��q ��F!A E� &��X�@� ������A����A9P��P@HEL�0�ҿ 5b`B�_BAS��RSR�6�CSH����1�Ǌ�2��3��4���5��6��7��8��}�ROO����Pf�PNLEA�cAB)�ܫ ��ACKu�IN2O�T��(B$UR0� =�_PU��!0��OU+�Pd�8j���� V��TPFWD�_KAR��� ��R�E(ĉ P�P�>QUE�:RO�p�`r0P1I� x�j�P�8f��6�QSEM��0t��� A��STYL�3SO j�DIX�&p�����S!_TMC�MANRQ��PE�NDIt$KEY?SWITCH����kHE�`BEA�TM83PE{@LEP��>]��U��F���SpDO_HOeM# O�@�EF�p�PRaB�A#PY�C�� O�!���OV_�M|b<0 IOCM��dFQ�h�HKYA D�Q�7��	UF2��M���p�c�FORC�3WAR�"�OM|@ � @S�#o0U)SP��@1�2&3&4RE���T�O��L�y��8UNLOv��D4K$EDU1  ��SY�HDDN�F� M�BLO�B  p�SN�PX_AS�� �0@�0��81$S{IZ�1$VA{�~��MULTIP-���# A� � $��� /4`��BS��0�C���&F'RIFBO�S����3� NF�ODBUP߰�%@3;9(���܋�Z@ x��SI���TEs�r�cSG%L�1T�Rp&�Н3xB��@�0STMTq2�3Pg@VBW�p�4�SHOW�5@�SmV��_G�� 3p�$PCJ�PИ���F�B�PHSP A�W�EP@VD�0WC�� ���A00 ��PB XG XG XGT$ XG5VI6VI7VIU8VI9VIAVIBVI@�XG�YF�0XGFVH���XbI1oI1|I1��I1�I1�I1�I1��I1�I1�I1�I1��I1�I1Y1Y2�UI2bI2oI2|I2�I2�I�`�X�I2p�X��I2�I2�I2�I2
�I2Y2Y�p�hbIU3oI3|I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3�IU3Y3Y4�i4bIU4oI4|I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4�IU4Y4Y5�i5bIU5oI5|I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5�IU5Y5Y6�i6bIU6oI6|I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6�IU6Y6Y7�i7bIU7oI7|I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7�I�7Y7T�VP� UD�y"ՠ��Q
<A62��t��R��CMD� ��Mb5�Rv�]��Q_hЁR���e����<�Y�SL���  � �%\2��+4�'��xW�BVALU���b��'���FH�ID�_L���HI��I���LE_��㴦��$0C�SAC��! h �VE_BLCK��1>%�D_CPU5ɧ  5ɛ �����C�� ���R " � �PWj��#0��LA��1SBћì���R?UN_FLG�Ś� ���ĳ ���������šH���Х��T�BC2��# � @ B��e �S�88=�FTDC�����V���3d�Q�TH�F�����R�L�ESERVE9��F���3�2�E��Н��X -$��LEN`9��F��f�RA��LW"G�W_5�b�1�њд2�MO-�T%S60U�Ik�0�ܱF�����[�DEk�21LA3CEi0�CCS#0�� _MA� j��z玤�TCV����z�T �������.Bi�'A�$z�'AJh�#EM5���J��@@i�V�z���2Q �0&@o�h��JK��VK9��{����щ�J0����J�J��JJ��AAL����������4��5�ӕ N1������J.�LD�_�1* v�CF�"% `�GROU���1�A�N4�C�#m REQ�UIR��EBU��#��6�$Tk�2�$���zя #�&{ \�APPR� �C� 0�
$OPE=N�CLOS��St��	i�
��&' �MfЩ���W"N-_MG߱7CB@��A���BBRK�@NOLD@�0RTMO_5ӆp1	J��P�����@���������6��1�@ )!�#�(� ������'��+#PATH ''@!6#@!�<#� � 9'��1SCA��l�6IN��UCJ�[1� C0@UM�(Y  ��#�"�����*���*���� PAYLOA�~J2LؠR_A	N^�3L��91�)�1AR_F2LSHg2B4LO4�!F7��#T7�#ACRL_@�%�0�'�$��H���.�$HA�2FL�EX��J!�) P�2�D߽߫��|�0��* :�� ��z�FG]D����z���%�F1]A�E�G4�@F�X�j�|���BE�� �����������(� �X�T*�A���@�XI��[�m�\At�T$g�QX <�=��2TX���emX �������������������+	�J>+ �-�K]o|�٠cAT�F�4�ELFP�Ѫs�J� *� J�EmCTR�!�AT�N�vzHAND_VB.��1��$7, $8`F2Avԍ��SWu	#-?� $$M*0. �]W�lg��PZ����A��� 1����:QAK��]AkAzP��LN�]DkDzePZ G��C�ST_hK�lK�N}DY�� � A����0��<7]A <7W1�'��d�@g`�P�������t"
"J"�. M��2D%"p�H��~�AS�YMj%0�� j&-��-W1�/_�{8�  �$�����/�/�/�/ 3J<�:9�/�89.�D_VI�v��>��V_UNI�ӛ��cD1J����╴�W< ��n5Ŵ�w=4��9���?�?<�uc�4�3d�%�H���/��j��0�DIzuO�� �k�>0 �`��I��A��#�� �@ģ���@���IPl� 1 � /�ME.Qp��9�ơT}�PT�;pG �+ Gt� ���'���T�0 $D�UMMY1��$�PS_�@RF�@ � G b�'FLA�@ YP(c|��$GLB_TP�ŗ����9 P�q��2 �X� z!ST9�� SBRM M21�_V�T$SV_�ER*0O�p����C)L����AGPO��f��GL~�EW>�3 �4H �$YrZBrW@�x�A1+�A���"j� �U&�4 �8`NZ�"�$GIn�p}$&� -�8 �Y�>�5 LH {��}$F�E��NWEAR(PN�CF��%PTANC�B	!JsOG�@� 6.@$JOINTwa�?pd�MSET>�7�  x�E��HQtpS�{r��up>�8� ��pU.Q?�� L?OCK_FOV06�ޅ�BGLV�sGL�t�TEST_XM�� 3�EMP��8���_�$U&@%�Fw`24� Y��5��h2�d��3��CE- |���� $KAR�Q}M��TPDRA)�����VECn@��kIU��6��HEf�OTOOL�C2V�D;RE IS3ER96��@ACH� �7?Ox �Q�29�Z�H I�  @�$RAIL_BO�XEwa�ROB�O��?��HOW�WAR�1�_�zROLMj��:qw�pjq� �@ O_Fkp�! d�l>�9��� �R O8B:� �@�	""�O%U�;�Һ�3ơ�r|�q_�$PIP��N&`H�l�@��~#@CORDEDd��p >f�fpO�� �< D ��OB ⁴sd���Kӕ����qSYS�ADqR��f��TCHt�� = ,8`ENTo��1Ak�_{�-$xCq_�f�VWVA��?> �  &���PREV_RT~�$EDITr&_VSHWRkq��(� &R:�v�D��JA��$�a$HEA�D�6�� �z#K�E:�E�CPSPD.�&JMP�L~��0R*P��?��1%&�I��S�rC�pNEx; �q�wTICK�Cb��M�13�3HN��@ @� 1Gu�!�_GPp6��0STY'"xLO��:�2|l2?�A t 
m MG3%%$R!{�=��S�`!$��w`��Ȃճ���Pˠp6SQ�U��E��u�TER�C�0��TSUtB ����hw&`gw��Q)�pO����@I�Z��{��^�PR`�kюB1XPU��ΞE_DO��, XS:�K~�AXI�@���UR�pGS�r� �^0�&��p_) �EET�BPm��o��0�Fo��0A|����Rԍ��a;�SR�Cl>@P��b _�yUr��Y��yU��yS ��yS���UЇ�U���U ���U�]��Ul[��Y�bXk�]Cm������YRSC�� D h�DS~0��Q�3SP���eATހ����A]0,2N�ADD�RES<B} SH�IF{s��_2CH����I��=q�TVsrI��E"���aT�Ce�
��
;�VW��A��F \��q� �0l|\A@�rC�_B�"R{zp�ҩq�TX_SCREE�Gv�=�1TINA����t{�c��A�b?�H T1�ЂB������I��A��BE�y RR�O������� B��Š�
�UE4I ��g�!p�S��RSyM]0�GUNEX(@~Ƴ�j�S_S�ӆ�� Á։񇣣�ACY��0� 2H�pUE�;�J�����@GM�T��Lֱ�A��O^	�BBL_| W8�N��K ��0s�OM��LE/r��� TyO!�s�RIGH���BRD
�%qCKG9R8л�TEX�@��>��WIDTH�� ��B[�|�< �U�I_��Hi� L 8K���_�!=r���R:�_��Y�1R�O6q�Mg0璴�U��h�Rm��L�UMh��FpERV�w �P���`�Nz��&�GEUR��iFP)�)� LP��(RE%@�a)ק�a�P!��f �5�6�7�8Ǣ#B�É@����tP�fW�S@�M�USR&�O <����U�Qs��FOC)��PRI�;Qm� :���TRI}P�m�UN��
��Pv��0��f%�p�'���@�0 Q�\���AG �0T� ��a>q�OS�%�R Po���8�R/�A� H�L4N���U¡��SU�g��¢5��OSFF���T�}�=O�� 1R���:��S�GUN��}6�B_SUB?Ҝ�В�SRTN�`TU0g2��mCOR| D�'RAUrPE�TZ�#'��VCC��	3V �AC36MFB�1�%d�PG �Ws (#��ASTEM�a����0PE��:T3G�X �\ �ڏMOVEz�A��A�N�� ���M���LIM_X��2��2� �7�,�����ı�
�BVF�`E���~��024Y��IB�7��
�5S��_Rp� 2�^�� WİGp�+@��}СP��3�ZGx ���3����A�ݠCZ�D#RID����Vy08��90� De�MY_UBYd���6��@��!��X��P_Sh��3��L�KBM,�$+0DEY(#E�X`�����UM_M�U� X����ȀUSн� ���G0`PACI���а@��:��`:,�:����RE/��3qL�+��:[^��TARG��P�r���R<�\ d�`��A��$�	��ARF��SW2 ��-���@Oz�%qA7p�yREEU�U�01�,�+HK�2]g0�0qP� N� �EAM0G�WOR���MR�CV3�^ ���O*�0M�C�s	���|�REF_��� x(�+T� ����������3_RC H4(a�P�І�hrj�pNA�5��0�_ ��2�����L@��n�@@OAU~7w6���Z�6�a2[��RE�p�@F;0\�c�a'2K�@WSUL��]��C��f0�^��� NT�� L�3��(6I�(6q�(3� L��Q5��Q5I�]7Jq�}�Tg`4D`�0�.`0�AP_HU�C�5SA��CMPBz�F�6�5�5�0_�aAR��a�1I\!X�9��GFS��ad� ��M��0p�U�F_x��B� �ʼ,R�O��Q��'����URF�3GR�`.�3IDp���)�D�;��A,��~�IN��H{D���V@AJ���S͓UWmi=�����TY&LO*�5���󾖄bt +�cP�A� �cCACH�vR�UvQ��Y���p�#CF�I0sFR��XT���Vn+$HO����P!A3�XB�f�(1 ���$�`VPxy� ^b_SZ3132he6K3he12J�eh� chG�chWA�UM�P�j��IMG9�uPAD�iiIMRyE�$�b_SIZ�$�P����0 ��ASY�NBUF��VRT�D)u5tqΓOLE�_2DJ�Qu5R��C���U��vPQuEwCCUlVEMV x�U�r�WVIRC�aIuVTPG���rv01s��5qMPLAqa�R�v�V0�c��� _CKLAS�	�Q�"��d  �ѧ%ӑӠ@}¾�$�Q���Ue |�0!�rSr��T�#0! �r�iI���m�vK�BG��VE�Z�PK= �v�Q��&�_HO�0��f � >֦3�@Sp��SLOW>�R=O��ACCE���!� 9�VR�#���p:����AD�����PA�V�j�� D����M�_B"���^�JMP�G ��g:�#E$SSC��x&�vPq��IhݲvQS�`qVN���LEXc�i T�`�sӂ��Q�FLmD �DEsFI��3�02���:����VP2�Vj� ��A��V�4[`MV_PIs��t����A�@��FI��|�Z ��Ȥ�����A���A���~�GAߥ1 LOO��1 JCB���Xcx��^`�#PLANE��R��1F�c�����pr�M� [`�噴��S����f����Af��R��Aw�״tU��pR�KE��d�VANC��EM�V���� �k���ϲ�BR;_AA� l��2�� ��p�#�����m h�@��O K�$����2��kЍ0OU&A�"eA�
p�pSK�T�M@FVIEM 2l� ��P=���n �<<��dK�UMM�YK1P��`D6�ȟ�CU��#A�U��o $��T�IT�$PR�����OP���V�SHIF�r�p`J�Qsԙ�fOxE[$� _R�`U�# ����s��q������ G�"G�޵'�T�$��SCO{D7�CNT Q i�l�>a�-�a�;� a�H�a�V���1�+�2u1��D���� w � SMO�U�q��a�JQ���%��a_�R[�r�n׍*@LIQ�AA/`��XVR��s�n�T�L���ZABC��t�t�c�
L�Z�IP��u���LV�bcLn"�is ��ZMPCFx�v�:�$�� ���D�MY_LN����s8���@y�w Ђ(a\�u� MCM�@Cbc�CART_�DP~N� $J71D��=NGg0S�g0�BUXW� ��U�XEUL|B yX���	��A=Z��x 	����m�YH�Db  �y 80���0EI3GH�3n�?(� H�r���$z ���X|�����$B� Kd'b��_��L3�RVS�qF`���OVC��2'�$|�>P&��
hq���5D�TR�@r �V�1�SPHX��!{ ,� *<��$R�B2 2 ����C!��  �@L�V+@b*c%g!`+�g"�`V*�,8�?�V+�/V.�/@�/?�/�/V(7%3@/ R/d/v/�/6?�/�/�?��?�?O4OOION;4 ]?o?�?�?�?SO�?�? �O_�O0_Q_8_f_N;5zO�O�O�O�Op_�O _o8o�_MonoUo�oN;6�_�_�_�_�_�o o%o4Uj�r�N;7�o�o�o�o�o � BQ�r�5���������N;8���� �Ǐ=�_�n���R����ş��ڟN;G N� џ�
����?���W�i�{��� ����ï�.�������A��dW�<�N� |�������Ŀֿ�ޯ ���0�B�_�R�d� 꿤϶����������� ��*�L�^��rτ� 
�������������&�8�J�l�~� `ҟ @�з�����ߩ��-����&� ,���9�{�����a� ��������������A 'Y���� �����a�#1�
��N;_M?ODE  ��/S ��[�Y�B���
/\/*	�|/�/R4CWORK�_AD�	��^T1R  ����� �/� _INTV�AL�+$��R_�OPTION6 ��q@V_DA�TA_GRP 2Y7���D��P�/ ~?�/�?�9��?�?�? �?OO;O)OKOMO_O �O�O�O�O�O�O_�O _7_%_[_I__m_�_ �_�_�_�_�_�_!oo Eo3oioWoyo�o�o�o �o�o�o�o/ eS�w���� ���+��O�=�s� a�������͏���ߏ ��9�'�I�o�]������$SAF_D?O_PULS� ��~������CAN_GTIM����Α�R ��Ƙ_��5�;#U!P"�1!��� �?E�W�i�{����� .�ïկ�����'(+~�T"2F��"�dR�I�Y��2�o+@a얿����)�u�� k0ϴ��_; ��  T� �� �2�D�)�T D��Q�zόϞϰ��� ������
��.�@�R߀d�v߈ߚ�/V凷�����߽���R�;�o ��W�p��
�t���Diz$� �0 � �T"1!�� ����������� ����*�<�N�`�r� �������������� &8J\n�� ������"4FX ��࿁� ������/` 4�=/O/a/s/�/�/�/@�/�/�/�!!/ �0޲ k�ݵu�0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ ok$o6oHo Zolo~o�o�o�o�o1/ �o�o 2DVh z�/5?����� ���&�8�J�\�n� ��������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	���-�?�Q�c�u��� ���`Ò�ϯ��� �)�;�M�_�q�����@����˿ݿ� �����3� ���&2�,��	1234�5678v�h!�B!��2�C
h���0�ϵ��� �������!�3�9ѻ� \�n߀ߒߤ߶����� �����"�4�F�X�j� |�h�K߰��������� 
��.�@�R�d�v��� ����������� *<N`r��� ����&�� J\n����� ���/"/4/F/X/ j/|/;�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�/�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ �?L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o=_�o�o�o�o �o�o 2DVh�z�����h� �����u�o.�@�R����Cz  B���   ���2�&� � _�
~���  	�_��2�Տ����_�%p������ďi� {�������ß՟��� ��/�A�S�e�w��� ������N������ +�=�O�a�s������� ��Ϳ߿���'�9�DK�_������<v��_��$SCR_G�RP 1
�� �� t{ ��� ���	 �����������������_������)�a�����&�DE� �DW8���l�&�G��CR-35iA� 9012345�67890��M�-20��8��C�R35 ��:�
������������� ��:֦�Ӧ�G���&������	��]�o������:���#H���>�����������&���ݯ:� �j����g������B�t����������9A����  @�`���@� ( ?��=��Ht�P
��F?@ F�`z� y������ � $H��Gs^p��B��7� �/�0//-/f/Q/ �/u/�/�/�/8���P�� 7%?����"?W?x-2?<���]?� H�1�?t�ȭ7��������?-4A , �&E@�<�@G�	B-1 3OZOlO-:�HA�H�O�O|O P�B(�B�O�O_���EL_DEFAU�LT  �����`SHOTSTR#]JA7R�MIPOWERFOL  i�/UYToWFDO$V /U�RRVENT 1�����NU �L!DUM_E�IP_-8�j!?AF_INE#P�_�-4!FT�_->��_;o!��`o ��*o�o!RPC_OMAIN�ojh�vo��o�cVIS�oii���o!TPpP�U�Ydk!
�PMON_PROXYl�VeZ�2r��]f��!R?DM_SRV��Y9g�O�!R��k���Xh>���!
�`M���\i���!R�LSYNC�-9�8֏3�!ROS̽_-<�4"��!
�CE4pMTCOMd���Vkn�˟!	��OCONS̟�Wl����!��WASR�C��Vm�c�!N��USBd��XnR� ��Noӯ�������!���E��i�0���WR�VICE_KL �?%�[ (%SVCPRG1��D-:Ƶ2ܿ�˰3�D	�˰4,�1�˰5T�DY�˰6|ρ�˰7�� ��˰�����9����ȴf�!�˱οI�˱ ��q�˱ϙ�˱F��� ˱n���˱���˱�� 9�˱��a�˱߉�� 7߱��_������ ��)����Q���� y��'���O���� w������� ��˰��İd�c�� ����=( as^����� �/�/9/$/]/H/ �/l/�/�/�/�/�/�/ �/#??G?2?k?V?}? �?�?�?�?�?�?O�? 1OCO.OgORO�OvO�O �O�O�O�O	_�O-_��_DEV �Y��MC:5Xd��GTGRP �2SVK ��bx 	� 
 ,�PK 5_�_�T�_�_ �_o�_'o9o o]oDo �ohozo�o�o�o�o�o �o5{�_g� �������� �?�&�c�u�\����� ��Ϗ���J\)��� M�4�q���j�����˟ ݟğ��%���[� B��f������ٯ�� �����3��W�i�P� ��t���ÿ���ο� ��A�(�e�L�ί�� RϿ��ϸ������ � �O�6�s�Zߗߩߐ� �ߴ������'�~ϐ� ]���h������ �������5��Y�@� R���v���������@� 	��?&cu\ ������� �;M4qX�� �����/�%// I/[/B//f/�/�/�/ �/�/�/�/�/3??W? �L?�?D?�?�?�?�? �?O�?/OAO(OeOLO �O�O�O�O�O�O�O�O�_iV �NLyٿ6 * 		S=?>��+c"_VU�@Tn_Y_B���B�2�J�j~Q�´~_g_�_�Q%JOGGING�_��^7T(?VjZ��Rf��Y��� /e�_%o7e�Tt�]/o �o{m�_�o�m?Qi�o��o;)Kq%��o�}os��� ���9�{`��)� ��%���ɏ���ۏ� S�8�w��k�Y���}� ��ş���+��O�ٟ C�1�g�U���y����� ��'����	�?�-� c�Q���ɯ����w��� s����;�)�_ϡ� ��ſOϹϧ������� ��7�y�^ߝ�'ߑ� ߵߣ��������Q� 6�u���i�W��{�� �����=��M���A� /�e�S���w������� �����=+a O������u�� �9']�� �M������ /5/w\/�%/�/}/ �/�/�/�/�/=/"?4? �/?�/U?�?y?�?�? �??�?9?�?-OO=O ?OQO�OuO�O�?�OO �O_�O)__9_;_M_ �_�O�_�Os_�_�_o �_%oo5o�_�_�o�_ [o�o�o�o�o�o�o! coH�o{�� ����; �_� S�A�w�e�������я ���7���+��O�=� s�a������П��� ��'��K�9�o��� ����_���[�ɯ��� #��G���n���7��� ������ſ����a� Fυ��y�gϝϋϭ� ������9��]���Q� ?�u�cߙ߇ߩ���%� ��5���)��M�;�q� _���߼��߅���� ��%��I�7�m���� ��]�����������! E��l��5�� �����_D �we���� �%
//���=/ s/a/�/�/�/��/!/ �/??%?'?9?o?]? �?�/�?�/�?�?�?O �?!O#O5OkO�?�O�? [O�O�O�O�O_�O_ sO�Oj_�OC_�_�_�_ �_�_�_	oK_0oo_�_ co�_so�o�o�o�o�o #oGo�o;)_M o����o�� ��7�%�[�I�k��� �������ُ��� 3�!�W���~���G�i� C����՟���/�q� V������w������� �ѯ�I�.�m���a� O���s�������߿!� �E�Ͽ9�'�]�Kρ� oϑ�����Ϸ�� ��5�#�Y�G�}߿Ϥ� ��m���i������1� �U��|��E��� ������	���-�o�T� �����u��������� ��G�,k���_M �q���� ���%[Im ���	���/ /!/W/E/{/��/� k/�/�/�/�/	??? S?�/z?�/C?�?�?�? �?�?�?O[?�?RO�? +O�OsO�O�O�O�O�O 3O_WO�OK_�O[_�_ o_�_�_�__�_/_�_ #ooGo5oWo}oko�o �_�oo�o�o�o C1Sy�o��oi �����	�?�� f�x�/�Q�+���Ϗ�� ���Y�>�}��q� _�������˟���1� �U�ߟI�7�m�[�}� ���ǯ	��-���!� �E�3�i�W�y�ϯ�� ƿ��������A� /�eϧ���˿UϿ�Q� ��������=��d� ��-ߗ߅߻ߩ����� ���W�<�{��o�]� ���������/�� S���G�5�k�Y���}� �������������� C1gU������ {����	?- c���S��� ���/;/}b/� +/�/�/�/�/�/�/�/ C/i/:?y/?m?[?�? ?�?�?�?? O??�? 3O�?COiOWO�O{O�O �?�OO�O_�O/__ ?_e_S_�_�O�_�Oy_ �_�_o�_+oo;oao �_�o�_Qo�o�o�o�o �o'ioN`9 ������A &�e�Y�G�i�k�}� ����׏���=�Ǐ1� �U�C�e�g�y���� ֟���	���-��Q� ?�a���ݟ��퟇�� ϯ��)��M���t� ��=���9���ݿ˿� �%�g�Lϋ���m� �ϑϳ�������?�$� c���W�E�{�iߟߍ� �������;���/�� S�A�w�e�������� ������+��O�=� s������c������� ����'K��r�� ;������� #eJ�}k� ����+Q"/a �U/C/y/g/�/�/�/ /�/'/�/?�/+?Q? ??u?c?�?�/�?�/�? �?�?OO'OMO;OqO �?�O�?aO�O�O�O�O __#_I_�Op_�O9_ �_�_�_�_�_�_oQ_ 6oHo�_!o�_io�o�o �o�o�o)oMo�oA /QSe�����%{,p�$SE�RV_MAIL + +u!��+q��OUTPUT��$�@�RV �2�v  $� �(�q�}��SAV�E7�(�TOP10� 2W� d �6 *_�π( _������#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u����������Ͽݷ��YP���'�FZN_CF�G �u�$�~����GRP� 2�D� ,�B   A[�+qD�;� B\�� � B4~�RB{21��HELL�C�u��j�k�2�|����%RSR�� �����
�C�.�g�R� ��v߈��߬�����	����-�?�Q��  �_�%Q���_����,p����Sޖ�g�2,pd��|���HK 1�� ��E�@�R�d� ���������������� *<e`r�~��OMM ������FTOV_E�NB�_���HOW_REG_UI��(�IMIOFWD�L� �^�)WAIT���$V1�r^�NTIM7���VA�_>)_UNIT��v��LCTRY�B�
�MB_HD�DN 2W� 2�:%0 �pQ/�q L/^/�/�/�/�/�/�/��/�"!ON_AL�IAS ?e�	f�he�A?S?e?w? �:/?�?�?�?�?�?O O&O8OJO�?nO�O�O �O�OaO�O�O�O_"_ �OF_X_j_|_'_�_�_ �_�_�_�_oo0oBo To�_xo�o�o�o�oko �o�o,�oPb t�1����� ��(�:�L�^�	��� ������ʏu�� �� $�Ϗ5�Z�l�~���;� ��Ɵ؟����� �2� D�V�h��������¯ ԯ���
��.�ٯR� d�v�����E���п� ��ϱ�*�<�N�`�r� ϖϨϺ���w���� �&�8���\�n߀ߒ� ��O����������� 4�F�X�j�|�'��� ���������0�B� ��f�x�������Y��� ������>Pb t������ (:L�p� ���c�� // $/�H/Z/l/~/)/�/ �/�/�/�/�/? ?2?�D?V?]3�$SMO�N_DEFPRO ���1� *SYSTEM*0�m6RECALL� ?}9 ( ��}tpdis�c 0=>147�.87.149.�40:13148� 8 �>2204y �1�95172]?�O+M}tpconn 0 �?�?�?��?�O�O4G
xyz�rate 11 �JO\OnO�O_#_6E�E61�?�A�O�O_ �_�_�NJ_\_n_�_o #o6_H_�_�_�_�o�o�4G9copy f�rs:order�fil.dat �virt:\tm?pback\Io�A�yo
/L0�bmd�b:*.*�o�o `�o��8C4x�d:\H�pZ�At�\�)� }5�ua� ��F�������JJ� \�n����#�6oHoZo ����������_X�j� |���2�D�֟��� ������B�ɟ[�m����"�5�G�12532ޯ������8C�? R�]�o����$�7Oɿ ۿ����Ϣϵ��NX� j�|���2�D�V��� �ϋߝ߰�T�f�x� 	��.�@�������� ��,ﾯP�b�t����)� }?��E2896 ���������8���S�\�n��� #6����������� ����Wi{1� C�U�������� Sew�/-?� ��/�/�/�O/a/ s/�/?(?;/�/�/�/ ?�?�?�/K?]?o?�? O$O7?I?�?�?�?�O�O�f8�o�oIO[AyO
__�l/?�ORI�O_�_�_�d3�ҏNM s_�_o(o�yG��_� �_o�o�o�O�OW_r_ �o':_�o^_�o����b�$SNP�X_ASG 2�����q�� P 0 �'%R[1]�@1.1��y?��s%�!��E�(�:� {�^�������Տ��ʏ ���A�$�e�H�Z� ��~���џ����؟� +��5�a�D���h�z� ����ů�ԯ���
� K�.�U���d������� ۿ������5��*� k�N�uϡτ��ϨϺ� �����1��U�8�J� ��nߕ��ߤ������� ���%�Q�4�u�X�j� ������������� ;��E�q�T���x��� ��������% [>e�t��� ���!E(: {^������ /�/A/$/e/H/Z/ �/~/�/�/�/�/�/�/ +??5?a?D?�?h?z? �?�?�?�?�?O�?
O KO.OUO�OdO�O�O�O �O�O�O_�O5__*_ k_N_u_�_�_�_�_�_ �_�_o1ooUo8oJo��ono�o�o�d�tPA�RAM �u}�q �	��jUP�d9p�ht���pOFT_KB_CFG  �c��u�sOPIN_S_IM  �{v�n��p�pRVQSTP_DSBW~�r"t�HtSR �Zy � &�!pINGS EL�_5SEM����vTOP_ON_?ERR  uCy~8�PTN Zu�k�A4�RN�_PR�D��`�VCNT_GP �2Zuq�!px 	r��ɍ���׏���wVD��RP 1	�i p�y��K� ]�o���������ɟ۟ ����#�5�G�Y��� }�������ůׯ��� ��F�C�U�g�y��� ������ӿ��	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�qߘߕߧ߹��� ������%�7�^�[� m����������� ��$�!�3�E�W�i�{� �������������� /ASew�� �����+ =Ovs���� ���//</9/K/ ]/o/�/�/�/�/�/�/ ?�/?#?5?G?Y?k? }?�?�?�?�?�?�?�?�OO)�PRG_CoOUNT8v�k��GuKBENB��FEM�pC:t}O_UPD �1�{T  
 4Or�O�O�O__!_ 3_\_W_i_{_�_�_�_ �_�_�_�_o4o/oAo So|owo�o�o�o�o�o �o+TOa s������� �,�'�9�K�t�o��� ������ɏۏ���� #�L�G�Y�k������� ��ܟן���$��1� C�l�g�y��������� ӯ����	��D�?�Q� c���������ԿϿ� ���)�;�d�_�q��=L_INFO 1��E�@ �2@����������� �ٽ`y*�d��h'���¿���=`y;MY?SDEBUGU@�@����d�If�SP_�PASSUEB?~x�LOG  �ƕ�C��*ؑ� � ��A��UD�1:\�ԘΥ�_M�PC�ݵE&�8�A���V� �A�SAV !�������X����SVZ�TE�M_TIME 1u"���@ 0��-�X��X�X�����$T1SVGU�NS�@VE'�E���ASK_OPT�IONU@�E�A�A�+�_DI��qOG�B�C2_GRP 2�#�I�����@� � C���<Ko�CF�G %z��� 8�����`��	� .>dO�s� ������* N9r]���� ���/�8/#/\/ n/��Z+�/Z/�/�/H/ �/?�/'??K?]�k? =�@0s?�?�?�?�?�? �?O�?OO)O_OMO �OqO�O�O�O�O�O_ �O%__I_7_m_[_}_ _�_�_�X� �_�_o o/o�_SoAoco�owo �o�o�o�o�o�o =+MOa��� ������9�'� ]�K���o��������� ɏ���#��_;�M�k� }��������ß�ן ��1���U�C�y�g� �������������� 	�?�-�c�Q�s����� �����Ͽ���� )�_�Mσ�9��ϭ��� ����m���#�I�7� m�ߑ�_ߵߣ����� ������!�W�E�{� i������������ ��A�/�e�S�u�w� ������������+ =O��sa��� ����9' ]Kmo���� ���#//3/Y/G/ }/k/�/�/�/�/�/�/ �/??C?��[?m?�? �?�?-?�?�?�?	O�? -O?OQOOuOcO�O�O �O�O�O�O�O__;_ )___M_�_q_�_�_�_ �_�_o�_%oo5o7o Ioomo�oY?�o�o�o �o�o3!CiW ������� ��-�/�A�w�e��� �������я��� =�+�a�O���s����� ��ߟ͟��o�-�K� ]�o�ퟓ�����ɯ����צ��$TBC�SG_GRP 2�&ץ� � �� 
 ?�  6�H�2�l� V���z���ƿ��������(�d��E+�?�	 H�C���>����G����C�  Aq�.�e�q�C��>�'�33��S�/]϶��Y��=Ȑ� C\ g Bȹ��B����>����P���B%�Y�z��L�H�0�$����J�\�n�����@�Ҿ������� ��=�Z�%�7�����?3�����	�V3.00.�	�cr35��	* ����
��������� 3��4�   {�CT�v�}��J2�)����~��CFG +ץ�'� *�������I����.<
�<bM �q������ �(L7p[� �����/� 6/!/Z/E/W/�/{/�/ �/�/�/.�H��/?? �/L?7?\?�?m?�?�? �?�?�? OO$O�?HO 3OlOWO|O�O����O ӯ�O�O�O!__E_3_ i_W_�_{_�_�_�_�_ �_o�_/oo?oAoSo �owo�o�o�o�o�o�o +O=s�E� ��Y����� 9�'�]�K�m������� u�Ǐɏۏ���5�G� Y�k�%���}�����ß şן���1��U�C� y�g�������ӯ���� ��	�+�-�?�u�c� ���������Ͽ�� �/�A�S�����qϓ� �ϧ��������%�7� I�[���mߣߑ߳� �����߷��3�!�W� E�{�i������� ������A�/�e�S� u������������� ��+aO�s ��e�����' K9o]�� �����#//G/ 5/k/}/�/�/[/�/�/ �/�/�/??C?1?g? U?�?y?�?�?�?�?�? 	O�?-OOQO?OaO�O uO�O�O�O�O�O�O_ __M_�e_w_�_3_ �_�_�_�_�_oo7o %o[omoo�oOo�o�o �o�o�o!3�o�o iW�{���� ���/��S�A�w� e�������я����� ��=�+�M�s�a��� ������ߟ�_	�� �_ן]�K���o����� ��ۯɯ���#��� Y�G�}�k�����ſ׿ ��������U�C� y�gϝϋ��ϯ����� ���	�?�-�c�Q�s� u߇߽߫�������� )��9�_�M����/� ���i������%�� I�7�m�[��������� ����������EW i{5����� ���A/eS �w�����/ �+//O/=/_/a/s/ �/�/�/�/�/�/?'? ��??Q?c??�?�?�? �?�?�?�?O�?5OGO YOkO)O�O}O�O�O�O��N  �@S �V_R�$TB�JOP_GRP �2,�E��  ?�V	�-R4S.;\��@�|u0{SPU �>��UT �@�@LR	 �C�� �Vf  C����ULQLQ>�s33�U�R����U��Y?�@=�ZC]��P��ͥR��P  B��W$o/g�C��@g�dDwb�^���ee�ao�P&ff�e=��7LC/kaB �o�o�P��P�efb_-C�p��^g`��d�o�PL�Pt<߿eVC\  �Q@��'p�`�  A��oL`�_wC�?BrD�S�^�]��_�S�`<PB���P�anaa`C�;�`L�w�aQox�p�x�p:��X�B$'tMP@�PCH S��n���=�P��x��trd<M�gE� 2pb����X�	�� 1��)�W���c���� ��������󟭟7�@Q�;�I�w���;d�V�ɡ�U	V3.�00RScr35QT*�QT�A��� E�'E��i�FV#F�"wqF>��F�Z� Fv�RF��~MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
�D���E'
EMK�E���E�ɑ�E�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F��v�F�u�<#�
/<t���ٵ=��_��V ��R�p�V9� ]ES/TPARtp�HFP�*SHR\�ABLE� 1/;[%�SDG�� �W�G�GȡG� WQG�	G�
�G�GȖ�QG��G�G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ�H����w�S]�CS !� ������������ �&�8�J�\�n����� �������� ]\�`�� 	��(�:�����
���.�@�w�NUM�  �EEQ��P	P ۰ܰw�_?CFG 0���)r-PIMEBF_�TTb��CSo�,V�ERڳ-B,R� 11;[ 8$��R�@� �@&  ������ �//)/;/M/_/q/ �/�/�/�/�/?�/? J?%?7?M?[?m?>�@ �?�?�?�?�?�?�?O #O5OGOYOkO}O�O�O �O�O�O�O�O__1_�C_U_g_y_�_�_l_��Y@cY�MI__CHAN8 c} cDBGLV���:cX�	`ETHERAD ?f�\`��?�_uox�oQ�	`ROUTV!	
!�d�o�l?SNMASKQhc>ba255.uߣ�'9ߣY�OOL�OFS_DIb���U;iORQCTROL 2		���~T�����#� 5�G�Y�k�}������� ŏ׏�����.���R�V�PE_DET�AI/h|zPGL_�CONFIG �8�	���/c�ell/$CID?$/grp1V�̟ ޟ����Ӏ�o?� Q�c�u�����(���ϯ ������;�M�_� q�����$�6�˿ݿ� ��%ϴ�I�[�m�� �ϣ�2���������� !߰���W�i�{ߍߟ���%}F�������@/�A�C�i�H�E� �����������?�� .�@�R�d�v������ ����������*< N`r���� ���&8J\ n��!���� �/�4/F/X/j/|/ �//�/�/�/�/�/? ?�/B?T?f?x?�?�? +?�?�?�?�?OO�? >OPObOtO�O�O�O����User �View ��}}�1234567890�O�O�O_#_5_�=T�P��]_���I2 �I:O�_�_�_�_�_�_X_j_�B3�_GoYoko@}o�o�o o�op^46o �o1CU�ovp^5�o�����	�h*�p^6�c�u�����������ޏp^7 R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3��O�M�_�q��������y  e��Yz���	��-� ?�Q���uχϙ�俽�@��������>��e� 5i��c�u߇ߙ߽߫� d������P�)�;�M� _�q��*�<��i��� ������)���M�_� q�������������� ��<�û��=Oas ��>����* '9K]f�Q� ������/� %/7/I/�m//�/�/ �/�/n<��^/?%? 7?I?[?m?/�?�?�?  ?�?�?�?O!O3O�/ <׹��?O�O�O�O�O �O�?�O_!_lOE_W_@i_{_�_�_FOXG9+_ �_�_oo(o:o�OKo po�o)_�o�o�o�o�o( ��	g�0�oM _q���No�� ��o�%�7�I�[�m� &l�n��Ə؏� ��� ��D�V�h��� ������ԟ柍�g� ڻ}�2�D�V�h�z��� 3���¯ԯ���
�� .�@�R���3uF�鯞� ��¿Կ������.� @ϋ�d�vψϚϬϾ� e�w���U�
��.�@� R�d�ψߚ߬����� ������*���w� ��v�������w� ����c�<�N�`�r� ����=�w��-����� *<��`r� ���������  ��1CU gy�������   -/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O�_!_3_E_W_i_� � 
��(  �>%( 	 y_�_ �_�_�_�_�_o	o+o -o?ouoco�o�o�o�Z* �Q &�J\n��� ���o���9�(� :�L�^�p�������� �܏� ��$�6�}� Z�l�~�ŏ����Ɵ؟ ���C�U�2�D�V��� z�������¯ԯ��� 
��c�@�R�d�v��� ��᯾�п�)��� *�<�N�`ϧ����Ϩ� ���������&�8� �\�n߀��Ϥ߶��� ������E�"�4�F�� j�|�������� ����e�B�T�f�x� ������������+� ,>Pb���� ������( o�^p���� ��� /G$/6/H/ �l/~/�/�/�/�// �/�/?U/2?D?V?h?pz?�?�/�`@ �2��?�?�?�3�7�P���!frh:\t�pgl\robo�ts\m20ia�\cr35ia.xml�?;OMO_OqO��O�O�O�O�O�O�O ���O_(_:_L_^_ p_�_�_�_�_�_�_�O �_o$o6oHoZolo~o �o�o�o�o�o�_�o  2DVhz�� ����o�
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟� ݟ��&�8�J�\�n� ��������ȯߟٯ�� �"�4�F�X�j�|��������Ŀ־�8.1� �?@88�?�ֻ�ֿ�3� 5�G�iϓ�}ϟ��ϳ� �������5��A�k��U�wߡ߿��$TP�GL_OUTPU�T ;�!�! ������� �,�>�P�b�t��� �����������(� :�L�^�p�������������2345678901�������� �"��BTf x��4�����
}$L^p ��,>��� / /$/�2/Z/l/~/�/ �/:/�/�/�/�/? ? �/�/V?h?z?�?�?�? H?�?�?�?
OO.O�? <OdOvO�O�O�ODOVO �O�O__*_<_�OJ_ r_�_�_�_�_R_�_�_ oo&o8o�_�_no�o �o�o�o�o`o�o�o "4F�oT|����\��}���� �0�B�T�e�@�������� ( 	 ��Џ������ <�*�L�N�`������� ��ޟ̟���8�&� \�J���n��������� ȯ���"������� *�X�j�F�����|�¿ Կ��C���ϱ�3�E� #�i�{�忇ϱ�S��� �������/ߙ�S�e� ߉ߛ�y߿���;��� ����=�O�-�s�� �ߩ��]�������� '����]�o������ ������E�����5 G%W}������ g���1�U g	w�{��= O	//�?/Q///u/ �/��/�/_/�/�/�/ �/)?;?�/_?q??�? �?�?�?�?G?�?O�? OIO[O9OO�O�?�O �OiO�O�O�O!_3_�O _i_{__�_�_�_�_��_�R�$TPOF?F_LIM >�op>:��mqb�N_SV`  �l�jP_MON7 <6�dop�op2l�aSTRTCHK =6��f� bVTCO�MPAT-h�afVWVAR >Mm��h1d �o ��oop`ba_D�EFPROG �%|j%ZERO ZUZAUN	��j_DISPLA�Y`|n"rINST�_MSK  t|� ^zINUSE9R�odtLCK�|}{QUICKMEJp��"rSCRE�p�6��btps�cdt�q��b*�_�.�ST�jiRAC�E_CFG ?�Mi�d`	�d
�?�u�HNL 2E@|i����k r ͏ߏ���'�9�K��]�w�ITEM 2�A�� �%$1�23456789y0����  =<��xП��  !���p��=��c��^� ���������.��� R��v�"�H�ί��Я ������*�ֿ��� r�2ϖ�����4�޿�� ����&���J�\�n��� @ߤ�d�v��ς���� ��4���X��*��@� �����ߨ����� ��T���x������ l��������,�>�P� ������FX��d�� ����:�p "��o���� �F6HZt~� �N/t/�/��// / 2/�/V/?(?:?�/F? �/�/�/j?�??�?�? R?�?v?�?QO�?lO�? �O�OO�O*O|O_`O  _�O0_V_h_�Ot_�O __�_8_�_
oo�_ @o�_�_�_Lodo�_�o �o4o�oXojo3�oN �or��o���s�S�B���z�g  h��z ��C�:y
 P�v�]�����UD1:\������qR_GR�P 1C��� 	 @Cp����$��H�6�l�Z�� |�����f���˟���ڕ?�  
��� <�*�`�N���r����� ��ޯ̯��&��J�8�Z���	�u����~�sSCB 2D� �����(��:�L�^�pς��|V_�CONFIG �E���@����ϖ�O�UTPUT F<�������6� H�Z�l�~ߐߢߴ��� ���������#�6�H� Z�l�~�������� ������2�D�V�h� z��������������� 
�.@Rdv� ������ )<N`r��� ����//%8/ J/\/n/�/�/�/�/�/ �/�/�/?!/4?F?X? j?|?�?�?�?�?�?�? �?OO/?BOTOfOxO �O�O�O�O�O�O�O_ _+O>_P_b_t_�_�_ �_�_�_�_�_oo'_ :oLo^opo�o�o�o�o �o�o�o $���� !�bt����� ����(�:�-o^� p���������ʏ܏�  ��$�6�G�Z�l�~� ������Ɵ؟����  �2�D�U�h�z����� ��¯ԯ���
��.� @�Q�d�v��������� п�����*�<�M� `�rτϖϨϺ����� ����&�8�J�[�n� �ߒߤ߶��������� �"�4�F�W�j�|�� ������������� 0�B�S�f�x������� ��������,> Pa�t����� ��(:L/x���k}g V�K���// &/8/J/\/n/�/�/�/ W�/�/�/�/?"?4? F?X?j?|?�?�?�?�/ �?�?�?OO0OBOTO fOxO�O�O�O�?�O�O �O__,_>_P_b_t_ �_�_�_�O�_�_�_o o(o:oLo^opo�o�o �o�o�_�o�o $ 6HZl~��� �o���� �2�D� V�h�z��������ԏ ���
��.�@�R�d� v���������Ϗ��� ��*�<�N�`�r��� ������˟ޯ��� &�8�J�\�n����������Ż�$TX_S�CREEN 1G�g�}ipnl/��gen.htmſ��*�<�N�`Ͻ�Panel se7tupd�}�dϥ� �����������ω� 6�H�Z�l�~ߐ�ߴ� +�������� �2�� ��h�z������9� g�]�
��.�@�R�d� �������������� }���<N`r� �;1�� &8�\�������QȾUAL�RM_MSG ?5��� �Ȫ -/?/p/c/�/�/�/�/ �/�/�/??6?)?Z?~%SEV  -��6"ECFG� I�� � ȥ@�  A��1   B�Ȥ
 [?ϣ��?OO %O7OIO[OmOO�O�O��G�1GRP 2J�; 0Ȧ	 ��?�O I_BBL�_NOTE K��:T���lϢ�ѡ�0RD_EFPRO %+ (%N?u_Ѡc_ �_�_�_�_�_�_o�_�o>o)oboMo�o\I�NUSER  �R]�O�oI_MENHIST 1L�9  ( _P���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1�oCUgy3�)
13/������p1��ue�dit(rTISC�HZUZAUN,A1�GK�]�o����|o ����ʏ܏� ���$� 6�H�Z�l�~������ Ɵ؟�������2�D� V�h�z������¯ԯ ���
��h9Rq��B� T�f�x���������ҿ ����ϩ�>�P�b� tφϘ�'�9������� ��(߷�L�^�p߂� �ߦ�5������� �� $����Z�l�~��� ��C�������� �2� �/�h�z��������� ������
.@�� dv�����_ �*<N�r �����[�/ /&/8/J/\/��/�/ �/�/�/�/i/�/?"? 4?F?X?C�U��?�?�? �?�?�?�/OO0OBO TOfO�?�O�O�O�O�O �O�O�O_,_>_P_b_ t__�_�_�_�_�_�_ �_o(o:oLo^opo�o o�o�o�o�o�o �o $6HZl~i?{? ������2� D�V�h�z����-� ԏ���
����@�R� d�v�����)���П� ��������N�`�r� ������7�̯ޯ�� �&���J�\�n�����������$UI_�PANEDATA 1N���ڱ�  	��}/frh/�cgtp/wid�edev.stm����%�7�I�Y�)Gpriρ�@�}����ϻ�������� ) �)��M�4�q߃�j� �ߎ����������%��7��[�7����     2ƓϘ��� ������E����:�L� ^�p������������ ����$H/l ~e������o� ݰܳ7�<N `r����-�� �//&/8/�\/n/ U/�/y/�/�/�/�/�/ ?�/4?F?-?j?Q?�? �?%�?�?�?OO 0O�?TO�xO�O�O�O �O�O�OKO_�O,__ P_b_I_�_m_�_�_�_ �_�_oo�_:o�?�? po�o�o�o�o�oo�o  sO$6HZl~ �o�������  �2��V�=�z���s� ����ԏGoYo�.� @�R�d�v�ɏ���� П������<�N� 5�r�Y�������̯�� �ׯ�&��J�1�n� ������ȿڿ��� �c�4ϧ�X�j�|ώ� �ϲ���+�������� 0�B�)�f�Mߊߜ߃� �ߧ��������� P�b�t�������� ��S���(�:�L�^� ���i�����������  ��6ZlS`�w�'�9�}��@�"4FX)� }��l����� /j'//K/2/D/�/ h/�/�/�/�/�/�/�/�#?5??Y?��C�=���$UI_POST�YPE  C��� 	 �e?�?�2QUICK�MEN  �;��?�?�0RESTO�RE 1OC��  ��L?��6OCC1O��m aO�O�O�O�O�OuO�O __,_>_�Ob_t_�_ �_�_UO�_�_�_M_o (o:oLo^oo�o�o�o �o�o�oo $6 H�_Ugy�o�� ���� �2�D�V� h��������ԏ ����w�)�R�d�v� ����=���П���� ��*�<�N�`�r��� �����ޯ���&� ɯJ�\�n�������G��ȿڿ�����7SC�RE�0?�=�u1sc+@uU2K�3K�4K�5Kĕ6K�7K�8K��2U�SER-�2�D�ksTMì�3��4��5�ĕ6��7��8���0N�DO_CFG �P�;� ��0PDA�TE ����None�2��_INFO 1QC�@��10%�[��� Iߊ�m߮��ߣ����� �����>�P�3�t���i���<-�OFFS_ET T�=�� ��$@������1�^� U�g������������ ����$-ZQcu���?�
�����UFRAME  �����*�RTO?L_ABRT	(��!ENB*GR�P 1UI�1Cz  A��~��@~���������0UJ�9MSK  M@�;-N%8�%��/��2VCCM��V��ͣ#RG�#Y�9����/����D�BeH�p71C����3711?�C0�$MRf2_�*S��괰	���~XC56 *�?�6�Y��1$�5����A@3C��. 	��8�?��OO KOx1FOsO�5�51ⴰ_O�O�� B����A2�DWO �O7O_�O8_#_\_G_ �_k_}_�__�_�_�_��_"o�OFoXo�%TCC�#`mI1�i���u��� GFS�»2aZ; �| 2�345678901�o�b�����o@��!5a�4BwB�`�56 311:�o=L�Br5v1�1~1�2 ��}/��o�a��# �GYk}�p�� �����ُ�1�C� U�6�H���5�~���ߏ����	���4�dSEGLEC)M!v1b3��VIRTSYN�C�� ���%�SIONTMOU�������F��#b�U��U�(�u FR:\�H�\�A\�� ��� MC��L�OG��   U�D1��EX����'� B@ �����̡m��̡  �OBCL�1�H�� �  =	 �1- n6 � -������[�,xS�A�`=��͗���ˢ��TRA�IN⯞b�a1l�
�0d�$j�T2cZ; (aE2ϖ�i�� ;�)�_�M�g�qσϕ� ���������	��F�STAT dmB~2@�zߌ�*j$i�\���_GE�#eZ;7�`0�
� 0}2��HOMIN� �fU��U�� ~�����БC�g��X���JMPERR� 2gZ;
   ��*jl�V�7������ ��������
��2�@��q�d�v�B�_ߠREr� hWޠ$LEX�ԹiZ;�a1-e��V�MPHASE  �5��c&��!OF�F/�F�P2n�jJ�0�㜳E1�@��0ϒE1!1?s#33�����ak/�@kxk䜣!W�m[�䦲�[����o3;� [ i{���� /�O�?/M/_/q/ ��/��//�/'/9/ �/=?7?I?s?�/�?�/ �/�?�??Om?O%O 3OEO�?�?�O�?�O�O �?�O�O�O__gO\_ �OE_�O�_�O�O/_�_ �_�_oQ_Fou_�_|o �o�_�oo�o�o�o�o ;oMo?qof-�oI �����7� [P��������� ˏ��!�3�(�:�i��[�ŏg�}������TD_FILTEW��n�� �ֲ:���@���+�=�O�a� s���������֯� ����0�B�T�f�x����SHIFTME�NU 1o[�<��%��ֿ����ڿ� ���I� �2��V�h� ���Ϟϰ�������3��
�	LIVE/�SNAP'�vs�fliv��E�����ION * U<b�h�menu~߃������ߣ���p����	����E�.ォ50�s�P�@� �Z�AɠB8z�z�!�}��x�~�P��� ���MERb���<�0���kMO��q���z��WAITDINE�ND������O9K1�OUT���SD��TIM����o�G���#����C���b������RELEASE������TM�������_�ACT[�����_DATA r�%L����xRD�ISb�E�$X�VR�s���$Z�ABC_GRP �1t�Q�,#�r0�2���ZIP�u'�&����[�MPCF_G 1	v�Q�0�/� �w�ɤ� 	|�Z/  85�`�/�/H/�/l$?��+ �/�/�/?�/�/???|r?�?  �D0 �?�?�?�?�?�;����x�]hYLI�ND֑y� ���� ,(  * VOgM.�SO�OwO�O�M i?�O�O^PO1_ �OU_<_N_�_�O�_�_ �__�_�_x_-ooQo�8o�_�o�oY&#2z� ���oC� e?a?>N|�oq��햋qA�$DSPH�ERE 2{6M� �_�;o���!�io |W�i��_��,��Ï ���Ώ@��/�v��� e�؏��p�����������ZZ�� � N