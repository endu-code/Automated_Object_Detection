��   !�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����CCPTP_�CFG_T  �P '$DAT�A_PATH �!$OUTPU�T>PART_N�AMEC $ED�GE\!$CLR�_VDB_BUF�  $x_S�IZ 9VER~�DEV_ID��H �VIS_REyS���P_DT��POS_OFS_�ENB�TAR_�D� �DEBUG�_MOD` � MAX_FC_PN���CUVS�EGLAP
TPP_� 
X
fH�f�Ac� L��CNS� �JUM�P_LEN_t$CURV�V�5T�T�MAT�?ABOVE_���$TOL_WP�R_CHH! EXP�SA "��ERR_H�� __LONG1L*2L&/REALY!l&g!��$s ASS ? ����!���Z��Z� � SIO�N�(  ��5�!IRTU�AL�/�!'2 �(Z�!FR:\) �:\����!UD1:?���!G?38D?q?��� ��� ��6��N�0u0  [�3 d�0г8���0  ?���BH  @�1�  >�0�2��3�?C