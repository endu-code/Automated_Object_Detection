��   ʇ�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DCSS_C�PC_T� �$COMMENT� $ENA�BLE 6 MO�DJGRP_NU�MKL\  ?$UFRM\] ?_VTX 6 � �  $Y�Z�1K $Z2�STOP_TYPK�DSBIO�ID�XKENBL_C�ALMD�USE_PREDIC? � &S. �c 8J\TC�~u
SPD_LI_0���SOL�&|Y0  � 1CHG_SIZO$APGESDIS��G�!C����Jp 	�J�� &�"��))$'2_SE��� XPANIN�  �STAT�/ D $F�P_BASE �$_ K�$!� �&_V�.H�#0:g%J- ��ZAXS\UPR�JLW7Se���&� | 
 �/�/�/D&?8?zh$�ELEM/ Tc ��2�"NOG<�0�3UTOOi�2�HAD�� $D7ATA"g%e�0  @@p:�0 _2 
&Pp%' � p!U*n   �FS�Cz�B�� �B(�F�D(�R|UC�DROBOT�H��CqBo�E�F$�CUR_2Rh$SwETU�	 l� ��P_MGN�I?NP_ASS�0 "@�� �3�8B7gP@U��^V�Sp!�h$T1�
`B|8�8�TM 0 �6P�+ Ke�1VRCFY�8
dD5F1� ��W��1$R��8SPH/ (�{ �CA�CA�CA3�BOX/ 8 �0������b'o�EjTUIR�0 � ,{ FR`ER��02 $�` ��a_S�b��gZN/ 0 �{9F0� -a0rZ	_0�_0�u0  @Q�Yv	�o:o� �$$CLLP ? ����q���Q��Q�pVERSwION�xZ0��5�qIRTU�AL��q' 2 ��xQ   ��Double �Parts Si�de�� �0�p����#PDM@DM�-�N��  ��@k����� W����0��q`��/�A�S�f D��|
�y�DJ@ D�p+������򫏽� r��a�W�u����ٟ �Z��~���Ɵ��F� {������� �2�h��� ��/���S�¯ԯ� ��
���ѿ@���d�v� ��=Ϭ�a�s�⿗ς� �*���N��߄�%� Kߺ��ρ��ϥ߷�N� 8���\�n�#��G�Y� k��ߏ������4��� ���|�1����9��� w��������B�T��� x�
?Q��u���� ,����b� ��_���� (:L/p%/7/� [/F/���//�/�/ H/�/?~/�/E?�/i? {??�/�? ?2?�?V? OO/O�?SO�?�?�O �?�O�O�O@O�OdOvO �O�O;_a_s_�O�__ _N_<_�_oo�_9o �_�_�_�opo�o�o&o �oJo\ono#�oGY �o}�o�o�4� �j�
���g�� �������ӏB�T�	� x�-�?�֏��u���� ���ϟ��b���� ��M���q�������� (�:���^���%�7��� [�ʯܯ� ���ǿٿ H���l�~���E�4�i��{���$DCSS�_CSC 2�!���Q  D�������*� �������A��S�4� ��X߭�|��ߠ����� �����<�a�0�B�� f���������'� ��K��o�>�P���t� ����������5 Y(}L^����'ɘ�GRP 2N�� ��,�	Z� ?*cN�r�� ����/)//M/ 8/q/\/�/�/�/�/�/ �/?�/�/7?"?[?F? ?j?�?�?�?�?�?�? �?!OOEO0OiOTO�O �O�O|O�O�O�O�O�O /__S_>_w_�_�_f_ �_�_�_�_�_oo=o (oaoso�oPo�o�o�o �o�o�o�o'K] o:�~��������5��_GS?TAT 2��1��,8����ô?5�|���?�  5*����Ҵ������}����D���bH^��z$�8t��;�.���/����Z�w0�I����3��4�����C-å�t�/�M'B���|�͈��X[D1'U�D�N䏖�������M��r�4��r������DK��D&+�����Ѐ/��u4�D��ZBbE� T�.�@���w�����ȑ ������ �F�X�6� |�������+Ű�%�ĕ ���ԯ� �
��>� @�R�t�������Կ� ���`���D�V�4�z� �Ϧ�࿶ϼ������� ��"��.�X�B�dߎ� xߊ��߮�l����߀<�N�,�r��b�ؑ��?���Ǚg��8(��� �,�Ǫ�4� ����Dr*@�m�aDC������z�1�/��ԀUؑ�����ԁC���������~��8�z��?�D��<:z?������B��Y�ſ"DE:ĕ=�����|�@?|�:z�+�����ު�|��:z(�=���B��a�נ�oDj��H�|�h�=�p�����A��bSD\�������2���m:����(C��=4��ſ&ؑ�� �����h�:L*p �`��������� �$N8J� n�����/� 2/D/�h/z/X/�/�/ �/�//�/?�/? .?0?B?d?�?x?�?�? �?�?�? /*O<O�/`O rOPO�O�O�O��
�� �������"�4�F�X� j�|������������� �O�O�Ojo�OZo�o �o�o�o�o�/O�? H2T~h�� ����� �
��o b�t�R�������Ώ�� �o4�
���@�*�L� v�`�r�������ʟ̟ ޟ �*���Z�l����� ����Ưد�O(o:o�O 
__._@_R_d_�_�_ �_���_�_�_�_oo ��No�Ϛϴ����� ��������8�B�� N�x�b߄߮ߘߺ��� ������&�P�:�� ���ς��������� *�d�:�@�F�p�Z�|� �������������� H2���z� ����X�j�(� :�L�^�p��������� ʿܿ� ��$�6�  2D~ϸ/�/��/ ? �/$?6?�F`?j\? ~?�?�?�?�?�?�?O �? OJO4OVO�Or�O �O?�O�O�O_._H? Z?�Oj_pOv_�_�_�_ �_�_�_o�_oBo,o Noxobo@_�o_�o�o �o&8v/�/�/X j|������ �//h/B/T/f/P bt���؏�0� �T�f�L_�o���o�� Ɵ��������� .�P�z�d������o� �D��(��L�^�x� ����Ư��������ܿ ���<�&�H�r�\� ~Ϩ�ί����<��� � ��0�V�4ߦ���ʏ� �������� *�<�N�`�r������ ��̏F��*��N�`� >�����|��������� ����,8bL ^�����v� " FX6|��� �������$/ / /B/D/V/x/�/�/ �/�/�??l>?P? .?t?�?p�����߸� ������ ��\�6�H� Z�l�~������? �?��?H_�?X_~_\_ n_�_�_��/�_�/�_ &oo2o\oFoho�o|o �o�o�o�o�o�o�_@ R0v�f���_ ��o���*�T� >�`���t��������� ޏ���8�J�(�n����^������u�$DC�SS_JPC 2��uQ ( D���#�� �@�G��(� }�L�^�p�ů��ӯ�� �ܯ1� �U�$�6�x� ��l�~�ӿ����ƿ� �?��c�2χ�Vϫ� zό��ϰ�����)��� 7��q�@ߕ�d߹߈� ���������7��� *��N��r������ �������E��&�8� ��\������������� ����@e4F� j|����+ �OsBT�x ������9// ]/,/�/P/b/�/�/�/ �/�/�/�/�/G??k? :?�?^?�?�?�?�?�? O�?�? OUO$OcO"�*ԕSݐ�@NO�O rODO�O�O_�O?__ $_u_H_Z_l_�_�_�_ �_�_�_�_;oo o^o �oVoho�o�o�o�o �o�o7
E.R d������� 3���*�{�N�`��� Ï������̏���A� �&�w�J���n����� ����ȟڟ�=��"� s�F�X�j�������ޯ �֯�9��]�0��� T�f�����ſ����ҿ �5���,�}�P�b� �φϘϪ�������� C��(�y�Lߝ�p��� �ߦ��������?���$�u�H�Z�HMOD�EL 2�K�xp�e�
 <��c���  g� ��l�����R�)� ;�M�_�q��������� ����%7� [m������ �a�J��!�	 w����/�� B//+/=/O/a/s/�/ �/�/�/�/�/�/?? '?t?K?]?�?EW�? �?O?�?�?LO#O5O �OYOkO�O�O�O�O _ �O�O6___l_C_U_ g_�_�_�_�_�_�_ o �?�?�?oo�_couo �o�o�o�o�o�o�o )vM_��� ����*���`� 7�I�[�1o��Uo���� k�ُ�8��!�n�E� W�i�{������ß՟ "�����/�A�S��� w���֯����ѯ��0� ˏ���x�O�a����� ��俻�Ϳ߿,��� b�9�KϘ�oρϓ��� ���������L�#�5� G����A�o߁����� ��$�����1�C�U� ��y����������� ��	�V�-�?���c�u� �������������� ��d;M�q�� ����N% 7I[m��� /���/!/3/	 �/-[/m/�/�/�/? �/�/?X?/?A?�?e? w?�?�?�?�?O�?�? BOO+OxOOOaOsO�O �O�O/�/�/�O�OP_ �O9_K_]_o_�_�_�_ �_o�_�_�_o#o5o �oYoko�o�o�o�o�o �o�o6l__ GY�A���� �D��-�z�Q�c�u� ��������Ϗ�.�� �)�;�M�_������� �}���ϟ<���%� 7���[�m�������� ǯٯ�8��!�n�E� W���{������ÿտ "����X����E� W�-ϛϭ�������0� ��+�=�O�a߮߅� ���߻��������� b�9�K��o���i� ��ϻ�����#�p� G�Y���}��������� ��$��Z1CU gy����� �	��h�1C� �����/�/ /d/;/M/�/q/�/�/ �/�/�/?�/?N?%? 7?�?[?m??U�?y �?�?&O�?O\O3OEO WOiO{O�O�O�O�O_ �O�O__/_A_�_e_ w_�_�_�_�_�_�_�_��:�$DCSS_�PSTAT ����_aQ    po6~j no (�o�oh�o�o�o | �`�``q�`7o0B�9�*c_elpa�~PdSETUP 	_i'B�"d�3�1�t�KiT1SC 2
4�zp�1Cz�3���+��uCP R�|��0D�?v��� �?����Џ����� �<�N�`�/�����e� ��̟ޟ����&��� J�\�n�=��������� گ��>d�!�3���W� i�{�J�����ÿ��� ���ڿ/�A��"�w� ��XϭϿ��Ϡ���� ���=�O�a�0߅ߗ� �������f���'� ��K�]�o�>���� ���������#�5�� Y�k�}�L��������� ������1C�߼� y������ 	�?Qc2� �hz���// )/�M/_/q/@/�/�/ �/�/�/�/Vh%?7? �/[?m??N?�?�?�? �?�?�?O�?3OEOO &O{O�O\O�O�O�O�O �O__�OA_S_e_4_ �_�_??�_�_j_o o+o�_OoaosoBo�o �o�o�o�o�o�o�o' 9]o�P�� ������5�G� �_�_}������ŏ׏ �������C�U�g� 6�����l�~�ӟ埴� 	��-���Q�c�u�D� ����������Z�l� )�;�¯_�q���R��� ��˿������7� I��*�ϑ�`ϵ��� �Ϩ����!���E�W��i�8ߍߟ߯��$D�CSS_TCPM�AP  ������Q W@ z�z�zЩz���z�z��z�z�	�  �z�z�z�z��z�z�z�z��z�z�z�z�Rz�z�z�z�z�Uz�z�z�z�U z�!z�"z�#z�U$z�%z�&z�'z�U(z�)z�*z�+z�U,z�-z�.z�/z�U0z�1z�2z�3z�U4z�5z�6z�7z�U8z�9z�:z�;z�U<z�=z�>z�?z��@��UIRO 2]����� � ��0�B�T�f�x��� ������������,>Py��y� ������	 -?Qcu��� ��Z�~�)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? �?
/�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�Or?_���UIZN 2.��	 �����L_ ^_p_u�G_�_�_�_�_ �_�_o�_,o>oPoo to�o�ogo�o�o�o�o �o(�oL^p� E����� �� �6�H�Z�)�~����� e�Ə؏ꏹ�� �2� ��V�h�z�I����� ԟ����
�ٟ.�@�R��_��UFRM R.����8}ߪ� ��{���ͯ�(�� L�^�9�����o���ʿ ��� �ۿ$�6��G� l�~ϕ��ϴ�S����� ��� ���D�V�1�z� ��g߰��ߝ�����
� ��.�@��d�v�Ϛ� ��K���������� <�N�)�_�����q��� ��������&8 \n���C�� ��"�FX3 |�i����� �/0//T/f/}t/ �/�/�/�/�/�/?? �/>?P?+?t?�?a?�? �?�?�?�?�?O(OO LO^Ou/�/�O�OEO�O �O�O __�O6_H_#_ l_~_Y_�_�_�_�_�_ �_�_ o2ooVohoO �o�o=o�o�o�o�o
 �o.@dvQ� �������*� �N�`�wo����5��� ̏�����ݏ�8�J� %�n���[�������ڟ �ǟ�"���F�X�2�