��   m�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING,��<$1_8k  �FMS*�t *v M_LIF��u,(8*x��M(DSTB0+_0>*_���*#�z&+CL_TIM>�PCCOMi��FBk M� �MAL_�EC�S��P!Q%XO �$PS� �TI����%�"r $D�TY?R. l*1E�ND14�$1�ACST1#4V22\93\9�4\95\96\6_O3VR\6� GA[7�2 h7�2u7�2�7�2�7�2ޜ8FRMZ\6DE��DX\6CURL� HSZ27Fh1DG u1DG�1DG�1DG�1DC�NA!1?( �sPL� + ���STA23TRQ_�M��/@K"�FSUX�JY�JZ�II�JuI�JI�D �$U1�SS  ����6Q����+PV�ERSI� 4W  �5GQ?IRTUAL3_EQ�' 1 TX W ��(P���_�_�_�Vm���څ �!� ���~����������R?����?��J�B�y4���=�t��7�Q��]�����V���u������?�� ��_�P�eygwe�YAQ�o�^A����O ���b I ������o�o�_�l/VSet�$�w�gAP�B�w�un�Q�� Su���}g`� ��`���	 j�����& ~�����j��b%���d�o#�5�G���=gL��R�y�?�z���@�����я��� ��+�=�O�a�s���� rU������ޟ:T  2��!�3� E�W�i�{���������<��ۯ����#�5��G�Y�k�}���������$$ 1�\��aP4DeJ�q��J�kpT�I��QӺN�=� �kD�EJ���:Ha�@��J`BB��@G{(�mA��1����mB�@kB�����`��C�+���Pk��.dP�o�Ϙ�ϸ��+�=ϟ���M�x���2ߡ�V�A�z���� @P�� P�֠՞՞� ����{Ђ�K�}g�L��3L�X�������L��c�MZQ�MZ�R<MZS�MZ�Z��3�8��H�L�VM�]+N�Rxq��td ���t�������6Q�Q� ������8N�S$T�i���i����/U ���� ��� x�
� x���������NQ���Q�sQ�WQ�BM�C��T�C���C����������E���������������������%����^��p��C���C�F�C��4�C���C�������� �6�g�� �7 �4�7 m�t ��ZN �X� ��W �Ts ��1�5���&N� �s�W �/4 �4� �59��m9������{��M��Q��� ��r�N�a�,a�$a� �2��ړ����� ���v�c+�{��M��*M��M��M��M�I����ѡ�š����}� t�� �0q� 1� �1�L 1ح��ρu��EA���@��s�����������������z���N����M���7��9��O�K�͋ w�3���n	 1	 i	 �� �Ġ��1g����F Av���q�����#���+��&��8��'H��>�HdUc

e�AIHJ��`KT��k}+����1sP����x��wbsP��E�Q���`h�sP�td��8f�������>� 2  ��?S�	-��sewasP!R?PO�sP������9��������l>�����h�i�A�s�sP좩�>����� �_����{� ⩀a��H楄��ssPU�bsP�sP�sP����(����������sPd��ͭM��AQ����4-8�ԵP�Ǡ_� =��WSsP��эi&F.�'ce�+�/`,�/�$����?�?���*���Ix�ڭD�@�^�0�g�0p�D��=��.�Ħ^��ħ��0��0�?������&J���L��.c��/m�@�z�0U��06�0G�0P�0�Y�?�s��0��?�t_?�.k�����?-���?-��?-���?-�x?����@��?����?)�?�~��?���?�q`�!@�?�r")@�z)@���z�w9@���z��������b?��>����I.��\�ž�v�u��l��ſ���]�2����!�{.��z�_��z�;y@�y@y�9@��@?���@���BA�=�_�@K��@5�@�D�@N=%��>�y�">�w�ޠ�@Gh�@_�@?�E�@ߍ@�ԍ@ʍ@�5Bh��b�hΪ�@���"�V��>�����,���m���;B���f���/?���?��׫�M?��:E�i�_��hճ�h�9�h�W�hѻ)P�m��B��B���9Q�ݫ�?��K��Jvh��Ju�MP}MP8?�����i���C͆?+��Wu�9P!5P
5PU5P 5P9P�� �,($not a� program�|?���_�_�_�_�_PLACE�_%o�_Io0hZERXmoTofo��o�o�o�o�o�o4dFRAM�o,7oP7�I�($A�q_POSPIC���xA��_q��� �#�`�G���k�}���x��ޏ��PLCLų��� �D1�ѐ?� � �>���?C��q�T�m�x�c� �������������� �>�P�