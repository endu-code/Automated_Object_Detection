��   :�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP �   �$8 A~O  ���z�����o VER�SIONw�  �5�IRTUALw�'�DEF\ � � �� ���ENA'BLE� �������LIST 1 ��  @!H�,��)���( yL^����� ��-/ /Q/$/u/H/ Z/�/~/�/�/�/�/�/ ?�/:? ?q?D?V?h? �?�?�?�?�?O�?7O 
OOmO@O�OdO�O�O �O�O�O_�O3___ U_<_z_`_�_�_�_�_ �_�_�W