��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER� q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS�	 DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� �DRE-  ? � �0�BB{F S{T� M�D|TRS$STD6XlQCWFA� 7X�QCW��"YV�"eS/ �A7 �  $�@TI�Nd@�0SULگ �R_@ g $}@ SW�@�RO�RR%	� �P�T� �@J�U� �SqFS4DN6
 �2P�0_@�cFOL[d!$�FIL� jjE�P��C�S�aDIG4R_C_SCA��c�INTTHRS�_BIdA�dSMA9L�bCOL�b9G�`� �� ��_IVTIM��$!0B"$S�?0xCCBDDN���-qI2wT2wDE�BUdA\!SCHN�"TOfa0�! �  Q0mr<0V� �;!�r~AUTTUN�� TRQa�uE�40N �qFS3A	XG  � 1eb}t��rI�v Q�agr7 �l �!�3@W�EIGH�q�2 �uS_5QF(�T2�W�A� 	pEsNTERVA�; - Q�� �S!�t�AS0S�$�J-_STA�p QJQg���1(���2��3��W���� �hqx��"COG_X��Y�Z�ҁCM��p?�p�܂RSLT�4��D��(D��	"_�p_�q7 � �~�b#0VR�OUNDCMVPE�RIODA�1PUnU3F2D�'TM1�� �Ƒ_D��G�AMMc1�TR�XI�K�K�K���CLbP�&O00A�DJ�GAu�UP�DB#I%0 ,$M"P30f��� d�:pG p�"��HCD�GV��#GVY��Z�J�DO5�,q��S��$R��E_8@{٣��pAPHBC<��$VF6�P�b�2L��蘨@IL[� ���;���;�d@��RG���NEW_���r�Q}���ڡ�5'OBOA@fY�sW2
/�G<�	����ȴ\��2�E�KP�NUCNPRGOV����@N`d_TW�c,�G�E^!NV2#C�c0@��WTS�TRL_�SKI2!$SJ��Q��NQpGW��J�	"��7 \ ;60FR]b� � CMDC���T�b���TO?��� �5گ���_�Ah 0 '��ALARM�_�*�wTOT6�FRZn l�,!Y 3��X!��m� ��X �Œ`X �ʕ�U#
��2��2
�X#Z���'FIX�8��F�"��IT�`IB�PN�_d��CH�%��_sDFL _�BF2N��ڶ�3����� ��3�"�����ʷ�� ����3��3
��X��DIA����/#B� ���%����� [1��g1�[���Z��#���!���%���$@0�@
p��7F��D�� HA�pU�5�����v�FSIW6 ��2PN@�`R>!��PHMP�`HCK %���>0G�'*#e 1A����pNT��^8H	��HUFRzs�3��A��UgvCa�$�v0Q ���4�@p@p �  sSI0� P��5�IRTU�_��� %SV 2���   �P6>0]@]	Q<�EF@ �o|P�  @p P� �//'/9/�K/U%@pd@p
m h K�/w/�/�/�(��$ ��/� �/�/?.8e" �/?J?\?r?8?�?|? �?�?�?�?�?�?>O4O bOO�OTO�O�OjO|O �O�O�O_�O(__\_ f_�_B_�_�_�_�_ o �_$o�_Ho>oo^b�/��ot��%�/�o�o�k�	MC: 56�78  Afs�dt1 78901234q#5w/  	q 6xzc.Ops�'���j l�o�o��� ������,�5�~DMM �)5�A ��x���𨏺�=���OR 2]	Q� ��m���_� tuB?�)DN�S�4D 
Q�!tY�d�!Ls|�q`rlƈ̀?�l�B����$ ONFIG� �(o� �� �����i!��� 2�,�
Hand g�uide��?�3����  �X���с��ь�g#?�=���A��ύ �������p�ݯ� (��L�7�p�[����m*������ʿ ܿ� ��$�6�H�Z� lɌ��ό��ϰ����Ϡ���
�C�E�I �2Q�(�0�� -�zՀ�Fտ���_`πB����d�C��  ��uq=#׽
_aNnk(��K�����̥@��=e��=D����_a�;����8I�y�_aIt$ �}$F�>���k"����Q�Fۀ3]儢ѯǯ���!�/�``+�����.������_a$�=���(4$����޷�>�E��B<�~w%�_a8E�y�5�;�jA��Ҝ{�Q�>��]�_a?��m��箑����<~u1�?�33����0�:�o����0�@����LSB�� ~uq�ӻ��m��S]���8��� ���t�	eF|���]���
�����n�O�;�.����3��'	�����B���4* 2/�V��%D�DH  *%v�+��^-���
�/��/u/~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?;)�7�?�?�o�?�8Jhq�?�?�zyjG�_FSIW Q��9��O�O �Ou�