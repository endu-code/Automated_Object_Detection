��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����CCSCB_�GRP_T  � � $COM�PMATEXP � 9RIX �  0$IN7NER��P0D_�OFFSETS�hCMPAzCO}FsFS_TYCSBFRAMES � Y IT_T�OL�RANGE_� �r�FTRATIOS�h_H_LIM�D �L�FSOOFST1�
2��  �$$CL�ASS  �S��3����(VERSION0w%�5D?IRTUAL0B�' 2 Q� �<  0 -��S��� ���  a����&�H��ٸ����� ���/��� ��B�,��4 @�=  ��D W!o%k!C@ %3 �1 �� BpI'Z/�/�-