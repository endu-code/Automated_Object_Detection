��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  /�  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81F3�K2> �! � �$SOFT�T�_IDk2TOTAoL_EQs $�0�0NO�2U SPI�_INDE]�5X�k2SCREEN_�(4_2SIGE0�_?q;�0PK_F�I� 	$TH{KYGPANE�4� � DUMMYE1dDDd!OE4LA�� R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B!SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C?CFS_UT~p0 "�1�3�#�ؗ`qX"�}R0  4F OIMCM�`O#S�` ��upi �_�p�EBA9!���M/� h�pIMPEE_F�N��N��0�@O��r�D_�~��n�Dy�F� dCCq_�r0  T� '��'�DI�n0"���p�P�$�I������F�t X� GRP0��=M=qNFLI�7��0UIRE��$g"~� SWITCH5��AX_N�PSs"C�F_LIM�� � �0EED���!��qP�t�`PJz_dVЦMODEh��.Z`�PӺ�ELBOF� ������p@� ���3���� FB�/��0�>�G�� �� WARNM��`/��qP��n�N�ST� COR-�0bFLTRh�TR�AT�PT1�� $ACC1a��N ��r$ORI�o"V��RT�P_S� C�HG�0I��rT(2��1�I��T�I1���� x pi#�Q��HDRBQJ; CQ�2L�3L�U4L�5L�6L�7L�U8L�9s!��O`S <F +�=�O�x�#92��LLECy�}"MULTI�b@�"N��1�!���0T��w �STY�"�R`�=l�)2`��8��*�`T  |� �&$��۱m��P�̱��UTO���E��EXT����ÁB���"G2� (䈴![0������<�b+�� "D"���ŽQ��H<煰kcl�9�#���1��ÂM�ԽP���" '�3�$ �L� E���P<��`A�$JOBn�T����l�TRIG3�% dK�������<���\h��+�Y���_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`�0Z���0��P_�P��n@ ( @F RO.���&�t�IT�c�NOM�
����S��`T)w@���Z�1P�d���RA�0��p2b"����
$T��.��MD3�T��`QU31���p(5!HGb��T1�*E�7��c�KAb�WAb�cA4#Y�NT���PDBG�D�� *(��PU�t@X��W���AX���a��eTAI^cB�UF��0!+ g� 7n�PIW��*5 P�7M�8M�9
0�6F�7SIMsQS@>KEE�3PATn�^�a" 2`#��"�L64FIX!, ���!d��D�12Bus=CCI�:FgPCH�P:BAD렀aHCEhAOGhA]HW�_�0>�0_h@�f�Ak� ��F�q\'M`#�"�:DE3�- l�p3G@��@FSOES]FgH�BSU�IBS9WC��.� ` ��MARqG쀳��FACLp�SLEWxQhe�ӿ��MC��/�\pSM_JBM����QYC	g�ex��R�0 ā��CHN-�MP�#$G� Jg�_� #���1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�f�JR���rSEGF�R�PIO� ST�RT��N��cPV5���!41�r��
r�>İ�b�B�O�2` +�[���,q E`&�,q`y�Ԣ}t���yaSIZ%���t��vT�s� �z�y,qRSINF}Oбc��@�k��`��`�`L��8� T`7�CRCf�ԣCC/�9��`a�uah�ub'�MIN��uaD�s�#�G�D�YC��C �����e�q0��� �SEV�q�F�_�eF��N3�s�ah��X�a+p,5!�#1��!VSCA?� A䕖s1�"!3 � �`F/k��_�U��g��]���C�� a�s��R>�4� �����N����5a�R�HA;NC��$LG��P�6f1$+@NDP�t�AR5@N^��a�q���c��ME�18���}0f��RAө�AZ �𨵰�%O��FCT K��s`"�S�PFADIJ�OJ�ʠ� ʠ���<���Ր��qGI�p�BMP�dp�p�Dba��AES�@�	�K�W_��BAS��� �G�5  zM�I�T�CSX[@�@�!62�	$X����T9�{sC��N��`�a~P_HEIG9Hs1;�WID�0�aVT ACϰ�1�A�Pl�<���EXP�g���|��CU�0M�MENU��7�T[IT,AE�%)��a2��a��8 P,� a�ED�E.`��wPDT��REM.���AUTH_KEGY  ������ ��b�O	�.a}1ERR9LH� �9 \� �q�-�OR�DB�_IDx�@l �PUN_O��>Y�$SYS0��4�g�-�I�E�EVx�#q'�PXWO��z �: $SK7!tf2%�Td�TRL��7; �'AC�`��nĠIND9DJ.D��_��f1��f���kPL�A�RWAj�D��SD�A��!+r||��UMMY9d҆F�10d�&���J�<��}1PR� 
�3�POS��J�= ��$V$^�q �L~�>��H��ܠK�?����CJ��@����ENE�@TƷ�A���_�RE�COR��BH �5 O�@=$LA�>$~�r2�R��`��q�b`�_Du��0R	O�@�aT[�Q��b�������! }У�PA�US���dETURYN��MRU� v CRp�EWM�b��AGNAL:s2$�LA�!?$=PX�@$P�y #A �Ax�C0 #ܠDO�`X�k�W�v��q�GO_AWAYF��MO�ae���]��CSS_CCSCB C �'N��CERI��гJ`u�QA0�}��@�GAG� R�0�`�`�{`��{`OF�q`�5��#MA��eX��A��LL�?D� �$���s�U�D)E%!`���O�VR10W�,�OR�|�'�$ESC_|$`�eDSBIOQ���l ��B�VIB&� �c,�����f�=pSSW���f!�VL��PL���AORMLO
��`�����d7%SC �bA1LspH�MPCh @�Ch �#h �#h 5�UU���C�'�C�'�#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$4�C��P3Wұ46$V7OLT37$$`�*�^1��$`O1*��$o��0RQY���2b4�0DH_TH�E����0SЯ4�7ALPH�4�`���7�@Q �0�qb7�rR�5�88� ×���"(��Fn�MӁ!VHBPFUAFLQ"Dt�s�`�THR��@i2dB�����G(��P�VP�����������1��J2�B�E�C�E�CPSu�Y@��Fb3��� H�(V�H:U�G�
X0��FkQw�[�Na�'B���C INHBcFILT���$��W �2�T1�[ ��$h���H YАAF�sDO��Y�Rp� fg �Q�+�c5h�Q�iSh�QPL���Wqi�QTMOU�#c�i�Q \��X�gmb��vi�h�biAi�fI�aHIG��ca	xO��ܰ��W�"vAN-u!��	#�AV�H!Pa8�$P�ד#p�R_:�A(�a��B�N0�X�MCN���f1[1�qVE�p��Z2;&f��I�QO�u�rx�wGldDN{G|d��a!F>!�9��aM:�U�'FWA�:�Ml��� X�Lu��$!����!l��ZO����0%O�lF��s�13�DI�W� @��Q���_��!�CURVA԰0rC	R41ͰZ�C<�r�H� v���<�`��<�(�f�CH�QR3�S���t0���Xp�VS_�`�$ד�F��ژ����-?NSTCY?_ E L����A1�t�1��U��24�2B�NI O7�����އDEVI|� �F��$5�RBT.xSPIB�P���#BYX����T���HNDG��G HC tn���L�@�Q�C���5��Lo0� H��閻�FBP�{tFE{�5�t�h�T��I�DO���uPMCS�v>�f�>�t�"HOTSWt�`s�?ELE��J T���e�2��2d5�� O� ��HA7��E��344�0>��A�K� �� MDL� 2J~PE��	A��@s��tːÈ�s�JÆ G!��rD"�ó�����&\�TO��W�	��/�ޅSLAV�L;  \0INPڐ����`%ن_CFd��M� $��ENU��OG��b�ϑ]Ռ�P�0`ҕ�]�I�DMA�Sa��\�WaR�#��"]�VE�$.a�SKI�STs��s$k$��2u���J��������	��Q���_S}Vh�EXCLUMq�J2M!ONL��D�YȔ�|�PE ղI_}V�APPLYZP���HID-@Y�r�_�M�2��VRFY��0��r�1�cIOC_f�� 1�����әO��u�LS���R$DUMMY3�!����S� L_TP/Bv�"���AӞ�ّ� N ���R�T_u�� �r�G&r[�O D���P_BA�`L�3x�!F ��_5�
��H������ ��� P $4 KwA�RGI��� q�2�O ��SGN�Z�Q �~P/�/PICGNs�l�$�^ �sQANNUN�@�T<�U/�ߴ�LAzp]	Z�d~�>EFwPI�@ �R @�F?IT~�	$TOTA%Š�d���!�M6�NIY�S+����E�A[�
DAYS\�ADx�@���	� �EFF_A�XI?�TI��0zC�OJA �ADJ__RTRQ��Up�!�<P�1D �r5̀Ll�T�p? ]P��"p��mtpd��V 0w�G������-��SK�SU� ���CTRL_CA��� W�TRA�NS�6PIDLE_PW���!��A��V��V_�l�V ?�DIAGS���X� /$2�_;SE�#TAC����t!�!0z*@��RRD��vPA���p ; SW�!�!�  ��o2l�U��oOH��3PP� ��IR�r���BRK'#��"A_A k���x 2x�9ϐZs2��%l�W�pt*��x%RQDW�%MS�x�t5AX�'�"��L?IFECAL���10��N�1{"�5Z��3{"dp5�ZU`}�M�OTN°Y$@FsLA�cZOVC@p��5HE	��SUPCPOQ�ݑAq� Lj �(C�1_X6�IEY
RJZRJWRJ�0TH�!�UC��6�XZ_ARl�p��Y2�HCOQ���Sf6AN��w$��ICTE�Y }`��CACHE��C9�M�PLAN���UFFIQ@@�Ф0<�1	��6
���MSW�EZ 8>w KEYIM�p��TM~�SwQq�wQ�#�����OCVIEܻ �[ A�BG�L��/�}�?� 	��?��D\p�ذST��!�R� �T� ��T� �T	��PEMA�If�ҁ��_F�AUL�]�RцĆ1�U�� �TR�E�^< �$Rc�uS�% IT��BUFW}�W��9N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTT(����sP��M��Ot�T�LwAX � ��XX~`9#�c_G�3
ЧYN_1�_�D���1 �2M�*��T�F��H@ ~g�`� 0p���Gb-sC_R�AIAK���r�t�RoQ8�u7h�qDSPq��rP��A�IM�c6�\����s2�U�@�A�s�M*`IP���s�!D��6�TH�@n�)�OyT�!6�HSDI3��ABSC���@ V`y��� �_D�/CONVI�G��H�@3�~`F�!�pd��psqSCZ"���sgMERk��qFB��Lk��pET���aeR�FU:@DUr`����x�CD,���@p;cJHR�A!��bp�ՔՔ+PSԕCJ���C��p���єSp�cH *�LX�:cd�Rqa�|  ����W��U��U���U�	�U�OQU�7R�8BR�9R��0T�^�1k�U1x�1��1��1��U1��1��1ƪ2Ԫ�2^�k�2x�2��2���2��2��2��2*ƪ3Ԫ3^�3k�x��3���o���3��3j��3ƪ4Ԣ�HsXTk!0�d <�  7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr�����.�2REM� Fj��B�OVM��A�T7ROV�DT�`-�MX<�IN��0,�NW!INDKЗ
w�<׀�p$DG~q3�6��P�5�!D�6�R�IV���2�BGEA-R�IO�%K�¾DN�p��J�82�PB@>�CZ_MCM�@�1���@U��1�f ,<②a? ���P�I�!?I�E���Q�4���`m���g�� _0Pfqg RI�9ej�k!UP2_ khh��cTD�p@���! a���-��wBAC�ri T�Ph�b�`�) OG���%���p��IFI��!�pm�>��	�PT��"��MR2��j ��Ɛ+"�� ��\��������$�B`�x%��_ԡ�ޭ_����� M������D�GCLF�%DGDMY%LDa��5�6P�ߺ4@��Uk���? T�FS#p�Tl P���e�qP�p$EX_����1M2��2� 3�5���G ���m ���Ѝ�SW�eOe6D�EBUG���%G�R���pU�#BKUv_�O1'� �@PO�I5�5�MS��OOfswS�M��E�b�Q�0�0_?E n �p� �TERM�yo�Q��ORI+��p��P�SM_����b�q��@TAr�r�C��UP�R�s� -�1�2�n$�' o$SEyG,*> ELTO���$USE�pNFIAU"4�e1���>#$p$UFR���0`ؐO!�0����OT�'��TAƀU�#NST�PAT��P�"OPTHJ����E�P8 rF�V"ART�``%pB`�abU!REL:�aSHFT��V!�!.�(_SH+@M$���"� ��@N8r�����OVRq��rSHI�%0��UN� �aAY#LO����qIl���p�!�@��@ERV]� �1�?:�¦'�2��0%��5�%�RCq��E�ASYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba���
5Po��0�p6OeR�MY� `GR��t2b5n� � ��8UPa�Uu Ԭ")�]��TOCO!S�1POP ��`�pC��������Oѥ`R%EPR3��aO�P�b�"ePR�%WU.X|1��e$PWR��3IMIU�2R_	S�$�VIS��#(AUDp��~�av" vh��$H���P_AD+DR��H�G�"�Q��Q�QБR~pDp1�w H� SZ�a��e`�ex�e��SE�l�r��HS��MNv?x ���%Ŕ��OL���p<Px��-��ACROlP<_!QND_C��גx�1�T �ROUPT���B_�VpQ�A1 Q�v��c_��i���iр�hx��i���i��v�AMCk�IOU��D�g�fsu^d�y $|�P_D��VB`b�PRM_�bi�H�TTP_אHaz{ (��OBJEr�l�P��$��LE�#��s`{ � \��u�AB_x�T~��S�@�DBGL�V��KRL�YHIoTCOU�BGY �LO a�TEM���e�>�+P'�,PSS�|�P�JQUERY�_FLA�b�HW(��\!a|`u@�3PU�b�PIO��"��]�ӂ/dԁ=dԁ�� _�IOLN��}�����CXa$SL�Z�$INPUTM_g�$IP#�P��L'���SLvpa~���!�\�W�C-�BMyF���pF_ASv��$L ��w �DF1G�U�B0m!���0HY��ڑ��ܓ��UOPs� `������[�ʔ[�і"�[PP�SIP�<�і�I�2��IP_MEsMB��i`� X��cIP�P�b{�_N�`����R�����bSP��p$FO�CUSBG�a��U=J�Ƃ �  � �o7JOG�'�DI�S[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A���APHIb�Qt�]�D� J7J\����� _KEYt�� �KՀLMO�Na���$XR���ɀ��WATCHa_��3���EL��b}Sy����s� ���!V�g� �CTR�3򲓥��LG�D�� �R��I�
LG_SIZ���J�q XIƖ�I�FDT�IH� _�jV�GȴI�F�%S O���q �Ɩ���v������K�S����w�kR�N����E�@�\���'�*�U�s�5��@L>�4�DAUZ�EA�pՀ�Dp�f��GH�B���BOO>��� C���P�IT���� ��RE=C��SCRN�����D_p�aMARG f�`��:���T�L���S�s��W�Ԣ�I�JGMO�MNC�H�c��FN��R�Knx�PRGv�UF���p0��FWD��HL.��STP��V��+�X��Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28�����Gh�0PO��������M8�Ģ��EX��TUIv�I��(�4�@� t�x�J0J�~�P��J0r��N�a�#ANA���O"�0VAIA��dC�LEAR�6DCS�_HI"�/c�O��O�SI��S��IGN_�vpq��uᛀT�d� DEV�-�LLA �°BUTW`��x0T<$U�EM��Ł��T��0�A�R��x0p�σ�a�@OS1��2�3�`�`� �ࠜh�AN%-���.-�IDX�DP�2MRaO��Գ!�ST���Rq�Y{b! �$E&C+��p�.&A&���`� L ��ȟ%Pݘ��T\Q�U�E�`�Ua��_ � �@(��`������# �MB_PN�@ R`r��R�w�TR�IN��P��BAS�S�a	6IRQ6�aMC(�� ���CLDP�� ETRQLI��!D�O9=4FLʡh2�Aq3z1D�q7��LDq5[4q5ORG�)�2� 8P�R��4/c�4=b-4�t� �rp[4*�L4
q5S�@TO0Qt�0*D}2FRCLMC@D �?�?RIAt,1ID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCESJ?R�EMhPa�͠��BD4�E�q`�`�F_A�J�C[��O�H� K��� \ȶ��bTf$� ��LI��q�SREQUIR�E�#MO�\�a�XD�EBU��,1L� M䵔 �p���P�c�AA,1N��
Q�qa�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N�a�NdPST9� w� 4��LOC��RI���EX�fA�NG��A,1ODA5Q䵗�@$��9�ZMF�����f��"���%u#ЖVSUPܡ%���FX�@IG=Go�� �rq�"���1��#B��$���p% #by��rx���vbPODATAK�pE;�ȥ��R��M��*� �t�`MD�qI��) �v� �t�A�wH�`���tDIAE��sAN�SW��th���uD���)��aԣ(@$`�[ PCU_�V6��ʠ�d�PLOr�$`�HR���B���B�p�t����,1RR2�E��  ��V�A�/A d$CALII�@��G~�2���!V��<$R�S�W0^D"��ABC~�hD_J2SE�Q\�@�q_J3M�
G�G1SP�,��@PG�Bn�3m�u�3p�@���JkC���2'AO)IyMk@{BCSKP^:�ܔ9�wܔJy�{BQ�ܜ�����`_A1Z.B��?�EL��YAOCMP�c|A)���RT�j���1�ﰈ��@1�������Z��SMG��pԕf� ER!��2a[INҠACk�p�����b�n _���@����D�/R��3DIU��CDH�@
�:#a�q$V�Fc6�$x�$���`0@���b��Á�E��H �$BE�LP����!ACCE�L���kA°IR�C_R�pG0�T<!�$PS�@B2L`���W3�طx9� ٶPATH���.�γ.�3���p�A_@��_�e�-B�`C�_MG�$D�D��ٰ��$FW��@�p����γ����D}E��PPABN�ROTSPEEu�����O0��DEF�>Q��`$USE)_��JPQPC��J�Y����-A 6qYN��@A�L�̐�L�M�OU�NG��|�O9L�y�INCU��a��¢ĻB��ӑ�AENCS���q�B�����D�IN�IY����p�zC�VE�����2�3_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��rPRC����MOS� �gTMOpp�@-GPE�RCH  M�OVӤ �����!3�yD�!e�]�6�<�� ʓAY���LIʓdWɗ��p:p3�.�I�TRKӥ�AY����?Q^�Ym�b��`p�CQ�� MOM�B?R�0u��D����y�0Â��D�UҐZ�S_BCKLSH_CY���o� n��TӀ���
c��CLALJ��A8��/PKCHKO0��Su�RTY� �q���M�1�q_
#c�_�UMCP�	C���SsCL���LMTj��_L�0X����E �� �� ���m�`h���6��PC��B��H� �P�ŞCN@�"XT����CN_b��N^C�kCSF����V6����ϡjY���nCAT�SH s�����ָ1���֙�0��������PA���_P���_P0� e�`��O1u�$xJG� �P{#�OG���TORQU(�p�a�~�����Ry������"_W ��^�����4t�
5z��
5I;I ;Iz�F��`�!��_8�1��VC"��0�D�B�21�>	P8�?�B�5JRK�<�2��6i�DBL_SMt�Q&BMD`_DLt�&BGRV4
Dt�
Dz��1H_���31�8J�COSEKr�EHLN �0hK�5oDt�jI��jI <1�J�LZ1�5Zc@y���1MYqA�HQBTH|WMYTHET09�NK23z�/Rn�r@[CB4VCBn�CqPASfaYR<4gQt�gQ�4VSBt��R?UGT	S���Cq��a��P#x���Z�C$DUu  ��R䂥э2�Vӑ��9Q�r�f$NE�+p!Is@�|� �$R�#Q�A'UPeYg7EBHBALCPHEE.b�.bS�E �c�E�c�E.b�F�c�j�FR�VrhVghd��lUV�jV�kV�kV�kUV�kV�kV�iHrh@�f�r�m!�x�kH�kUH�kH�kH�kH�i�OclOrhO��nO��jO�kO�kO�kO*�kO�kO�FF.bTQ𰉔E��egSPBA�LANCE��RLmE�PH_'USP���F��F��FPFULC�3��3��E��{1�l�UTO_p ��%T1T2t���2NW�����ǡ��5�P`�擳�T�OU�|��� INSEG���R�REV��R���D3IFH��1���F�1�;�OB��;C���2� �b�4LC�HWAR��;�AB�W!��$MECH`]Q�@k�q��AXk��P��IgU�i�� �
���!����ROBF��CR��ͥ*��C��_s"T �� x $WEI3GHh�9�$cc�2� Ih�.�IF ќ�'LAGK�8SK��nK�BIL?�OD��LU��STŰ�P䑄; � ����������
�Ы�L��  �2�`�"�DEBU�.�L&�n��PMMY9��NA#δ9�g$D&���$��܅ Q �DOu_�A��� <	� ��~��L�BX�P��N��+�_7�L�t�O�H  �� %"��T���ѼT������TICK/�C�TE1��%������N��c�Ã�R L�S����S�����PROMP�h�E� $I�R� X�~ ���!�MCAI�0��j���_9�C���t�l�R�07COD��FU`�+�ID_" =����耿G_SUFF<0 �3�O����DO��ِ��R��Ǔن�@S����!{������	��H)�_FI��9n��ORDX� �����36��X���Ɩ�GR9�S��ZD�TD��t�ŧ�4 *�L_NA�4���K��DEF_I[�K���g��_����i��Ɠ�š���IS�`i �萚�����e����4�0i�DPg����D� O�>�LOCKEA!u���ϭϿ���{�u�UM z�K�{ԓ�{ԡ�{��� ��}��v�Ա��g� �����^���K��@�����!w�N�P'� ��^���,`�W\�[6R�
��TEF��� �OULO�MB_u�0�V�ISPITY�A��!OY�A_FRId��(�SI���!R������3����W�W��0��0_,�EAS%��!��& "���4p�G�;� h ��7�ƵCOEFF_O m���m�/�G!%�S.�߲CA5�����u�GR` � �� $R� �X]�TME�$R�s�Z�,/,)�ER�T;�:�n���  ]�LL�:�S�_SV�($~����@����� "SETU��MEA��Z�x0��u������ � l� �� ȰID�" ���!*��&P���*�F�'����)3��#���"�5;`*���REC���!���MSK_���� P	�1_USER��,��4���D�0��VEL,2�0���2�5S�I��0�MT�N�CFG}1� � ���Oy�NO�RE��3��2�0SI����� ��\�UX�-�ܑPDE�A $KEY_��}��$JOG<EנSVIA�WC�� 1�DSWy���
��CM7ULT�GI�@@�C��2� 4 p�#t�+�z�XYZ���쑡���z� �@_ERR��� ��S L��-���@��s0BB/$BUF-@X1��MOR�� H	�CU�A3�z�1Q��
��3���$���FV��2TbG��� � $S1I�@ G�0VO B`�נOBJE&�!FA�DJU�#EELA�Y' ���SD�WOU��мE1PY���=�0QT i�0�W�DIR$ba�pےʠGDYNբHeT�@¥�R�^�X����O�PWORK}1�},�SYSBU@p 1SOP�aR�!�j�U�k�PR��2�eP�A�0�!�cu� 1OP���UJ��a'�D^�QIMAG�A	���`i�IMACrIN�,�bsRGOVR!D=a�b�0�aP�`s@ʠ� �^uz�LP��B�@��!PMC_QE,�Q��N@�M�r�Ǳ��1Ų��=qSL�&�~0���$OV�SL\G*E��*E2y�Ȑ�_=p�w��>p �s���s	�����=q�#}1� @�@;���MOE�RI#A��
N� �X�s�f�ՠ���P�L}1�,RTv�m�A�TUSRBTRC_T(qR��B ������$ �Ʊ��,�~0� !D��`-CSALl`�`SA���]1gqXE�� �%���C��J�
�Ʊ�UP(4����PX���؆�q��3�w� ��PG�5� $SUB���������t�JMPWAI�TO��s��LOyCF8t�!D=�CVF	ь��y���R`�0��CC�_CTR�Q�	�I�GNR_PLt�D�BTBm�P��z�B�W)����0U@���I�G�a��Iy�TNL�N��Z�R]aK� N��B�0�PE�s���r܊�f�SPD}1� L	�A�`gఠ�S��CUN�{���]�R!�BDLY�2���tP^��H_PK�E��2?RETRIEt��2f�b)���FI�BǼ ����8� �2��0DBGLV~�LOGSIZ$C��KTؑUy#u�D�7�_�_T1@�EMB�@C\1A����R��|D�FCHECKK��R�P�0����@�&�(bLEc�" PA�9�T���P�C߰P4N�����ARh�0Ґ��Ӯ�PO�BORMATTnaF�f1�h���2�S��UX�y`	��LB��4� � rEITCH����p19PL)�AL_ � $���XPB�q� C,2Dx�!��+2�J3D���� T�pPDCK�yp��oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYL�OA��m�_1t�2<t���J3AR�����դ֏�laTIA4��5��6,2MOM�CP�����������0BϐAD��������PUBk`R��;����;���.��z4�` I$PI\Ds�o�@�1yՕ�w�2�w�Z��I��I��I���p� ���n���y�e`��9S)bT�SPEED� G��(�Е��/��� Е�`/�e�>��M�<�ЕSAMP�6V0��/���ЕMO�@ 2@�A��QP���C�� n�����������LRf`�kb�ІE9h�EIN 09��7S.В9
�yPy�GAMM�%S���D$GE�T)bP�cD]��2
��IB�q�I�G$HI(0;A��LR�EXPA8)LWVM8z)���g���C5�CHKhKp]�0�I_�� h`eT��n�q���eT,���� ��$�� 1�iPI>� RCH_D�313\��30LE�1�1\��o(Y�7 �t�MSW�FL �M��SCRc�7�@�&��%n�f�;SV���PB``�'�!�B�sS_SAaV&0ct5B3NO]�C\�C2^�0�mߗ� uٍa��u���u:e;��1���8��D�P��� ������)��b9� �e�GE�3��V������Ml�� � F�YL��QNQSRlbfqXG�P�RR�#dCQp� �S:AW70�B�B[�CgR:AMxP�KCL�H���W$�r�(1n�g�M�!o��� �F�P@}t$WP�u�P r��P5� R<�RC�R��%�6@�`��� ��qsr X��	OD�qZ�Ug�ڐ>D�� ��OM# w�J?\?n?�?�?��9��b"�d�]�_��� |��X0��bf��qf@��q`�ڏgzf��EڐN� Ag�"�ܰ���FdPB��PM��QU�� � =8L�QCOU!5�7QTHI�HOQBp7HYSY�ES��q�UE�`�"�O��ˋ  �P�@\�U)N���Cf�O�� P��Vu��!�����OGRAƁcB22�O�tVuITe �q^:pINFO����h�{�qcB�e�OI�r�� (�@SLEQ@S��q��p�vgqS�ލ�� 4L�EN�ABDRZ�PTIO�Nt�����Q���)�G�CF��G�$JX�q^r�� R����U�g�5BOS_E9D����� �F��P�K��E'N9U߇وAUT$1܅COPY�����n��00MN���PWRUT8R �Nx�;OU��$G[rf�}
e�RGADJ����*�X_:@բ$P�����P��W��P��`} ��)�}�EX�kYCDR|�NS.�9�F@r�LGO�#��NYQ_FREQ�R�W� �#�h�TsL�Ae#����ӄ �CcRE� s�IF�ᶕsNA��%a�_}Ge#STATUI`<e#MAIL������q t�������EwLEM�� �/0><�FEASI?�B ��n�ڢ�1�]� � I�p��Y!q]�Lt#A�ABM���E�pr<�VΡY�BASR҈Z��S�UZ��0�$q���RMS_TR;�qb ���SY��	�ǡ��$���>C��Q`	� 2� _�TM������̲��@ �A��)ǅ�i$D�OU�s]$Nj���P�R+@3���rGRIyD�qM�BARS �sTY@��OTO�Rp��� Hp_}�!����d�O�P/�� �s �p�`POR�s���}���SRV��),����DI&0T��Ѡ�� #�	�#�4!�5*!�6!�7!�8�e��F�2��Ep$VALUt��%��ֱ��>/��� ;�1ėq�����(_�AN��#�ғ�Rɀ(���T�OTAL��S��P�W�Il��REG#EN�1�cX��ks0(��a���`TR��R��_S� ��1ଃV �����⹂Z�E��p��q��Vr���V_Hƍ�DA�S����S_�Y,1�R4�S� AR��P2� ^�IG�_SE	s����å_�Zp��C_�Ƃ�EN�HANC�a� T ;�������GINT�.��@FPs^İ_OVRsP�`@p�`��Lv��o��7�p}��Z�@�SLG�
AA�~�25�	��Dd��S�BĤDE�1U�����TE�P���� !Y��
��J��$2�IL_M`C�x r#_��`TQ�`���q���'�BV�CF�P_� 0�M�	[V1�
V1�2�U2�3�3�4�4�
�!���� � m�A�2IN~VIB�P���1�2�2��3�3�4�4��A@-�C2���=p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KEEP_HNADD!�!`$^�j)C�Q�� �$��"	��#O�a_$�A�!�0�#i��#REM�"�$��½%�!��(U}�e�$HPW�D  `#SBWMSK|)G�qU�2:�P	�COLLAB� �!K5�B�� 4��g��pITI1{�9p#>D� ,�@F�LAP��$SYNT �<M�`C6���UP_DLYAA�ErDELA�0ᐢ�Y�`AD�Q� ��QSKIP=E� i���XpOfPNTv�A�0P_Xp�rG�p �RU@,G��:I+�:IB1 :IG�9JT�9Ja�9Jn��9J{�9J9<��RA=s� X���4��%1�QB� NFLIC�s�@J�U�H�LwNO_H�0�"?��R�ITg��@_PAz�pG�Q� ��
^�U��W��LV�d�NGRLT�0_q���O�  " ��OS��T_�JvA V	�APPR�_WEIGH�sJg4CH?pvTOR��vT��LOO��]�+�"tVJ�е�ғA�Q�U��S�XOB'�'�{�J�2P���7�X�T �<a43DP=`Ԡ\"<a8�q\!��RDC��LW� �рR��R�`� �RV��jr�b��RGE��*��cN�F�LG�a�Z���SP9C�s�UM_<`^2TH2NH��P.a� 1� m`E�F11��� l�Q �!#� <�p3AT � g�S�&�Vr�p�tMq��Lr���HOMQEwr�t2'r�-@?Qcu��w3'r�������w4'r�'�9�K�]�o����w5'r뤏��ȏPڏ����6'r�!�@3�E�W�i�{��7'r힟��ԟ����8'r��-�?�Q�c��u��S$0�q�p �� sF��`)a�"`P�����`/���-��IO[M�I֠���*�POWE�� ��0Za�0p��� �5��$DS=B GNAL���0�Cp��*laS23�23�� �~`���� / ICEQP��P1Ep��5PIT�����OPBx0��FLOW�@TRvP��!U�֤�CU�M��UX�T�A��w�ERFA�C�� U��vɲCH��� tQ b _��>�Q$����OM��A�`T\�P#UPD7 A�c2t�T��UEX@����U EFA: X"�1�RSPT�����T ��PPA�0o�6�`EXP�IOS���)ԭ�_���%��FC�WR�A��ѩD�a�g֕`ԦFRIENDsaC2UF7P�����TOOL��MYH� C2LENGTH/_VTE��I��Ӟ�$SE����U�FINV_����RGI�{QIT�I5B��Xv��-�G2-�G17�w�SG�DX��_��UQQD=#@���AS��d~C�`���q�� �$$Cz/�S�`������S0f�����VERS�I� ��f��5��I���������AAVM_Y�2 �� 0  �5���C�O�@�r� �r�	 ����S0�����������������
?QY�BS����1��� <-��� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O�iCC�@XLMT���C�  ���DIN�O�A�Dq�EKXE�HPV_���ATQz
��LA�RMRECOV ��RgLMD/G *�5�O�LM_IF *��`d�O�_�_�_�_�j�_'o9oKo]onm, 
��odb��o��o�o�o^��$� <z, A   2D{��PPINFO u[ �Vw��������`�� �����*��&�`�@J���n�����DQ� ���
��.�@�R�d��v���������a
PP�LICAT��?��P��`�Handling�Tool 
� �
V8.30P/�40Cpɔ_LI�
883��ɕ$?ME
F0G�4��-
398��ɘ�%�z�
7DC3�ɜ
��NoneɘVr�|��ɞ@6d�� Vq_ACTI�VU��C죴�M�ODP���C�I��HGAPON���n��OUP�1*�� i�m����Қ�_����1*�  �@�������� Q���Կ�@�
������ ����5�Hʵl�K�?HTTHKY_�� /�M�SϹ�������� �%�7ߑ�[�m�ߝ� �ߵ����������!� 3��W�i�{���� ����������/��� S�e�w����������� ����+�Oa s������� '�K]o� �������/ #/}/G/Y/k/�/�/�/ �/�/�/�/�/??y? C?U?g?�?�?�?�?�? �?�?�?	OOuO?OQO cO�O�O�O�O�O�O�O �O__q_;_M___}_ �_�_�_�_�_�_kŭ��TOp��
�DO_CLEAN9��pc_NM  !{血�o�o�o�o�o��D?SPDRYRwo��HI��m@�or� ��������p&�8�J���MAXݐ Wdak�H�h�XWd��d���PLUGGpW�Xgd��PRC)pB�`�kaS��Oǂ2DtSEGF0�K� �+��o�or�����������%�LAPOb�x�� �2�D� V�h�z�������¯ԯ|�+�TOTAL��|��+�USENUO��\� e�A�k­�R�GDISPMMC�.���C6�z�@@$Dr\�OMpo�:�X��_STRING �1	(�
��M!�S�
��_�ITEM1Ƕ  n������+�=� O�a�sυϗϩϻ����������'�9��I/O SIGN�AL��Try�out Mode�ȵInpy�Simulateḏ�Out��O�VERRLp = �100˲In �cycl�̱P�rog Abor���̱u�Stat�usʳ	Hear�tbeatƷM?H Faul	��Aler�L�:�L� ^�p��������� ScûSaտ�� -�?�Q�c�u������� ��������);pM_q��WOR.� û������ +=Oas�� �����//'.PO����M �6/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~?��?�?�?�?H"DEV P.�0d/�?O*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_PALT	��Q� o_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o��o�o�o�_GRI m�û9q�_as� �������� '�9�K�]�o�������'�R	�݁Q��� �)�;�M�_�q����� ����˟ݟ���%�x7�I�ˏPREG�^ ����[�����ͯ߯� ��'�9�K�]�o����������ɿۿ�O���$ARG_� D �?	���0���  w	$O�	[D��]D��O�e�#�SB�N_CONFIG� 
0˃����}�CII_SAV/E  O������#�TCELLSE�TUP 0�%�  OME_IO�O�O�%MOV_qH������REP���J��UTOBAC�K�����FRA:\o� �Q�o���'`��|o��� � �� f�o������*�!�3�`�Ԉ�� f����������o� {��&�8�J�\�n��� ���������������� "4FXj|�������끁�  ��_i�_\A�TBCKCTL.�TMP 6.VD� GIF PHD�_q��N�t�#��f�INI�P�o���c�MESSAG�����8��ODE_D����z���O�0�c�PAU�SM!!�0� (�73�U/g+(Od/�/x/�/�/�/�/ �/�/???P?>?t?�1�0$: TSK  �@-��T�f�UPD�T��d�0
&XWZD_ENB����6STA�0��5�"�XIS��UNT� 20Ž� �� 	 ��z���en�g�-뷛��S�o�U@��H����xH�Oo�}CUw�g�^����.�O�O�O�O/_2F�MET߀2CMP�TAA��@��$A-�@����@���@����]5��5��(d5��P5��r�5F*5��338]SCRDC�FG 1�6K�Ь�Ź�_ �_oo(o:oLo��o�Q���_�o�o�o�o�o �o]o�o>Pbt����o9�i�GR`<@M/�s/NA��/�	i��v_E�D�1�Y� 
� �%-5ED�T-�'�GET�DATAU�o�9��u?�j�H�o�f��\��A��  ���2�&�ȏE�D����~�ŏ׏m����3 ��&��J�\�ߟJ�����9�ǟ�4���ϯ �\����]�o�����5N������\�w�@�)�;�ѿ_��6� ��gϮ�\�CϮ������+��7��V�3�z� \��z�����i����A8�ߜ���]����F�ߟ�5����9~������]����`Y�k�����CR� !ߖ���W�q���#�5����Y��p$�NO_D�EL��rGE_U�NUSE��tIG�ALLOW 1���(*S�YSTEM*S�	$SERV_G�R�V� : REGƟ$�\� NU�M�
��PMU|B ULAYNP�\PMPA�L�CYC10�#6 $\UL�SU�8:!��Lr�BOXOR=I�CUR_���PMCNV��10L�T4�DLI�0��	�� ��BN/`/r/�/�/�/�/�/���pLAL_?OUT �;����qWD_ABOR�=f�q;0ITR_�RTN�7�o	;0NgONS�0�6 
H�CCFS_UTI�L #<�5CC�_@6A 2#; h ?�?�?O#O6]�CE_OPTIO�c8qF@RI'A_Ic f5Y@�25�0F�Q�=2qz&}�A_LIM��2.� ��P��]B��KX�P
��P�2O�Q��B�r�qF�PQ5T1�)TR�H�_:JF_�PARAMGP 1�<g^&S�_��_�_�_�VC�  +C�d�`�o!o�`�`�`�`�Cd��Tii:a:e>e�Ba�GgC�`� D_� D	�`�w�?��2HE ON�FI� E?�aG_Pv�1#; � ��o1CUg|y�aKPAUS�s1�yC ,�� �������	� C�-�g�Q�w�������Ы�я���rO�A��O�H�LLECT�_�B�IPV6�ENp. QF�3�NDE>�� �G�71�234567890��sB�TR����%'
 H�/%)�� �����W���0�B��� f�x���㯮���ү+� ����s�>�P�b��� �������ο��Kπ�(�:ϓ�^�|��B!�F� �I|�IOG #��<U%e6`�'�9�K���TR�P2$��(9X�t�Yކ�`%�̓ڥH��_�MOR�3&�=�>�@XB��a� �A�$��H�6�l�~���~S��'�=�r_A? �a�a`��@K��RʭdP��)F�haÃ-�_�'�9�%
@�k��G� ��%Z�^%��`�@c.��PDB��+���cpmidbg��	�`:��@�eTR���p��N  �f�,	���]ܭ@s<�^���sg�$��fl�q��ud1:��:J��?DEF *ۈ���)�c�buf.txt�����_L64FIX ,������l/[Y/ �/}/�/�/�/�/
?�/ .?@??d?v?U?�?�?��?�?�?�?,/>#_E -���<2ODO`VOhOzO�O6&IM���.o�YU>����d�
�IMC��2/�����dU�C��20��M�QT:Uw�Cz � B�i�A����A���Au�g�B3�*CG��B<�=w�i�B.���B���B���5B�$�D��%B���ezVC��q�C�v�D����D-lE?\D�n�j����29"��22o��D|����� �𺪢�C�C���e�
�xObi�D4cdv`D��`/�`v`s]�E�D D�` �E4�F*� ?Ec��FC��u[�F���E��f�E��fFކ3�FY�F�P3��Z��@�33 ;?��>L���Aw��n,a@��@e�5!Y���a���`A��w�=�`<#���
��?��ozJRSMOFST (�,bI+T1��D @3��
�c�����a��;��b�w?���<��M�NTESTR�1O�CR@�4�4�>VC5`A�w�Ia�+a�aORI`CTPBՖU�C� @4����r��:d����qIj?�5��qT_�?PROG ��
��%$/ˏ�t��NUS/ER  �U�������KEY_TBL'  ����#a��	
��� !"�#$%&'()*�+,-./��:;�<=>?@ABC��GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?�����������LCK�
����S�TAT/��s_AU�TO_DO ��	�c�INDT_ENBP���Rpqn�`�sT2����STOr`쓯�XC�� 26����8
SONY XC-56��"b����@��F(� А�H�R50w���>�P�7<b�t�Aff����ֿ� Ŀ����C� U�0�yϋ�fϯ��Ϝ���������-ߜ�TR�L��LETEͦ ���T_SCRE�EN ���kcs���U�MMENU 17�� <ܹ���w� ��������K�"� 4��X�j������ ������5���k�B� T�z������������� ��.g>P� t������ Q(:�^p� ���/��;// $/J/�/Z/l/�/�/�/ �/�/�/�/7?? ?m? D?V?�?z?�?�?�?�? �?!O�?
OWO.O@OfO��OvO�O�O(y��RE�G 8�y�����`�M�ߎ�_MAN�UAL�k�DBC�O��RIGY�9�DBG_ERRL��9�ۉq��_�_��_ ^QNUML�I�pϡ�pd
�
�^QPXWORK 1:���_5oGoYo�ko}oӍDBTB_NN� ;������ADB_A�WAYfS�qGC�P 
�=�p�f_A!L�pR��bbRY�[�t
�WX_�P 1<{y�n�,�%oc�Pl��h_M��ISO���k@L��sONTImMX��
���v�y
��2sMOTN�END�1tREC�ORD 1B��� ���sG�O� ]�K��{�b�������� V�Ǐ�]����6�H� Z���������#�؟ ������2���V�ş z��������ԯC��� g��.�@�R���v�� ��	���п���c�� ��#ϫ�`�rτϖ�� ��)ϳ�M���&�8����\�G�Uߒ��8�������K� �����6��%RC7�n����ߤ������A�4���$���H�3�A�~��;��������9���]������|��B#Zl���zTO�LEREN\�rB��'r�`L��^PC�SS_CCSCB' 3C>y�`IP�� }�~�<�_` r�K�����/�{��5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O��O�O�O�O_�~�L5L� D��&qET|�c�a C[�C��PZP^r_ A�� p� �sp�x�QGPt[	 A�p�Q�_�[? �_�[oU�p�P�pSB�V�c�(a�PWoPio{h+�o�X�o�oY��[	r�h�LW��N:p����}�6ګ�c��aD@VB���|�G���+��K� �otGhXGr�So�����eB   =���Ͷa>�tYB��� �pC�p�q�aA"�H�S�Q-��q����ud�v�����AfP w` 0���D^P���p@�a
�QAXTHQ����a a"W>� �a9P��b�e :�L�^�h�Hc�́PQ�RFQ�PU�z�֟ �o\^��-�?��c��u����zCz��ů�b2�Щ�RD�;����l)*��� �S̡0��]�0�.��@���EQ�p��F�X� ѿUҁп�VSȺ�NSTCY 1E��]�ڿ��K� ]�oρϓϥϷ����� �����#�5�G�Y�k��}ߏߒ��DEVI�CE 1F5� MZ�۶a��	� ��?�6�c���	{䰟�����_HNDGD �G5�VP���R�LS 2H�ݠ��/��A�S�e�w����� ZPARAM I��FgHe�RBT [2K��8р<�߬WPpC�C��,`¢�P�Z�z��%
{�C��2�jMTLU0,`"nPB, s ��M� }�gT�g��F
B��!�bc y�[2Dchz� ���/��/gT�#I%D��C�`� b!�R��A���A,��Bd��kA�;���_C4kP��!2�C��$Ɓ�]��ffA�À��+B�� �| ���/�/�T (��54a5 �}%/7/d?/M?_? q?�?�?�?�?�?O�? OO%O7OIO�OmOO �O�O�O�O�O�O�OJ_ !_3_�_�_3�_�_�_ �_�_o�_(ooLo^o Ё=?k_IoS_�o�o�o �o�o�o�o#5 G�k}���� ���H��1�~�U� g�y�ƏAo�Տ��� 2�D�/�h�S���go�� ��ԟ����ϟ��� R�)�;���_�q����� �����ݯ�<��%� 7�I�[�m�������� �}�&��J�5�n�Y� �ϤϏ��ϣ�ѿ�� ����F��/�Aߎ�e� w��ߛ߭��������� B��+�x�O�a��� ���������,���%� b�M���q��������� ������L#5 �Yk}���  ��61CU g������� �	//h/���/w/�/ �/�/�/�/
?�/.?@? I/[/1/_?q?�?�? �?�?�?�?�?OO%O rOIO[O�OO�O�O�O �O�O&_�O_\_3_E_ W_�_?�_�_�_�_�_ "ooFo1ojoE?s_�_ �om_�o�o�o�o�o0 f=Oa�� �������� b�9�K���o���Ώ�� [o��(��L�7�I����m������$DC�SS_SLAVE L���ё���_4�D  љ��C�FG Mѕ��������F�RA:\ĐL-�%04d.CSV���  }�� ���A� i�CHq�z�������|�����  �����Ρޯ̩ˡҐ�-��*����_C�RC_OUT �N������_F�SI ?њ ����k�}��� ����ſ׿ ����� H�C�U�gϐϋϝϯ� �������� ��-�?� h�c�u߇߽߰߫��� ������@�;�M�_� ������������� ��%�7�`�[�m�� �������������� 83EW�{�� ����/ XSew���� ���/0/+/=/O/ x/s/�/�/�/�/�/�/ ???'?P?K?]?o? �?�?�?�?�?�?�?�? (O#O5OGOpOkO}O�O �O�O�O�O _�O__ H_C_U_g_�_�_�_�_ �_�_�_�_ oo-o?o hocouo�o�o�o�o�o �o�o@;M_ �������� ��%�7�`�[�m�� ������Ǐ������ 8�3�E�W���{����� ȟß՟����/� X�S�e�w��������� �����0�+�=�O� x�s���������Ϳ߿ ���'�P�K�]�o� �ϓϥϷ��������� (�#�5�G�p�k�}ߏ� �߳����� ����� H�C�U�g����� �������� ��-�?� h�c�u����������� ����@;M_ �������� %7`[m �������/ 8/3/E/W/�/{/�/�/ �/�/�/�/???/? X?S?e?w?�?�?�?�? �?�?�?O0O+O=OOO�xOsO�O�O�O�O�C��$DCS_C_F�SO ?�����A P �O�O_?_:_ L_^_�_�_�_�_�_�_ �_�_oo$o6o_oZo lo~o�o�o�o�o�o�o �o72DVz �������
� �.�W�R�d�v����� ��������/�*� <�N�w�r��������� ̟ޟ���&�O�J� \�n���������߯گ ���'�"�4�F�o�j� |�������Ŀֿ�������G�B�T��OC_RPI�N_jϳ� ���ς��O����1�Z�,U��NSL��@&�h� ����������"��/� A�j�e�w����� ��������B�=�O� a��������������� ��'9b]o �������� :5GY�}� �����/// 1/Z/U/g/y/�/�/�/ �/�/�/�/	?2?-??? Q?z?u?��ߤ߆?�? �?�?OO@O;OMO_O �O�O�O�O�O�O�O�O __%_7_`_[_m__ �_�_�_�_�_�_�_o 8o3oEoWo�o{o�o�o �o�o�o�o/ XSew���� ����0�+�=�O� x�s���������͏ߏ ���'�P�K�]�o������ �PRE_C�HK P۫�A� ��,8�2��� 	 8�9�K���+�q��� a�������ݯ�ͯ� %��I�[�9����o� ��ǿ��׿���)�3� E��i�{�YϟϱϏ� ����������-�S� 1�c߉�g�y߿��߯� ���!�+�=���a�s� Q���������� ����K�]�;����� q�������������# 5�Ak{� �����C U3y�i��� ���/-/G/c/ u/S/�/�/�/�/�/�/ ??�/;?M?+?q?�? a?�?�?�?�?�?�?�? %O?/Q/[OmOO�O�O �O�O�O�O�O_�O3_ E_#_U_{_Y_�_�_�_ �_�_�_�_o/ooSo eoGO�o�o=o�o�o�o �o�o=-s �c������ �'��K�]�woi��� 5���ɏ�������� 5�G�%�k�}�[����� ��ן�ǟ����C� U�o�A�����{���ӯ ����	��-�?��c� u�S�������Ͽ῿� ����'�M�+�=σ� ��w�����m������ %�7��[�m�K�}ߣ� �߳��߷����!��� E�W�5�{��ϱ��� e�������	�/��?� e�C�U����������� ����=O-s ����]��� �'9]oM� ������/� 5/G/%/k/}/[/�/�/ ��/�/�/�/?1?? U?g?E?�?�?{?�?�? �?�?	O�?O?OOOO uOSOeO�O�O�/�O�O �O_)__M___=_�_ �_s_�_�_�_�_o�_ �_7oIo'omoo]o�o �o�O�o�o�o!�o 1W5g�k}� �����/�A�� e�w�U�������я� �o����	�O�a�?� ����u���͟���� �'�9��]�o�M��� ������ۯ��ǯ�#� ůG�Y�7�}���m��� ſ�����ٿ�1�� A�g�E�wϝ�{ύ��� ����	�߽�?�Q�/� u߇�e߽߫ߛ����� ���)���_�q�O� ����������� ��7�I���Y��]��� ������������!3 WiG��}� ���%�A� 1w�g���� ��/+/	/O/a/?/ �/�/u/�/�/�/�/? �/9?K?�/o?�?_? �?�?�?�?�?�?O#O OGOYO7OiO�OmO�O �O�O�O�O_�O1_C_ %?g_y__�_�_�_�_ �_�_�_o�_+oQo/o Ao�o�owo�o�o�o�o �o);U__q �������� %��I�[�9����o� ��Ǐ�����ۏ!�3� M?�i��Y������� ՟�ş����A�S� 1�w���g�����������ӯ�+�=��$D�CS_SGN �QK�c��7m�� 16-MA�Y-19 10:�20   O�l�4�-JANt�08:�38}����� N.DѤ�����������M4�o���Im��P�Zۘq��  O�VE�RSION �[�V3.5.�13�EFLOG�IC 1RK���  	����P�?�P�N�!�P�ROG_ENB � ��6Ù�o�U?LSE  TŇ��!�_ACCLI�M����Ö���WRSTJNT��c��K�EMO�x̘��� ���INIT S.�G�Z����OPT_SL ?�	,��
 	�R575��Y�74j^�6_�7_�50��1��2_�@ȭ��<�TO  Hݷ���V�DEX��d�c����PATHw A[�A\��g�y��HCP_CLNTID ?��6� @ȸ�����IAG_GRP� 2XK� ,`����� �9�$�]�H������1234567�890����S�� |�������!�� ��H���;�dC�S���6�� ���.�R v�f��H�� //�</N/�"/p/ �/t/�/�/V/h/�/? &??J?\?�/l?B?�? �?�?�?�?v?O�?4O FO$OjO|OOE��O y��O�O_�O2_��_�T_y_d_�_,
�B^ 4�_�_~_`Oo�O &oLo^oI��Tjo�o.o �o�o�o�o �O'�_ K6H�l��� ����#��G�2� k�V���B]���Ǐُ �������(��L�B\�Drx�@��P�C����4  �79֐�$�� >���:�����ߟʟܟ����CT_CON�FIG Y��|Ӛ�egU����STBF_TTS��
��b����Û�:u�O�MAU��|�~�MSW_CF6��Z��  �OCoVIEW��[ɭ������-�?�Q� c�u�G�	�����¿Կ ������.�@�R�d� v�ϚϬϾ������� ߕ�*�<�N�`�r߄� ߨߺ��������� &�8�J�\�n���!� �������������4��F�X�j�|����RC£\�e��!*�B^�� ����C2g{��SBL_FAUL�T ]��ި�G�PMSKk��*�TDIAG ^:��աI��UD�1: 6789012345�G�BSP�-?Qcu �������/�/)/;/M/� ��
@q��/$�TR'ECP��

��/ ?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOi/{/xO�/�UMP_OPTIcONk���ATR¢tl��	�EPMEj���OY_TEMP � È�3B��J�P�AP�DUN�I��m�Q��YN_?BRK _ɩ��EMGDI_STaA"U�aQSUNC_S;1`ɫ �FO�_�_�^
�^dpOoo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{�E��� ��y�Q��� �2� D�V�h�z������� ԏ���
��.�@�R� d��z�������˟� ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i����� ����ÿݟ����� /�A�S�e�wωϛϭ� ����������+�=� O�a�{�iߗߩ߻�տ ������'�9�K�]� o����������� ���#�5�G�Y�s߅� ������i������� 1CUgy�� �����	- ?Qk�}����� ����//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?u ?�?�?�?��?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_m?w_�_�_�_ �?�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9Ke_ W����_�_�� ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�]oy����� ���ӟ���	��-� ?�Q�c�u��������� ϯ����)�;��� g�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�_�i�{ߍ� �߹����������� /�A�S�e�w���� ����������+�=� W�E�s������ߧ��� ����'9K] o������� �#5O�a�k} �E������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? GYc?u?�?�?��? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_Q?[_m_ _�_�?�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /I_Sew��_� ������+�=� O�a�s���������͏ ߏ���'�A3�]� o�������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �9�K�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� �������ߑ�C�M� _�q߃ߝ��߹����� ����%�7�I�[�m� ������������ �!�;�E�W�i�{��� ������������ /ASew��� ����3�! Oas������ ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?+=G?Y?k?!? ��?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	_#?5? ?_Q_c_u_�?�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o-_7I[m �_������� �!�3�E�W�i�{��� ����ÏՏ����% /�A�S�e�q����� ��џ�����+�=� O�a�s���������ͯ ߯����9�K�]� w���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� '�1�C�U�g߁��ߝ� ����������	��-� ?�Q�c�u����� ������m��)�;�M� _�y߃����������� ��%7I[m ������� �!3EWq�{� ������// //A/S/e/w/�/�/�/ �/�/�/�/�/+?=? O?i_?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O�? �$ENETMODE 1aj5��  0054_F[�PRROR_PR_OG %#Z%6��_�YdUTABLE  #[t?�_�_��_gdRSEV_N�UM 2R  ��-Q)`dQ_A�UTO_ENB � PU+SaT_NON>a b#[EQ(b_  *��`��`%��`��`4`+�`�o8�o�oZdHIS%c1�+PSk_ALM 1]c#[ �4�l0+�o;M_qȃ��o_b``  �#[aFR�zPT�CP_VER �!#Z!�_�$EX�TLOG_REQ��f�Qi,�SIZ\5�'�STKR�oe��)�TOL  �1Dz�b�A= '�_BWD�p���Hf��D�_DI�� dj5SdDT1<KRņSTEPя�|P��OP_DOt��QFACTORY�_TUN�gd<�D�R_GRP 1e#YNad 	���FP���x̹� ��� ��$�f?�� ���ǖ��ٟ �ԟ���1��U�@� y�d�v�����ӯ�����LW
 J�n��,��tۯ�j�U����y�B�  B�������$  A@<��s�@UUUӾ��������E�� E��`F@ F�5�U/�,��L����M��Jk��Lzp�JP���Fg�f�?� � s��9�Y9�}�9��8�j
�6��6�;���A����O ��� �� I �������[FEAT?URE fj5���JQHan�dlingToo�l � "
P�Englis�h Dictio�nary�def�.4D St��ard�  
�! hAnalog I/OI׿  !
IX�g�le Shift�I�d�X�uto �Software� Update � rt sѓ�ma�tic Back�up�3\st���ground� Edit��f�d
CamWera`�Fd�e���CnrRndIm����3�Comm�on calib� UI�� Eth�e�n��"�Mon�itor�LOA�D8�tr�Relgiaby�O�ENS��Data Acq�uis>��m.f�dp�iagnos���]�i�Docum�ent ViewyeJ��870p��ual Chec�k Safety�*� cy� �han�ced Us��F�r����C �xt�. DIO :�f�i�� m8���en]d��ErrI�L���S������s  t� Pa�r[�� ����J944�FCTN Men�u��ve�M� J9�l�TP InT�f�ac{�  744���G��p Mas_k Exc��g�� R85�T��Proxy Sv��  15 J�i�gh-Spe��S�ki
� R738�Г��mmuni�c��ons�S R7��urr�T�d��022��aю�connect 2�� J5��Incr���stru,Қ�2� RKARE�L Cmd. L���ua��R860~hRun-Ti��EnvL�oa��K^U�el +��s���S/Wѹ�7�Li�cense���r�odu� ogBo�ok(Syste�m)�AD p�MACROs,>��/Offs��2�NDs�MH��9 ����MMRC�?�ޙ�ORDE� ec_hStop��t? n� 84fMi$�,|� 13dx��]�p��׏���Modz�_witchI�VP��?��. sv<��2Optm�8�2��fil��I ��z2g 4 !+?ulti-T������;�PCM gfunY�Po|����4$�b&Regir� r �Pri���FK+7���g Nu�m SelW  �F�#�� Adj9u���60.��%�|� fe���&tatu�!$6���%���  9 J6�RDM Robo}t)�scove2�� 561��Rem�U�n@� 8 (|S�F3Servo���ҩ�)SN�PX b�I�\d�cs�0}�Libr<1��H� �5б f�0��58��S�o� tr�ssag�4%G 91�p Ȓ�&0���p/Iތ�  (ig TM�ILIB(MӋ�Fgirm����gd7����s�Acc�����0�XATX�Hel	n��*LR"1���Spac�Arqu>z�imulaH��ѹ Q���Tou�Pa��I��T��c���&��ev. f.�svUSB �po��"�iP�a��  r"1Unexcept��`0i$�/����H59� VEC&�r��[6����P{��RcJPRIN<�V�; d T@�TSP CSUI՚� r�[XC��#W�eb Pl6�%d# -c�1R�@4dp�����I�R66?0�FV�L�!FVGrid~K1play C�`lh@����5RiR�R�.@���R-35i�A���Asci�i���"��� 51�f�cUpl� � �(T����S��@r�ityAvoid�M �`��CE��r9k�Col%�@�GuF� 5P��j}P�����
 B�L�t� W120C C� o���!J��P��y��� �o=q�b @DCS- b ./��c��O��q��`�; ���q�ckpaboE4�D�H@�OTШ�mai'n N��1.�H��Gan.��A> aB!GFRLM���!i ��~�MI Dev� s (�1� h8j��spiJP��� �@��D�Ae1/�r���!hP� M-2� i��߂^0i�p6�P}C��  iA/'�?Passwo�qT�ROS 4����q�eda�SN��ClAi����G6x Ar��� 47�!���5s��DER��Tsu�p>Rt�I�7 (9M�a�T2DV�
�3D Tri-���&��_8;�
�A�@Def?����{Ba: deRe p 4t0��e�+��V�st64MB �DRAM�h86�΢FRO֫0�A;rc� visI���n��7| ), <�b�Heal�wJ�{\h��Cell`�2�p� �sh[���� Kqw�c� - ��v���p	VCv�t�yy�s�"Ѐ6�ut��v�m��"�xs ���TD_0��XJ�m�` 2��a[��>R tsi�MA3ILYk�/F2�h�|�ࠛ 90 H��(F02]�q�P5'����T1C��5����FC��U�F9�Gig�EH�S�t�0/A� cif�!2��boF��dri=c ��OLF�S����" {H5k�OPT �򆧊49f8���cCro6��@��l�A�pA�Syn.(RSS) 1L�\1y�rH�L� (2x5�5��d�pCVx9����e�st�$SР��> \�pϐSSF�e$�tex�D o���A��	� BP���a�(R;00�Qirt��:���2)�D��1�e�V}Kb@l Bui, 9n��WAPLf�į0��Va�kT�XCG�M��D��L����[CcRG&a�YBU��YKfL��pf��k�7\sm�ZTAf�@�О�Bf2�и��V�#�s���� r���CB���
f���W�E��!��
���T�p��DT�&4 1Y�V�`��EH�����
�61Z��
�R�=2�
�E (Np��F��V�PK�B���#��GHf1`?G���H��р?I�e ����L�D�L��N��7\@s@���`���M��Odela<,��2�]M�� "L[P� �`?��_�%�����5S��-F�TSO��W�J57��VG�F�|�VP2֥ 5\b�`0&�cV:����T;T� �<�c�e,?VPD���$T;F��DIu)�<I�a\so<"��a-�6Jc6s6�4L��M�V9R�h���T�ri�� ���5�` �f@�@�������P
� �����`��Img PdH�[l��I/A  VP�S��U��Ow��!%S�Skast�dpn)ǲt�� S�WIMEST�BFfe�00��-Q� �_p�PB�_�Rued�_�T�!�_�S ��_bOH573o2c2��-oNbJ5N�Iojb)�	Cdo�cxE��o�_�l p��o�TdP�o�c�B�o r�2.rٱ(Jsp�EfrSEo�f1�}Ξr3 RGoeEL	S��sL����s�� ���B	��S\ $�F�3ryz�ftl�o~�g�o���������?�����P  �n�&�"�l ��T�@<�^�蒐Y��e�u8Z���alib��Γ��ɟ3����埿�\v ��e\c�6�Z�f�T�v�'R VW���8S��UJ91����i�ů[c�91+o�w8���847�:��A4�j���Q��t6�m���vrc.����HR����ot�0ݿ��  d��8ޯ�460�f>eS0L�97��0�U�ЄϦ�60.� g �н�+��'�ܠ�Ϻ��8co��DM߱U"������ߕpi�߲T!� ��na;�� @���u%��ⅰI�loR�d��1a5a9gϱŭ���95����R����1��?��o��#��1A�/���vt{�UWeǟ���ￇ�73[���7�ρ�C3 W��62K�=f	R���8��������d����2�ڔ�����@�@" "http�����t87 �� v R7��78����4�� ��TTPT�#	���ePCV4/v߀�jL�Q�Fa7��$N�0�/2�rIO�)/;/M/N6.sv3�64i�o|S�l? torah?p*�|`�?��AM/�?�
??.?0�k/��1 �JO��� ,O�tro����[P��OB4c.0K?�g'�)�24g?��� (B�Od�\i�OA5sb�?U_�?vAi�/i��/�/Wn��`�o%�Fo�4l�$opf��oXF I)xoΚcmp\7��mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@����naO��4*O0wi��%P�?"�bsg@?�]7�YEM���8wo2VJ�/ե11?o��3DMs�BC��!7J�\���(�52�XFGa AP�ڟ<�v�`/şaqs����'/Of��1�	9�VRK���ph�fքH5+�=�IN/�¤SkiW�/�I�F��_�%��fsH�I�O�l����"<�`���$�`����\jԿ8z5bO�vrouς�93(�ΤH (DϮ� �?sG��|��F�Ou��������D)O��*�3 P$�FӅ�k��ϻ���럴� �PL��ʿ���pbox�ߦeboL���Sh �>�R.�b0wT{����fx6 ��P��D��3��#_&I\m;YEe�OԆ�M�hxW�=Ete,���dct\���O$AkR������Xm*���ro3��D�l��j9��V'�  FC���|@�քy f?6KARE0�_�~ (Kh��.ccf���WpoO�_K�up��a���<H/j#- Eqd/�384���$qu�o�@�/ o2o?Vo<�7C�)�s�NJԆ�|?�3l\sy�?�40�?�Τwio�u]?�w58�?,F�$OJ�
?&Ԇ"io�!�V��u&�A��PR�ߩ5,� s��v1\  H552B��Q21p0R{78P510.R�0  nel �J614Ҡ/WATUP��\d8P545*�H8R�6��9VCAuM�q97PCRImP�\1tPUIF�C8Q2?8  ingsQy0X��4P P63P @P� PSCH��D�OCVڀD �PCS�U���08Q0=PqpV?EIOCr���v P54Pupd�P�R69aP���PSET�pt\hPQ`Qt��8P7`Q�!MA�SK��(PPR�XY���R7B#PO�CO  \pppb36���PR�Q��b�1Pd60Q$cJ53�9.eHsb��v�LCH-`(�O�PLGq\bPQ0t]`��P(`HCR��t4`S�aund�P'MCSIP`e0aPle�5=Ps�p(`DSW � �  qPb0`�aPa��(`PRQ`Tq�RE`(P�oa601P<cPCM�PHcR0@q\j23b�V�`E`�S`UPvisP`E` c�`�UPcPRS	a�bJs69E`sFRDmP�sRMCN:eH9y31PHcSNBARan�rHLB�USM�q�c�Pg52�fHTyCIP0cTMIL�eh"P�`eJ �PA�P�dSTPTX6p967PTEL�p��P�`h�`
Q8P8$Q48>a0"PPX�8P95�P`�[�95qqbUEC�-`F
PUFRhmPfahQCmP90ZQ�VCO�`@PVI�P%�537sQSU�IzVSX�P�SWE�BIP�SHTTIPthrQ62aP�!tP�G���cIG؁�`c��PGS�eIRC�%��cH76�P�e� Q�Q|�Ror��R5�1P s:P�P,t53�=P8u8=Py�C�Q6�]`�b�PI��q52]`sJ56E`s��L�PDsCL�qPt5�7\rd�q75UP c�R8���u5P sR55]`,s� P8s���P�`CP�PP�SJ7]7P0\o�6���cRPP�cR6�ap0�`�QtaT�79P`�364�Pd87]`�d90P0c��=P,����5�9ta�T91P�� ��1P(S���Qpa�i�P06=P- C
�PF�T	���!aLP� PTS�pL�CABR%�I БIQ` ;��H�UPPaintPM�S�Pa��D�IP|�S{TY%�t\patP�TO�b�P�PLSR76�`�5�Q��Wa�NN�Paic�qN9NE`�ORS�`�cwR681Pint'�'FCB�P(�6x�-�W`M�r��!(`OB^Q`plug�`L�awot �`OPI-���PSPZ�PPGڤQ7�`73ΒPRmQad�RL��W(Sp�PS��n�@��E`�� �PTS-�� W��P�`�apw�`��P`cFsVR�PlcV3D%��l�PBVI�SAP�L�Pcyc+PAP�V1�pa_�CCG^IP - U��L�Pwrog+PCCR�`��ԁB�P �PԁK�=�"L�P��p��(h�<�P��h�̱�@g�=Bـ
TX�%�n��CTC�ptp��<2��P927"0ҝP�s2�Qb��TC-�r�mt;�	`#1ΒT�C9`HcCTE�Peurj�EIPp.p/��E�P�c��I�useZ��Fـvrv�F%���TG�P� CP��%��d -h�H-�Tr�a�PCTI�p��T=L� TRS���p��@נ��IP�PTh�Mn%�lexsQTMQ`�ver, �p�SCp:���F��Pv\e�PF�IPSV"+�H�$c�j�ـtr�aCTW8-���CPVGF-��S�VP2mPv\fx����pc�b��e��bV=P4�fx_m��-���SVPD-��SVP]F�P_mo�`V�Z cV��t\��LmP�ove4��-�sVKPR�\|�tPV�Qe5.W`V6�*u"���P}�o`���`��CV�K��N�IIP��CV�����IPN9�Gene���D��D�R�D(����  ��f谔��pos.��inaEl��n��DeR��d�`��d�P��omB���on,���R�D�R��\��TXf��D$b���omp�� "NȔ�P��m���! ��=C-f����=�FXU�����g �F��(��Dt IIД�r�D��u�� "x����Cx_ui 0X������f2��h	Crl2��D,r9�ui�Ԣ� it�2c�0co��e�"����ا(.{)� ���� ﯶ� IQn�Q �I[ ���_= wo���,bD� ���|GG� �����4 ��e� vʷ�� ��&� 2��Z uz������� ��TW�&q~q 5��޷&�o? ;0{��  �2� ��y� ����W&��� ?Ȼ3� A��ew�/> �\�3&�T��� 77߽� ���� �w��� ֵ��&8 �l1���S�) ��{�d *J� �F's ~���� 6:0� ���,��s�- Q��v� ���� �,�T �Z�BLx6���6 ݀�6���Pa�r ��s>�E��j�6dsq��F  ��������ЁDhel������ti-�S�� �Ob��Dbc`f�O�����t OFT��P<A�_�V �ZI��D��V\�qWS|��= dtle�E�an�(bzd��t�itv�Z�z�Ezt XWO H6�6܋��5 H�6H6�91�E4܀TofksqtF� Y682��4�`�f804�E9�1�g�`30oBkmo�n_�E��eݱ�� wqlm��0 J�f�h��B�_  ZD�TfL0�f(P7�EcklKV� �6|�ƁD85��ّ�m\�b����xo�k�ktq��g2.g���y�LbkLVts��IF�bk������I�d I/f��GR8� �han�L�`�Vy��%��%ere�����io�� ac.�- A�n�h��.�cuACl�_�^Cir��)�g��	.�@�& G��R630���p v�p�&H�f���un��R57v�OJavG�`Y���owc��-AS�F��O��7���S�M�����
afN��rafLa�Qvl�\F c�w a�`��?VXpoV �30���NT "L�FFM ��=����yh	a�G-�uw�� �m2.��,�t��̹�6lԯ��sd_�MC'VČ���D���fsl�m�isc. � H552�2��21&dc.pR78�����0�708J�614Vip OATUu�@�OL�w545ҴINTL��6�t8 (V�CA���sse�CRI��ȑ��U�I���rt\rL�2�8g��NRE��.�f,�63!��,�S�CH�d Ek�DO#CV���p��C,�<��L�0Q�isp��EcIO��xE,�54�����9��2\sl,�SET���lр�7lt2�J7�Ռ?MASK��̀?PRXY҇�ҹ7���OCO��J�6l�3�l�� (SVl�A�H�L�@Օn��539Rsv�v��#1��LCH����OPLGf�ou�tl�0��D��HC]R
svg��S@��h��CSa�!�{�50��D�l�5!�lQ��DSW��S����̀���OP����7��P�R���L�ұ�(Ssgd���PCM�Զ�R0 \s��5P՝���0���n�qԋ AJ�1��N�q�2���PRSa���69��� (AuF�RD�Խ��RMC�N���93A�ɐC�SNBA�F9N� HLB��� M���4���h�2A�95�z�HTCaԈ�TM;IL6�j95,��o857.,PA1��ito��TPTXvҴ JK�TEL���piL�� XpL�80�I)��.�!��P;��J95��s "N����H�UEC��77\cs�FR��<Q���C��57\{VcCOa�,���IP1�jH��SUI�	C�SX1�AWE9Ba��HTTa�8�R62��m`��G�P%�IG %tut�KIPGSj�| R�C1_me�H7�6��7P�ws_�+�?x�R51�\�iw�N���H�53�!��wL�8!�h�R66��H���Ԡ�8��@;J56��1�P��N0��9�j��L�F��R5`%�A|�5qԉr�`,�8 5��{16�5!��@�"5��H84!�29��0��P�J���n B[�J377!Ԩ�R6�5h3�n���y36P��3R6 ��-`;о Ԩ@��wexeKJ87���#J90!�stu�+�~@!䬵�k90�kop�B���D�@!�p�@|BA�g*�0n@!��Q��06!�@"[�F�FaP�6��́v,�TS� NC[ЗCAB$iͰl1I��R7��@q�y�wCMS1�rog+Q1M�� �� TY$x�wCTOa�nv\+���1�(�,�6�co�n�~0��15��JNN�%e:��P��9GORS%x���8A�w815[�FCBaUnZQ�P!��p{��C�MOB��"G��O�L��x�OPI�$\�lr[�SŠ�T	D7��U��CPRQR9R	L���S�V�~`����K�ETS�$1��0����3�Ԩ�FVuR1�LZQV3D$� ���BVa�SAP�L1�CLN[�PV��	rCCGaԙ��sCL�3CCRA�/n "W!B�H�7CSKQn\0�pX��)�0CTPn����Qe��p!$bCt�aT0U�pCTC��yЋRC1�1 (<�s��trl,�r��
TX��TCaersrm�r�MC"�sܡ�#CTE��nr5r�REa�XPj�^���rmc�^�a"��P�QF!$���$p� "�rG1�tTG�$c8��QH�$SC�TI�! s��C;TLqdACK�Rpt)��rLa�R82���M��YPk�.���OF ��.���e�{�CN���^�1�"M�^�aԀС�Q`US��!$��M�QW�$m�VGFޑ$R MH��P2�� H5� ΐq���ΐ�$(MH[�VP��uoY����$)��Dv��hg��VPF��"MHG̑`e!�+�V/vpcm�N���p��N��$�VPRqdL)��CV�x�V� `"�X�,�1�($TIa��t\mh��K��eCtpK�A%Y�VP%�ɠ�!PN���Ge{neB�rip�����8��extt���Y�m�"� (��HB���)�� x�������Ȣ�res.�yA�ɠ�n����*���p��@M�_�NĀ6�L���Ș�yAv`L�Xr�Ȉ2��"R;ʎȽ\ra��	P�� 7h86��Gu+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr�Ȩ2��L�1��n2�h� �0XL�XR}�RI{�e� L�x���c�Ș����N�vx�L��"��2\�r�]�N�82�d ���b�ɉa��y1��/��k�@���A��ruk8�ʘ L�sop��H��}�ts{�����sx��9��j965���Sc��h��5 JI9�{�
�PL�J	ween��t I[
.x�com��Fh�L��4 J��fo.��DIF+�6�Q����rati|��p�ڙ1�0�
R8l߾�M �����P��8� �j�mK�X�HZ��$��N�oڠ�ș3�q��vi���890�~�l Sl�yQ���tpk�xb�j �.�@�R�d������,/n(�8�8�0����
:�O8�<�Q}�C�O���PT��O (��.�Xp|�~H���?��v �wv���8�22�pm���7322��j7�^Ϙ@ƙ���cf�=Yv9r���vcu�� �O�O�O�O_#_5_7�93Y_��wv4{_��_w�ʈ�ust_�_�cus�_�Z�� oo,o>oPo�io���nge��(pLy747�jWelʨHM;47ZKEq {����[m�MFH�?�(wsK�8J�n����o��fhl;��wmf���? :�}(�4	<g J{��I�I)̏މw��X�7c74kﭏ/7ntˏ2݊e+���se�/�Caw��8�ɐ��EX �\�!+: �p��~�0e0��nh�,:Mo+�<xO��1 "K�O��\a��#0��.8����{h�L?�j+�mo�n�:��t�/�st�?-�w�:���)�;੬(=h�;
d Pxۻ�{:  ���c �J0��re��}��STD�!�treLAN�G���81�\tq�d�������rc�h.������htwv�WWָ�� R79��"Lo�51 (�I�W�ph�Ո�4�aww�� �vy �62�3c�h a?�ctAi�֘!�X�iؠ�t ��n,�։�����j��"AcJP@�3p�vr{��H�6��!��- S�eT� E3�) G�J�934��LoW�4 (S������ <���91 ��8!4�jA9�所+���y�
��v	�btN�ite{�R ��I@Ո����� P�������	 ����Z�vol��X ��9�0<�I�p���ld*���F�864{��?��K�	�k扐�֘1^�wmsk��M�q�Xa�e�����p��0RBT��1ks.OPCTN�qf�U$ RTCamT��y�� U��y��U��UlU6L�T�1Tx��D��SFq�Ue�6T���USP W�b# DT�qT2h�T��!/&+��TX�U\j6&�U U�UsfdO&�&ȁ�T���662DPN�bi��%�Q�%62V��$���%�� �#(�(6To6eG St�%��#5y��$�)5(To�%tT0�%5�W6T���%�#�#orc��#I��8�#���%cct�6ؑ�?�4\W6965q"p6}"�#\j536����4�"�?kruO O,Im?Np�C ��?t�0<O�;�ea �%���?
;gcJ7� "AV�?�;av�sf�O__&_8WtpD_V_0GT�F|_:U�cK6�_�_r�O�3e�\s�O2^y`O:�m�igxGvgW! m��%��!�%T�$E �A{6�po6��#37N�)5R5_2E���$�0���$Ada�Vd ���V�?;Tz7�_�e7�DDTF9���#8��`�%��4y�ted Z@�A}�@�}�04N�}�}���}�#dc& }����u �6�v��v1�u1\�b�u$2}���}� R�83�u�"}��"}�v�alg���Nrh �&�8�J�Y�o�ue��� j70�v=1���MIG�uerfa ��{q���E�N�ءEYE�ce A���񁏯pV�e�A! ���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b��T��/E In�B�  8W�|��537g��.��(MI�t�Ԇ1r��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y��ac���2���Rɏ �jo��2�� dj�d�8r}� og\�k�0��g��wm�f�Fro/� E�q'�4"}�3 J8��oni[���0�}Ĵ�� o� ��$ʛ��m@�R�e��{n�Д�V�o�������  ����=⣆"POS\��<��ͯ menϖ��6��OMo�43��� ��(Coc� An`[�t���"e�a\�v�p��.��cflx$�le��8�hr�trv�NT� CF+�x E/�t	qi�M��ӓxc��p�f�lxX����Z�cx��
0 lh��h8��mo���=� H���)� (�vSER,���g�0߆0\r�vX�= ���I � - �t�i��H��VC�8�28�5��L"�RC��n G/���w��P�y�\v�vm "o�lϚ�x`��=e�:ߠ-�R-3?������vM [�AX/2��)�S�rxl�v#��0��h8߷=� RAX�A�����9�H�E/Rצ�����h߶"RXk��F��˦85��2L/��xB885_�q�R�o�0iA��5\rO�9�K��v����q8���.�n "�v��88��8s�i ?� 9 ��/�$�y O�MS"���&�9�R H74&�`�745�	p��p��y'cr0C�c�hP0� j�-�a%?o��6D9;50R7trl��wctlO�APC����j�ui"�L��� � ����^ࣆ!D�A��qH��&-^7���� λ�616C�q�7914h���� M�ƔI��99��(���$FEAT_�ADD ?	����Q%P  	�H._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������������ &8J\n���������TD�EMO fY   WM _������� �//%/R/I/[/�/ /�/�/�/�/�/�/�/ ?!?N?E?W?�?{?�? �?�?�?�?�?�?OO JOAOSO�OwO�O�O�O �O�O�O�O__F_=_ O_|_s_�_�_�_�_�_ �_�_ooBo9oKoxo oo�o�o�o�o�o�o�o >5Gtk} �������� :�1�C�p�g�y����� ��܏ӏ���	�6�-� ?�l�c�u�������؟ ϟ����2�)�;�h� _�q�������ԯ˯ݯ ���.�%�7�d�[�m� ������пǿٿ��� *�!�3�`�W�iϖύ� ������������&�� /�\�S�eߒ߉ߛ��� ��������"��+�X� O�a��������� ������'�T�K�]� ���������������� #PGY�} ������ LCU�y�� ����/	//H/ ?/Q/~/u/�/�/�/�/ �/�/???D?;?M? z?q?�?�?�?�?�?�? 
OOO@O7OIOvOmO O�O�O�O�O�O_�O _<_3_E_r_i_{_�_ �_�_�_�_o�_o8o /oAonoeowo�o�o�o �o�o�o�o4+= jas����� ���0�'�9�f�]� o���������ɏ��� ��,�#�5�b�Y�k��� ������ş����(� �1�^�U�g������� ��������$��-� Z�Q�c����������� ��� ��)�V�M� _όσϕϯϹ����� ����%�R�I�[߈� ߑ߫ߵ�������� �!�N�E�W��{�� ������������ J�A�S���w������� ������F= O|s����� �B9Kx o������/ �/>/5/G/t/k/}/ �/�/�/�/�/?�/? :?1?C?p?g?y?�?�? �?�?�? O�?	O6O-O ?OlOcOuO�O�O�O�O �O�O�O_2_)_;_h_ __q_�_�_�_�_�_�_ �_o.o%o7odo[omo �o�o�o�o�o�o�o�o *!3`Wi�� ������&�� /�\�S�e�������� ������"��+�X� O�a�{���������� ߟ���'�T�K�]� w����������ۯ� ��#�P�G�Y�s�}� �������׿��� �L�C�U�o�yϦϝ� ���������	��H� ?�Q�k�uߢߙ߫��� �������D�;�M� g�q���������� 
���@�7�I�c�m� �������������� <3E_i�� �����8 /A[e���� ����/4/+/=/ W/a/�/�/�/�/�/�/ �/�/?0?'?9?S?]? �?�?�?�?�?�?�?�? �?,O#O5OOOYO�O}O �O�O�O�O�O�O�O(_ _1_K_U_�_y_�_�_ �_�_�_�_�_$oo-o GoQo~ouo�o�o�o�o �o�o�o )CM zq������ ���%�?�I�v�m� ��������ُ��|�;�  2� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as��������'9  :>Ugy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w����� ����я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ �������(/=C6Y k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ������/�A��$FE�AT_DEMOIoN  E��q���>�Y�INDE�Xf�u��Y�IL�ECOMP g�������t�T���SETUPo2 h����?�  N ܑ���_AP2BCK �1i��  �)B���%�C�>���1�n�E����)� ��M�˯�������<� N�ݯr������7�̿ [��ϑ�&ϵ�J�ٿ Wπ�Ϥ�3�����i� �ύ�"�4���X���|� ��߲�A���e���� ��0��T�f��ߊ�� ����O���s����� >���b���o���'��� K���������:L ��p����5�Y �}�$�H�l ~�1��g� � /2/�V/�z/	/ �/�/?/�/c/�/
?�/ .?�/R?d?�/�??�? �?M?�?q?O�?O<Ot���P� 2�*.VRCO�O�0*�O�O�3�O�O�5�w@PC�O_�0F'R6:�O=^�Oa_�KT���_�_&U�_�\�h�R_�_�6*.F�zOo�1	(SoElx�_io�[STM �b��o�^+P�o�m�0�iPendant? Panel�o�[H�o �g�oYor�ZGIF|��e�pOa��ZJPG ��*��e���z��JJS�����0@���X��%
JavaSc�riptُ�CS�ʏ1��f�ۏ %�Cascadin�g Style ?Sheets]��0�
ARGNAME�.DT���<�`\@��^���Д៍�АDISP*ן���`�$�d��V�e��C?LLB.ZI��=��/`:\��\������Collabo�鯕�	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V� 9���ϝ�$�4i����V���zό�!ߘ�TP�EINS.XML�(�@�:\<����C�ustom To�olbar}��PASSWORD��~�>FRS:\���� %Pass�word Config��?J���C� ��"O��3�����i��� ��"�4���X���|�� ���A���e����� 0��Tf���� �O�s��> �b�[�'�K ���/�:/L/� p/��/#/5/�/Y/�/ }/�/$?�/H?�/l?~? ?�?1?�?�?g?�?�?  O�?�?VO�?zO	OsO �O?O�OcO�O
_�O._ �OR_d_�O�__�_;_ M_�_q_o�_�_<o�_ `o�_�o�o%o�oIo�o �oo�o8�o�on �o�!��W�{ �"��F��j�|�� ��/�ďS�e������ ���T��x������ =�ҟa������,��� P�ߟ񟆯���9��� �o����(�:�ɯ^� ����#���G�ܿk� }�ϡ�6�ſ/�l��� ��ϴ���U���y��  ߯�D���h���	ߞ� -���Q߻��߇��,���$FILE_D�GBCK 1i������� ( �)
�SUMMARY.�DG,���MD:�`����Dia�g Summar�y���
CONSLOG��y����$����Consol�e log%���	?TPACCN���%g�����TP �Accounti�nF���FR6:�IPKDMP.ZIP����
��)�����Excepti�on-����MEMCHECK�������8�Memor?y Data���LN�)�RI�PE���0��%� Pack�et LE���$ySn�STAT*�#� %~LStatus�i	FTP�/��/�:�mmen�t TBD=/� �>)ETHERNE�/o�/�/���Ethern�U<�figura�L��'!DCSVRAF1//)/B?�0� verify �allE?�M(=5DIFF:? ?�2?�?F\8diff��?}7o0CHGD�1�?�?�?LO X�?sO~3&�
I2BO8)O;O�O bO�O�OGD3�O�O�OT_� �O{_
VUPDATES.�P��_��FRS:\��_�]��Upda�tes List��_��PSRBWLOD.CMo���R�o�_9�PS_RO�BOWEL^/�/:GIG��o>_�o��GigE ��n�osticW�N��>�)�aHADOW�o�o�ob��Shadow ?Change���8+"rNOT�I?=O��N?otific�"���O�A�PMIO�o��h��f/���o�^U�*�UI`3�E�W��{�UI������B���f��_� ������O������� ��>�P�ߟt������ 9�ί]�򯁯�(��� L�ۯp������5�ʿ ܿk� Ϗ�$�6�ſZ� �~��wϴ�C���g� ��ߝ�2���V�h��� ��߰���Q���u�
� ���@���d��߈�� )��M��������� <�N���r����%��� ��[����&��J ��n��3�� i��"�X� |��A�e� /�0/�T/f/��/�/�/=/�/�/�$�$�FILE_�PPR��P��� �����(MDONLY 1i5~�  
 �z/ Q?�/u?�/�?�?t/�? ^?�?O�?)O�?MO_O �?�OO�O�OHO�OlO _�O_7_�O[_�O_ �_ _�_D_�_�_z_o �_3oEo�_io�_�oo �o�oRo�ovo�o A�oew�*� �`����&�O�~�*VISBCK,8|1;3*.VDV�|���FR:\o��ION\DATA�\��/��Vi�sion VD filȅ��&� <�J�4�n������3� ȟW������"���F� ՟�|������m�֯ e������0���T�� x������=�ҿa�s� ϗ�,�>���b��� ϗϼ�K���o��� ��:���^����ϔ��*�MR2_GRP �1j;�C4�  B�}�	 �71������E�� �E�  F@ F�5U�������L���M���Jk�Lzp��JP��Fg�f�?�  S�����9�Y9}��9��8j
��6��6�;֞�A�  ���BmH��B���B���!$����������<���@UUU#��� ��Y�D�}�h������� ��������
C��_CFG k;T M����]�NO :�
F0� � \�R�M_CHKTYP  0�}�00�0��OM_MsIN	x���5v0X� SSBd]l5:0���bx�Y���%TP_DEF_OW0�x�9�IRCO�M��$GENOVRD_DO*�62�THR* �d%d�_ENB�� �RAVCr��mK�� ��� ��/3�/��/�/n�� �M!OUW -s��}��ؾ��8�g�;?�/x7?Y?[?  C��0ý���(7�?�<B�?B����2��*9�.N SMTT#t[)���X�4�$HOST�Cd1ux�̹�?�� MCx��;zOx�  �27.0�@1�O  e�O�O	__-_ ;Z�O^_p_�_�_�LN_�HS	anonymous�_�_�_oo"1o yO��FhFk�O �_�o�O�o�o�o�o J_'9K]�o�_ �����4o�Xo joG�~�o^������� ŏ�����1�T� ��y���������� �,�>�@�-�t�Q�c� u���������ϯ�� �(�^��M�_�q��� ��ܟ� �ݿ��H� %�7�I�[Ϣ�ϑϣ� �����l�2��!�3� E�Wߞ���¿Կ���� 
�������/�v�S� e�w��������� ����+�r߄ߖ�s� ����߻��������� ��'9K]����� �����4�F�X� j�l>��}��� ���//1/T ��y/�/�/�/�/.D~\AENT 1v
;� P!J/?  ��/3?"?W?? {?>?�?b?�?�?�?�? �?O�?AOOeO(O�O LO^O�O�O�O�O_�O +_�O _a_$_�_H_�_ l_�_�_�_o�_'o�_ Koooo2o{oVo�o�o �o�o�o�o5�oY .�R�v��zQUICC0���3��t14��"�����t2��`�r�ӏ!ROUTERԏ���#�!PCJ�OG$���!1�92.168.0�.10��sCAMgPRTt�P�!d�11m�����RT폟������$NAME �!�*!ROB�O���S_CFG� 1u�) ��Auto-started/FTP&��= ?/֯s����0�B� �f�x���������S� �����,������ ���ϼ�ޯ�������� �ʿ'�9�K�]�oߒ� ߥ߷���������SM%y�{�U� �ό���������� 
��.�@�c���v���0���������z�%� 7�I�K�8�\n� ��k����� 3�FXj|�� ��a��7 /M*/</N/`/r/9 �/�/�/�/��/�/? &?8?J?\?�m?�� �?�//�?�?O"O4O �/XOjO|O�O�O�?EO �O�O�O__0_w?�? �?�?�O�_�?�_�_�_ �_o�O,o>oPoboto �_o�o�o�o�o�o K_]_o_L�o�_�o� ����o� ��$� 6�Y�Y�~��������ƏZ�_ERR �w3�я�PDUS_IZ  g�^�p����>�WRD� ?r�Cq� � guestb�Q�c�u��������`�SCDMNGR�P 2xr����H�g�\�b��K� 	P01�.00 8`� /  � �  � B  ���� ���H�W��L��L��L�����O8�����Xl�����a4�  ��Ȥ� �8����\���)�`�;F�������d��.�@�R�ɛ_GROUUېy������	ӑ���QUPD'  ?u����İ�TYg����T�TP_AUTH �1z�� <!iPendan���-�l���!K?AREL:*-�6�H�KC]�m��U��VISION �SET���ϴ�! �����R�0��H�B߀��f�x��ߜ߮���C?TRL {�����g�
��FF�F9E3��AtF�RS:DEFAU�LT;�FAN�UC Web Server;�)�� ��9�K��ܭ����������߄WR_CONFIG |ߛ� ;��IDL_CPU_PCZ��g�B�I�y� BH_�MINj�)�}�?GNR_IO���g���a�NPT_SOIM_D_������STAL_SCR�N�� ���TPM?ODNTOL������RTY��y����F �ENO���Ѳ]�OLNK 1}��M�������|�eMASTE���ɾeSLAVE �~��c�O_CcFGٱBUO�|O@CYCLEn�>T�_ASG 19ߗ+�
 �� ��//+/=/O/a/�s/�/�/�/�/��N�UM��
@I�PCH�^RTRY_CNZ���@P�������� @kI�+E�z?E��a�P_MEMBE�RS 2�ߙ� 5$���2���ݰ7��?�9a�SDT_I�SOLC  �����$J23_D�SM+�3JOB�PROCN��JOmG��1�+�d8�?��+D�O�/?
�LQ�O __/_�OS_e_w_�_`�O Hm@��E#?>&BPOSREQO��?KANJI_����a[�MON ����b�yN_goyo@�o�o�o�Y�`3�<�� ��e�_ִ��_L����"?`EYLO�GGINLE��������$LANGUAGE ��<T� {q�LeGa2�	�b���g��xP��  �J�g�'��b����>�MC:\RSCH\00\<��XpN_DISP �+G�H��O�O߃gLOCp�Dz����AsOGBOOK �������������X����� Ϗ����a�*��	p�����!�m���!���=p_BUFoF 1�p���2F幟���՟D�� Collaborativǖ��� F�=�O�a�s������� ֯ͯ߯���B�9��K���DCS �>z� =���'�f���?ɿۿ���H@{�I�O 1�� ~?9Ø��9�I�[�m� �ϑϣϵ��������� �!�3�E�Y�i�{ߍ�@�߱��������E��TMNd�_B�T�f� x������������ ��,�>�P�b�t���p����L��SEVD0���TYPN�1�$6���QRS�"0&��<2FL 1�"�J0���������GTP�:pOF�NGN�AM1D�mr�tUP�S�GI"5�aO5��_LOADN@G� %�%DF_MOTN�y�� �MAXUALRM��'���(��_PR�"4F0d��1�B_�PNP� V 2��C	MDR0W771ߕ�BL"�8063%�@ A�_#?�ߒ|/�C���z�6��/���/P�o@P 2��+ ��ɖ	T 	t  ��/�%W? B?{?�k?�?g?�?�? �?O�?*OONO`OCO �OoO�O�O�O�O�O_ �O&_8__\_G_�_�_ u_�_�_�_�_�_o�_ 4ooXojoMo�oyo�o �o�o�o�o�o0B %fQ�u��� �����>�)�b� M�����{�������� Տ��:�%�^�p�S������D_LDXDISApB�MEMO_APj�E ?C
 �,�(�:�L�^�p�������ISC 1�C ����4 �������4��X����C_MSTR ����w�SCD 1���L�ƿH��տ ���2��/�h�Sό� wϰϛ��Ͽ���
��� .��R�=�v�aߚ߅� ���߻�������<� '�L�r�]����� ���������8�#�\� G���k����������� ����"F1jU g������ �B-fQ�u���h�MKCF�G ����/�#L_TARM_��7"0�0N/V$>� METPUᐒ3ۆ���ND� AD�COLp%A {.CM�NT�/ �%� ����.E#>!�/4��%POSCF�'��.PRPM�/9S�T� 1��� 4=@��<#�
1� 5�?�7{?�?�?�?�? �?�?)OOO_OAOSO �OwO�O�O�O�O_�A��!SING_CH�K  �/$MODAQ,#����.~;UDEV 	���	MC:o\HS�IZEᝢ��;UT�ASK %��%�$1234567�89 �_�U9WTR_IG 1���l3%%��9o��"ocoFo5#F�VYP�QNe��:S�EM_INF 1��3' �`)AT&FVg0E0po�m)�a�E0V1&A3&�B1&D2&S0�&C1S0=�m)�ATZ�o;"tH@?g�a[o�xA�@�z���� �o >��o'��K�� �����я:�L� 3�p�#�5���Y�k�}� �����$�[�H��� ~�9�����Ưد���� ����ӟ�V�	�z��� ����c�Կ����
�� .���d��)�;��� ��q�������˿<� ��`�G߄ߖ�IϺ�m� ϑϣ����8�J�� n�!ߒ�M�������h_NITOR� G� ?�[   	?EXEC1�/�U25�35�45�55�T�P7�75�85�9�0�Қ�4��@�� L��X��d��p��@|�������2��U2��2��2��2��U2��2��2��2U23��3��3@��;QR_GRP_S�V 1��k (��A�z�4�~��K������?�K:z�j]�Q�_D��^�PL_NAME !3%�,�!Def�ault Per�sonality� (from FwD) �RR2�� 1�L6(L�?�,0	l d������� �//(/:/L/^/p/ �/�/�/�/�/�/�/ZX2u?0?B?T?f?x? �?�?�?�?\R<?�? �?O O2ODOVOhOzOp�O�O�OZZ`\R��?�N
�O_\TP �O:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o Ho_)_~o�o�o�o�o �o�o�o 2DV hz�[omo��� �
��.�@�R�d�v����������Џ� �Ef  Fb�� F7���   #��!��d�� @�R�6�t�������l���ʝ����� ݘ����"�@�F��d���� "𩯹�ݐ�A�  ϩU[��$n�B�E� �� � �@D�  �?��� �?�@��A@��;f��FH� ;��	l,�	 |䒑j�s�d�>倀� ��� K(���Kd$2K ���J7w�KY_J˷�ϜJ��	�ܿ�� @I����_f�@�z���f�γ�N�������	Xl���������S�ĽÔ��I �����5��� � ����A?oi�#�;����� ���l�  �Ϫ�-���ܛG�G�Ѳ5��@n�@a �  �  ���ܟ*�͵	'�� � H�I�� �  ��Рn�:�Èl�ß�=��̈́�в@�ߚЕ����/�"����̷NP�  ',���-�@
�@����?=�@A���B�O  Cj�a�Be�yCi��#�B�޸�ee��^^ȹBР��P��`��̠�����ADz՟ �n�3��C�i�@�R�pR�Y����  �@o� ���  ���?�ff������n� ɠ#ѱy 9G
(���I�(�@u�P~����t�t���>�����;�Cd;���.<߈<��g�<F+<L �������,�d�,��̠?fff?��?�&&��@��@�x��@�N�@���@T�H �ِ�!-�ȹ�|� �
`������� //</'/`/r/]/�/��eF���/�/�/��/m?��/J?�(E��G�#�� FY�T?�?P?�?�?�? �?�?O�?/OO?OeO k��O�IQOG�?�O 1?�OmO_0_B_T_������A_�_	_��_�_�_ o��A��A0n0 bФ/o C�_Uo8�_�Op��؃o�o��o�o���W����v�oC�E� q�H�d��؜a@q���e�F�BµWB]��NB2�(A���@�u\?��D�������b��0�|�uR�����
x~�ؽ���Bu*C��$�)`�$� ���GC#����rAU�����1�e�G�D�I�mH��� I:�I��6[F���C��I��J��:\IT�H
?~QF�y��p��*J�/ I�8Y�I��KFjʻCe�o��s� ����Џ���ߏ�*� �N�9�r�]������� �����۟���8�#� \�G�����}�����گ ů���"���X�C� |�g�����Ŀ����� ��	�B�-�f�Qϊ� uχ��ϫ�������� ,��P�b�M߆�qߪ� ���߹�������(�� L�7�p�[����������s($���3�:����$���3Ï��d�,�4���@�R�wa����xl�~�wa���e��<��wa4 �{�������(L:ueP�P~�A�O�������	����G2W}h ������/�@��O�O7/m/[(d=� s/U/�/�/�/�/�/?��/1??U?C?y?�= � 2 Ef9gF[b��77�9fB)a,a)`C9A`�&`w`@-o�?w`e�O)O�?MO�Ow`�?�?�O�O��O�O9c?�0�A7hJt4w`w`!w`xn
 �O9_K_ ]_o_�_�_�_�_�_�_��_�_o#ozzQ ���h��G���$�MR_CABLE� 2�h ��a�T� @@��0�Ae��a�a�a���`��0�`C�`�aO�8�tB�n��d��`�aE�4��E�#�o�f#��0��0�DO���By`������bED4�E�c,��o�g8�  ���C�07n�d4
vے�0� �b��XE�Z&�l�`y`
q�C�p�bHE�
v{#g�5D�Ү�qz�lҠ`��0�q�p�b0�
v�%c����b=%	E;h��u/o�c-��4t H�\�?�9�K�]�o�ԏ Ϗ��
�ɏۏ@���?�:�eo �a����������b����� �����`�	 ����@������%� �*�0�6� ��ݐ�����`��	������@������*�,� ,�-�\cOM ��ii��3�� �  ( �%% 23456�78901i�{� �f�����������1�����
��`��not sen�t3�����;��TESTFEC�SALGR  eH�qiG�1d.�š
:�� �DCbS�Q��c�u��� 9UD�1:\maint�enances.Gxml��ֿq� �=��DEFAULT-�i4\b�GRP 2�M� � =��a�{�p  �%Fo�rce�sor check  ��
�b�z��p����h5-[ �ϻ������ϖ��D�%!1st c�leaning �of cont.� v�ilatiCon��}�Rߗ+��@[�ߔߦ߸����mech�cal,`������0��h5k�@�R�d�v������(�rolle _Ƶ����/����(�:����Ba�sic quarterly��������,����������M�F�M��:C@"Gp P�a�b`i4��� ����#C���M"��{Pbt����Supp~q�grease���?/&/8/hJ/\/��C+ ge��_. batn�y`/��/h5	/�/�/�/`? ?_�ѷen'�!v��/�/��/��?`�?�?�?�?�G=?O�qp"CrB1O��0�/`OrO�O�O�O�Xt$��Lf��C-m��A�O:�OO$_6_H_�Z_l_�t*cabYl�Om���S<m��Q�_:�
_�_�_o o0oo)(Ӂ/�_�_���_�o�o�o�o�o�;O@hau1�l�2r xm�<qC:��op�������ReplaW�f Uȼ2�:�._4� F�X�j�|�m�$%��� o�������#���
�� .�@���d���ŏ׏�� ��П����U�*�y� ����r���������	� q��?�߯c�8�J�\� n���ϯ�����ڿ)� ���"�4�Fϕ�jϹ� ˿������������ [�0�ϑ�fߵϊߜ� ������!���E�W�,� {�P�b�t����߼� ����A��(�:�L� ^������������ �� $s�H���� ��q�����9 ]o�Vhz� ��U�#�G/ ./@/R/d/��/�/� �//�/�/??*?y/ N?�/�/�?�/�?�?�? �?�???Oc?u?JO�?�nO�O�O�O�O+J�r	 H�O�O__6M2_ @OBE:_p_>_P_�_�_ �_�_�_ o�_�_oHo o(oZo�o^opo�o�o��o�o�o �o :z� �bA?�  @�q _����Fw�� �H* �** @q>v�p 2T�f�x�:�������ҏ��eO^C7�Տ #�5�G�	�k�}���ُ ���c�����W�� C�U�g���ß)����� ӯ���	��-�w��� ��9�������m�Ͽ���=�O�E	A�$�MR_HIST �2�>uN�� 
� \$�Force se�nsor che�ck  1234?567890q�3�����ß�N�}SB� -3�19.8 hou�rs RUN 9�.�Y�!1st �cleaning� of cont�. ventilation0Äϖ�Ԩ�-�Y���me;ch��cali�%���4��o�DN��t��95��1�|���rolleh��+�=�O��Y�B�asic qua?rterlyߒ� �߶�
O4�F��(�� ����b�t������ �����M�_����:�����p���:�SKCFMAP  >u�Q��r5�������ONREoL  .��3���EXCFEN���:
��QFN�CXJJOGOVLIM8dNá ��WKEY8��_PAN7����ԧ�����SF?SPDTYPxC���SIG�:��TO1MOT�G���_CE_GRP [1�>u\�D �����/Ⱥ� �/�/U//y/0/ n/�/f/�/�/�/	?�/ ???�/c??\?�?P? �?�?�?�?�?O)OO�MO,���QZ_ED�IT5 )TCO�M_CFG 1����[�O�O�O 
>�ASI �y3�!
__+[_O_ċ�>O�_bHT_/ARC_Uք�T_MN_MOD�E5�	UAP�_CPL�_gNO�CHECK ?^�� �� o .o@oRodovo�o�o�o �o�o�o�o*!�NO_WAIT_�L4~GiNT�A���EUwT_ERMRs2���3��Ʊ J�����>_)�V�|MO�s��}x:O�v���8�?������ l��rPA�RAM�r�����j���5�5�G� =  r�b�t�s� X������������֟0�0����b�t������SUM_RSPACE�����Aѯ�ۤ�$ODRDS�P�S7cOFFS?ET_CARt@�_��DIS��PE?N_FILE:�7��AF�PTION�_IO��q�M_�PRG %��%�$*����M�WOR�K �yf ���춍����������	 �������gT��R�G_DSBL  ���C�{u��R�IENTTO7 f��C� A ��UT_SIM_D�y���V�LCT ��}{B �<٭��_PEX�P=�n�RAT�W dc���UP ���`���e�w�]߬�ߩ��$�2r��L6(L?�>��	l d���� ��&�8�J�\�n�� ������������� "�4�F�X���2�߈� ������������*�<w�Tfx� ������J`�ˣG���Tz�Pg�� ����/"/4/F/ X/j/|/�/�/�/�� �/�/??0?B?T?f? x?�?�?�?�?�?�?�? �/�/,O>OPObOtO�O �O�O�O�O�O�O__`(_:_��O��y_�]2ӆ��_�^�_�_ �W^]^]��/ooSog�Hgrohozo�o�o �o�o�oF`�#|`�A�  9y�����OK�1�k������<o�EA�nq? @D�  �q��4��nq?��C��s�q|1� ;�	l���	 |�Q�s��r�q>��u ��sF`H<zH~��H3k7GL��zHpG��99l7�k_B�T�F`SC4��k�H���t���-�Ae���k������s��� � �ሏ����EeBVT���dZ�џ���ڏ ���q-�Fk�y�{jFbU���n@}6�  ����z�Fo��Be	'�� � ��I� �  �:p܋=���ڟ웆�@���B�,�D��B���g�AgN����  '|���g���B��p�BӀC�׏����@  #��Bu�&�ee^�^^މB:p 2���>�m�6p�Z���Dz?o}�܏�������׿������Ǒ��� ~f�  � �M�z��*�?�ff�_8�J�ܿ 3pϑ�ñ8�Чϵʖq.·�	(����P���'��s��tL�>��/�;�C�d;��.<���<�g�<F+<L ��^oiΚr�d@��r6p?fff�?�?&�п�@���@x��@��N�@���@T싶�Z���ћtމ �u�߈w	�x��ti�>� )�b�M��q����� ��������:�%�^��������W���S�E��  G�aF�� Fk��������� 1U@yd�� ����q��	�� {�A��h����D�a��ird��A{�/w/J/5/n/vA�A���":t�/ C�^/�/Z/ ލ?����/�/1??���Wҵ���g��pE�! ~1�?04�0
1ή1@IӀ��B���WB]�NB2��(A��@��u\?��������������b�0�|�uR����
�>��ؽ��B�u*C��$��)`�? ����GC#����rAU�����1�eG���I��mH�� I�:�I�6[Fߍ��C4OI���J�:\IT��H
~QF��y�Ol@�*J��/ I8Y�I���KFjʻC ��-?�O�O__>_)_ b_M_�_�_�_�_�_�_ �_o�_(oo%o^oIo �omo�o�o�o�o�o  �o$H3lW� {������� 2��V�h�S���w��� ��ԏ�������.�� R�=�v�a�������П ����ߟ��<�'�`� K�]���������ޯɯ���&�8�#�\��3(�J���3:a���9���J�3��c4������������1�����ڿ��1����e���14 �{2�2�r�`ϖτ�(�Ϩ��%PR�P���!�h�!�K�6�o�Z�����u�|ߵ� �����������3�� W�B�{�f�4���������d�A����!�� 1�3�E�{�i��������������  2 �Ef�7Fb�7���6B�!�!� C9� �� �0@�/`r@������#x�@�+=�3?, TV�8v��0�0���0�.
  D�����// %/7/I/[/m//�/�:� ��ֻ�G����$PARAM�_MENU ?�2�� � DEFP�ULSE�+	W�AITTMOUT��+RCV? �SHELL_W�RK.$CUR_oSTYL� 4<�OPTJJ?PTB�_?Y2C/?R_DECSN 0�Ű<�?�? �?�?�?OO?O:OLO�^O�O�O�O�O�O�!S�SREL_ID � .�����EUS�E_PROG �%�*%�O0_�CCC�R0�B���#CW_H�OST !�*!HT�_=ZT��O_�S�h_zQ�S�_<[_TGIME
2�FXU� ?GDEBUG�@�+��CGINP_FLgMSKo5iTRDo�5gPGAb` %l��tkCHCo4hTY+PE�,� �O�O �o#0Bkfx �������� �C�>�P�b������� ��ӏΏ�����(��:�c�^�p�����7eW�ORD ?	�+
? 	RSc`��/PNS��C4�sJOv1��TE�P�COL�է�2�Z�gLP 3������OjTRACEC�TL 1�2�.�! ��Ғ�|��q�DT Q�2��Ǡ��D � ��ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� �����Я0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~�T �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�?��3�$PGTRA�CELEN  ��1  ����0��6_UP ����A�@�1@�1_�CFG �E��3�1
@�<D�0<DZO<C�0uO$B�DEFSPD e�/L�1�0��0�H_CONFIG� �E�3 ��0�0d�D��2 	�1�APpDsA�A�0ۂ�0IN'@TROL �/MOA8pE�QPE�E��G��A<D�AILI�D(C�/M	bTGR�P 1ýI �l�1B  ������1A�33�FC� F8� _E�� @eN	�A��AsA�Y�Y�A�@� 	 vO�Fg�_G ´8cokB;` baBo,o>oxobo�o�1�>о�?B/�o�o~�o =%<��
C @yd��"������  Dz @�I�@A0�q� ����� ��ˏ���ڏ���7� "�4�m�X���|���Ú�)ґ
V7.1�0beta1HF� @����A�q��Q  6�?� �BܠP��p �C��&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@���f�������ҡ�R��ܣ�Rљ���1��i������t�<B!CeQKNOW_�M  lE7FbTSoV ĽJ�B oC_�b�t��������������1�]aSM�S�.�K ���	NB�0?���ĿK�|��-�bb� �A�RP����0��X���bQMR�S��T�iN���d���V]{ST�Q1 1�K
 4MU�iǨj� K�]�oߠߓߥ� ��������2��#�h� G�Y��}�������
������,�27�I��1�<t�H��PA3^�p�����,�4��������,�5(:,�6Wi{�,�A7����,�8�p!3,�MAD�6� F,�OVLD  KD�xO.��PARNUM  ��MC/%�SCH
� E
9'!G)�3Y%UPD/��E�/>P�_CMP_��0�@�0'7E�$ER/_CHK�%5H�&��/�+RS���bQ_#MO�+?=5_'?O��_RES_G6�� :�I�o�?�?�?�?O �?O7O*O[ONOOrO@�O�O�{4]��<�? �Oz5���O__|3  #_B_G_|3V b_�_�_ |3� �_�_�_|3� �_ �_o|3Oo>oCo|2�V 1�:�k1!��@c?�=2THR_INRc0i!}�o5�d�fMASS�o �Z�gMN�o�cMO�N_QUEUE C�:�"�j0��O�N� U1Nv�+Dp�ENDFqd?`yEX1Eo`u� BEnpP>AsOPTIOMwm;�DpPROGRAM7 %$z%Cp}o�(/BrTASK_I���~OCFG ��$��K�DAT5A��T���j12/ď֏������ +�=�O�a��������x��͟��INFO�͘��3t��!�3�E� W�i�{�������ïկ �����/�A�S�e�Pw�����Θ� '�ضFJ�a K_N��8T��˶ENBg ڽ�w1��2��GN�2��ڻ P(O��=���]ϸ��@���v� ��u�uɡdƷ_EDIT �T�����G�WERFL�x�c)��RGADJ �^��A�  $�?j0�0��a�Dqձӆ5?�?��ʨ�	<u�)%e�������FӨ�2�R��	HJ;pl�G�b_�>�p�Aod�t$��*�/� **:@�j0�$�@�5Y�T���^��q�߈b~� L��\�n����� ����������4�F� t�j�|����������� ��bLBT� x����:�� $,�Pb�� �/����/~/ (/:/h/^/p/�/�/�/ �/�/�/V? ??@?6? H?�?l?~?�?�?�?.O �?�?OO O�ODOVO �OzO�O_�O�O�O�O �Or__._\_R_d_�_@�_�_�_�_�_�f	g� io�pWo�o{d�o��~o�ozoB�PR�EF �Rږp��p
�IORIT�Y�w[���MPDcSP�q��pwUT6�|���ODUCT3������OG��_TG��8��ʯr�TOENT 1���� (!AF�_INE�p,�7��!tcp7�_��!udN���!�icmv��ޯrX�YK�ض���q)�� ,�����p� �&�	��R�9�v�]� o�����П�����ퟐ*��N�`�*�sK���9}�ߢ���Ư B,�/6쒯���������At�,  �Hp��P�b�t����u��w�HANCE C�R��:�wd��连�2s�9Ks���PORT_NUM��s�p���_CARTREP{p|�Ω�SKSTA�w� d�LGS)��ݶ��tӁpUnothing��������{��TEM�P ޾y��'e���_a_seiban�o\��olߒ�}� �ߡ���������"�� �X�C�|�g����� ���������	�B�-� f�Q���u��������� ����,<bM �q��������(L�VER�SIyp�w} �disable�dWSAVE �߾z	2600/H768S?��!ؿ����/ 	�5(�r)og+^/y�e@{/�/�/�/�/�*�,D/? �p���_�p� 1�Ћ� �����Wh?z?��W*pURGE��B��p}vgu,�WF�0DO�vƲ�vW%��4(��C�WRUP_DE?LAY �\κ5�R_HOT %�Nf�q׿GO�5R_NORMAL&H�r6O<�OZGSEMIjO�O|�O(qQSKIPF3	��W3x=_98_ J_\_]�_�_{_�_�_ �_�_�_�_	o/oAoSo owoeo�o�o�o�o�o �o�o+=aO q������� �'��7�]�K��������)E�$RA{����K/�zĀÁ_PoARAM�A3��Kw @.�@`�6�1�2C<��y���C�6$�BÀB�TIF�4`�RCV�TMOUu�c�]�ÀDCRF3��I� �+UC��AqD��2=\��(?��]�w
�ޅ���4���+_���;�Cd�;��.<߈�<�g�<F+<L���Ѱ��d�u�L�������ϯ� ���)�;�M�_����RDIO_TYP�E  M=U�k�E�FPOS1 1�N\�
 x4/��� ��+�$/<��$υ� pϩ�D���h��ό�� '������o�
ߓ�.� ��Rߌ�������5� ��Y���i��*�<�v� ��r���������U� @�y����8���\��� ��������?��c��^��2 1�KԿ�X�T�x��3 1����n�Y�S4 1� '9K�/�'/�S5 1����/�/�/�/:/S6 1�Q/c/u/�/-??|Q?�/S7 1��/��/
?D?�?�?�?d?S8 1�{?�?�?�?�WOBO{O�?SMASK 1L��O�D�GXNO���F&�^��MOTEZ�Ż��Q_ǁ�%]pA݂���PL_RANG�!Q]�_QOWER ��ŵ�P1VSM�_DRYPRG �%ź%"O�_�UT?ART �^�ZUME_PRO�_��_4o��_EXEC?_ENB  ��#�e�GSPD`O`Wh�ՅjbTDBro�jR�M�o�hINGVE�RSION �Ź#o�)I_A�IRPURhP ��O(�MMT_�@T�P#_ÀOBOT�_ISOLC�N�TV@A'qhuNAM�E�l��o�JOB_�ORD_NUM �?�X#qH768  j1wZc@�r�r�V�s��r�;?�r?�r�p�ÀPC_TIME�u�a�xÀS232�>R1�� L�TEACH PENDANw�:GX��!O Ma�intenanc�e Consj2䊏��"��No UseB�׏�������1�C�y�V�NPqO�P@�YQ�c�S�CH_L`��%^ �	ő��!�UD1:럒�R�@VAIL�q@�Ӏ��J�QSPACE�1 2�ż ���YRs�i�@Ct�YR�Ԁ'{��8�?��˯����"��� 7�2�c�u�����G��� ߯ѿ򿵿�(��u �AC�c�u�����Ͻ� ߿���ϵ��(��=� _�qσϕ�C߹����� �߱��$��9�[�m� ߑߣ�Q������߭� �� ���	�W�i�{�� ��M�������5��� .S�e�w�����I �������* ?as��E�� ���/&//;/] o������/2/ �/?"?�/7?Y/k/}/ �/�/O?�/�/�?�?�?�O0OOKA��*�SYPpM*�8.�30261 yB5�/21/2018� A �WPfG|��H�_TX`� !$COMME�$USAp� $ENAB�LEDԀ$IN�N`QpIOR�B�@R�Y�E_SIGN_4�`�AP�AIT�C�B�WRK�BD<�_T�YP�CRINDX�S�@W�@%VFRI�{�_GRPԀ$�UFRAM�rSRT�OOL\VMYHO�L�A$LENG�TH_VTEBTI�RST�T  �$SECLP�XUFINV_POS�@�$MARGI~�A$WAIT�`f�ZX2�\�VG2�GG1�AI�@�S�Q	g�`_WR�BNO_U�SE_DI�BuQ_�REQ�BC�C]S$CUR_TCQP��R"a^f �GP_�STATUS�A @ �A3`�BLk�H$zc1�h�P@����@_�FX ��@E_MLT_�CT�CH_�J�`CMO�@OL�E�CGQQ'$W�@w�b#t�DEADLOCK�uDELAY_C�NT�a3qGt�a$~wf 2 R�1[1$X<�2[2
�{3[3$Zwy�q%Y��y�q%V�@�c�@�b$iV�`�RV�UV3oh|>b�@ � �d��0arMSKJ�Lg�WaZ�C`NRK�PS_oRATE�0$����S
`�Q�TAC��P#RD���e�S*��a�4�b  �DG�A� 0�P�flp bquS2ppI�#`
`��P 
�S\` � �A�R_E�NBQ �$�RUNNER_A)XI�<`ALPL�Q�R�U�THICQ$�FLIP7��DTF�EREN��R�IF'_CHSU�IW��%V)�G1����$Př�A�Q�Pݖ_JF��PR_P�	�R�V_DATA�A�  $�ET�IM���$VAL�U$�	�OP_ �  �A � 2 �SC�*�	� �$ITP_!�SQ]PNPsOU}�o�TOTL��o�DSP��JOGsLIb��PE_PKpRc�Of�i��PX]P�TAS�$KEPT_MIR��¤"`�M�b�APq�aE �@�y�q�g@١c�q�;PG�BRK6�x�t��L�I��  ?�pSJ�q�P�ADEz��ܠBSOCz�MO�TNv�DUMMY{16Ӂ$SV�`�DE_OP��SFSPD_OVR
����@LD����OmR��TP8�LE���F������OV��S!F��F����bF�d��ƣ&c)�fQc�LCH�DLY��RECOQV���`��W�PM���gŢ�RO������_\F�?� @v�S ��NVER�@�`OFeS�PC,�CSWDٱ�c�ձ���B����TR�G�š�`E_FD}O��MB_CM}���B��BLQ�¢	�dQ�̄Vza�BUP�dg��G
��AM�`��@`KՊ�e�_M!��d�AMf�Q��T$SCA����DF����HBKd�v���IO�U��I'R��PA ����������p��і�?DVC_DB�S!�@x�Q�!�s�d�9�1A���9�3A��ATIEO�0��͠��US����WaAB��R+c��`tá`DؾA��_A�UXw�SUBCP	UP���S�`����3��жc���3�FLA<�B�HW_Cwp"��Ns&�]sAa��$/UNITS�M�F�ATTRIz�Z��CYCL�CNEC�A���FLTR_�2_FI��TARTUPJp����A���LP������_SCmT*cF_F�F_P����b�FS��+�K�CHA/Q��*�d�RSD��Q����Q�v��_TH�PROr���հEMPJ���G�9T� �Q�DI�@y�RAI�LAC/�bMX�L!Of�xS��ځ����X�����PR#�S`a�pp�C� =	��FUNC���RIN`QQP� fԱRA)]R ��pAƠ��AWAR֓F��BLZaWrAkg�ngDAQ�B�rkLD�र&q�dM�K���TI����j��$�@RIoA_SW��AF��Pñ#��%%�p9r�1��MOIQ���D�F_~P(�PD"L�M-�FA�PHRD]Y�DORG�H; �_QP�s%MULS�E~Pz���*�� J⼺Jײ��FAN?_ALMLVG��!�WRN�%HARD�P��UcO�� K2$SHADOW]��kp�a02��� STOdf�+�_^�w�AU{`�R��eP_SBR �z5���:F�� �3_MPINF?�\�8�4��3REGV/1DG�+cVm �C�C�FL(��?�DA`iP���Z`�� ������Z�	 �P(Q]$�A$Z�Q V�|@�[�
� ���EG߀o���kAAR���㌵2�axG��wAXE��ROB���RED��W�QD�_�Mh�SYA��AF��FS�GWRI�P~F&��STR����E�˰E"H�)��D�a\2kP�B6P��=V��Dv�O�TO�1)���AR�YL�tR�v�3���F�I&�ͣ$LINQKb!\��Q�_3S���E��QXYZt2�Z5�VOFF��R�R�R�XxPB���ds�G�cF�I�03g�������_J��'�ɲ�S&q�R0LTV[6���aTB�ja�"�bC���DUt�F7�TUR� !X��e�Q�2XP���gFL�E���x@�`��U9Z8���� 1�	)�K��Mw��F9���劂����ORQj��G;W3���#� Ґd ���uz����1�t'OVE�q_�M��ё ?C�uEC�uKB�v'0�x -�wH��t���&  `��qڠ�B�ё�u�q��wh�ECh����ER��K	�EP����AT�K�6e9e0�W���AXs�'� �v�/�R ����! �� ��P��`��` �3p�Yp�1�p� � �� �� (�� 8� � H�� X�� h�� x�� ������DEBU�$%3�I���RAB���ٱ�sV��� 
d�J、 ��@񘧕�������Q ���a���a��3q��Yq�+$�`%"<�cLAB�0b�u�'�GROh���b<��B_s ��"Tҳ*`�0A�u��u8q�p1}�ANDGp��@�����U��p1�� �р�0�Qθuݸ��PN�T0���SERV9E �Z@ $`EmAV�!�PO�� ����nP!�P@�$!Y@  $>�TRQ�b
=��BG�K�%"2\��� ?_  l��5�ND6ERRVb(�I��qV0`;���TOQ:��7�L�@
�R��e G�%�Q�� <�50F�G ,�`�z�>��RA� 2 �d!�����S� � M��pxU ����O�CuG�  >��COUNT6Q��FZN_CFGF�G 4#��6��TG4 �_�=�����Î�VC/ ���M �"���$6��q ��FA E� &��X�@��ِ����A����AP���P@HEL�0��� 5b`B_wBAS��RSR�6��CSH����1T�Ǌ�2��3��4��U5��6��7��8��}�ROO����P�P3NLEA�cAB)ë n��ACKu�INO�T��(B$UR0� �=�_PU��!0��OU+�Pd�8j��� �V��TPFWD_�KAR��� ��RE�(ĉ P�P�>QUE�:RO�p�`r0P1I� x�j�P�f��6�QSEM��0���� A��STYL�SO j�DIX�&�Ӹ���S!_TMCM�ANRQ��PEN�DIt$KEYSWITCH���k�HE�`BEATmM83PE{@LE��(>]��U��F���SpDO_HOM�# O�@�EF�pPARaB�A#PY�C� �O�!���OV_Mx|b<0 IOCM�d�FQ��h�HK�YA D�Q�7��U�F2��M���p�cFwORC�3WAR�"���k�OM|@ � @S�#o0U)SP��@1�2&3&4�E��T�O��L�<��8UNLOv�D4�K$EDU1  {�SY�HDDNF�� M�BLOB�  p�SNP�X_AS�� 0�@�0��81$SI=Z�1$VA{��ſMULTIP-��# A� � $��� /4`�B�S��0�C���&FRIFBO�S���3�� NF�ODBU P߰�%@3;9(����nZ@ x��SI���TEs�r�cSGL�1T�Rp&�Н3B�<�@�0STMTq�3�Pg@VBW�p�4S�HOW�5@�SV���_G�� 3p$�PCJ�PИ���FBZ�PHSP AW��EP@VD�0WCw� ���A00�� PB XG XG XG$ �XG5VI6VI7VI8*VI9VIAVIBVI� XG�YF�0XGFVH��TXbI1oI1|I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1Y1Y2UIU2bI2oI2|I2�I2�I�`�X�I2p�X�IU2�I2�I2�I2�I�2Y2Y�p�hbI3�oI3|I3�I3�I3��I3�I3�I3�I3��I3�I3�I3�I3�Y3Y4�i4bI4�oI4|I4�I4�I4��I4�I4�I4�I4��I4�I4�I4�I4�Y4Y5�i5bI5�oI5|I5�I5�I5��I5�I5�I5�I5��I5�I5�I5�I5�Y5Y6�i6bI6�oI6|I6�I6�I6��I6�I6�I6�I6��I6�I6�I6�I6�Y6Y7�i7bI7�oI7|I7�I7�I7��I7�I7�I7�I7��I7�I7�I7�I7jY7T��VP� �UD�y"ՠ��
�<A62��t�RN��CMD� ��M5��Rv�]��Q_h�R����e����<�YS�L���  �  �%\2��+4�'��<W�BVALU��b���'���FH�ID_YL���HI��I����LE_��㴦��$0C�SAC�!� h �VE_BLCK��1%�D_CPU5ɧ 5ɀ� �����C�� ��R� " � PaWj��& ��LA�1�SBћì���RUN_FLG�Ś�����ĳ ����������HЃ��ХĞ�TB�C2��# � @ B��e �S�8�=�FTDC����`V���3d�Q�THF������R�L�ESERVE9��F���3�2�E��Н�Xw -$��LEN90��F��f�RA��W"&G�W_5�b�1��дM2�MO-�T%S60U�Ik�0�ܱF�����[�DEk�21LACEi0�CCS#0�� _MA� j��z��GTCV����z�T� ������.Bi�'A�z�'AJh�#EM5���JH��@@i�V�z��с2Q �0&@o�h��JK��VK9��{����щ�J0����JJv��JJ��AAL��P�������4��5��� N1������.�%LD�_�1n0лCF�"% `�G�ROU���1�AN�4�C�#m REQUsIR��EBU�#���6�$Tk�2$����zя #�& �\�APPR� C�� 0�
$OPEN��CLOS�S�t��	i�
��&' �MfЩ���W"-'_MG߱7CB@�pA���BBRK@�NOLD@�0RT�MO_5ӆp1J��P������ ��������6��1��@ 8"�(�� �����x'��+#PATH''�@!6#@!�<#� � '��1SCA���66IN��UCJ�[1Z� C0@UM�(Y � �#�"�����*���*��~� PAYLOA~�J2LؠR_AN^�3L��91�)1�AR_F2LSHg2B4LO4�!F7�#|T7�#ACRL_� �%�0�'�$��H��.��$HA�2FLE�X��J!�) P�2�D߽߫���0>��* :���� z�FG]D����z���%�F1]A�E�G4�F� X�j�|���BE��� ����������(��X �T*�A���@�XI�[�Hm�\At�T$g�QX<� =��2TX���emX�� �����������������+	�J>+ ��-�K]o|�٠A1T�F�4�ELFP�Ԫs�J� *� JE�mCTR�!�ATN��vzHAND_�VB.��1��$,� $8`F2Av�Ƌ�SWu	#-� $$M*0.� ]W�lg��PZ�����A��� 1����:A(K��]AkAz���LN�]DkDzP2Z G��C�ST_K�4lK�N}DY���  A����0��<7]A<7�W1�'��d�@g`�P �������":8J"�. M�2D�%"��H����ASYIMj%0�� j&-��-W1�/_�{8� �$ �����/�/�/�/ 3J<�:9�/�89�D_VI�v����V_UNI�ӛ��cD1J����╴�W<�� n5Ŵ�w=4��9��?H�?<�uc�4�3��2%�H���/�j�L�0�DIzuO��q��k�>0 �`
��I��A��#���@�ģ���@��IPl� �1 � /�M�E.Qp��9�ơT}�PT�;pG �+ �Gt� ���'��T��0 $DU�MMY1��$P�S_�@RF�@  tG b�'FLA@ �YP(c|��$GLB_TP�ŗ����9 P�q��2 XX� z!ST9�� �SBRM M21_�V�T$SV_E�R*0O�p����CL�����AGPO��f�G�L~�EW>�3 4\H �$YrZr!W@�x�A1+�A���"tj� �U&�4 8`yNZ�"�$GI�p7}$&� -� �Y�>�5 LH {���}$F�E��NE+AR(PN�CF��%P�TANC�B	!JO�G�@� 6.@?$JOINTwa?p{pe �MSET>�7  x�E��HQtp�S{r��up>�8�k �pU.Q?�� LOCK_FOV0�6���BGLV�sG�Lt�TEST_X9M� 3�EMP��q���_�$U&@�%�w`24� Y��5Љ�2�d��3��CE�- ���� $KAR��QM��TPDRA8)�����VECn@���IU��6��HE�f�TOOL�C2Vv�DRE IS3ErR6��@ACH��� 7?Ox �Q�2�9Z�H I�  �@$RAIL_B�OXEwa�RO�BO��?��HOWWAR�1�_�zROLMj��:qw��jq� �@ O_Fkp! d�l>��9����R O8B:���@�	""�O%U�;�Һ�3ơ�r|�q_�$PIP��N&`H�l�@��~#@CORDEDd��p >f�fpO�� �< D ��OB ⁴sd���Kӕ����qSYS�ADqR�qf��TCHt�� = ,8`ENTo��1Ak�_{�-$xCq_�f�VWVA��?> �  &���PREV_RT~�$EDITr&_VSHWRkq��(� &R:�v�D��JA��$�a$HEA�D�6�� �z#K�E:�E�CPSPD.�&JMP�L~��0R*P��?��1%&�I��S�rC�pNEx; �q�wTICK�Cb��M�13�3HN��@ @� 1Gu�!�_GPp6��0STY'"xLO��:�2|l2?�A t 
m MG3%%$R!{�=��S�`!$��w`��Ȃճ���Pˠp6SQ�U��E��u�TERyC�qO�TSUtB ����hw&`gw�Q)�pO����@�IZ��{��^�P�R�kюB1XPU����E_DO��, XuS�K~�AXI�@���UR�pGS�r � ^0�&��p_) ��ET�BPm��o���0Fo��0A|����Rԍ��a;�S=R�Cl>@P� �b_�yUr��Y��yU�� yS��yS���UЇ�U�� �U���U�]��Ul[��Y�bXk�]Cm������YRSC�� 7D h�DS~0��fQ�SP���eATހ��A]0,2N�AD�DRES<B} S�HIF{s��_2C�H�p�I��=q�+TVsrI��E"����a�Ce�
��
;�V8W�A��F \��qA��0l|\A@�rC��_B"R{zp�ҩq�T�XSCREE�Gzv��1TINA����t{�c��A�b?�H T1�ЂB��р��I��A��BE�y RRO������ B���� �UE4I ��g�!p�S��R�SM]0�GUNEX0(@~Ƴ�j�S_S�ӆ@��Á։񇣣�ACY򼯂0� 2H�pU�E;�J�����@G+MT��Lֱ�A�нO*BBL_| W�8���K ��0s�OM��LE/r��� �TO!�s�RIGHΓ�BRD
�%qCKsGR8л�TEX�@|����WIDTH��� �B[�|�<��I�_��Hi� L 	8K���_�!=r���R:�_��Y����)O6q�Mg0紐�U��h�Rm��LUqMh��FpERVwD �P���`�N���&�GEUR��F4P)�)� LP��(R	E%@�a)ק�a�!���f �5�6�7�8Ǣ#B�É@���t�P�fW�S@M��USR&�O �<����U�Qs�FsOC)��PRI;Q�m� :���TRIP>�m�UN����Pv��0��f%��'8���@�0 Q���.�AG �0T� �aL>q�OS�%�RPo���8�R/�A�H�L4����U¡�S�U�g��¢5��OF�F���T�}�O�� 1R����ĝS�GUN�->6�B_SUB?���N,�SRTN�`TUg2���mCOR| D�R�AUrPE�TZ�#'��VCC��	3V �AC36MFB1��%d�PG �W �(#��ASTEM�0����0PE��T3�G�X �\ ��M�OVEz�A��AN��� ���M���LIM_X��2��2�� 7�,�����ı�
�BVF�`E�+�~��04Y��IB�7���5S��_Rp� 2���/ WİGp0p���}СP��3�Zx# ���3����A�ݠCZ�DRID����Vy08�90�� De�MY_UBYd���6��@��!q��X��P_S���3��L�KBM,��$+0DEY(#EX�`�����UM_MUb� X����ȀUS��� ���G0`PACI���а@��:��:0,�:����RE/�3qDL�+��:[��/TARG��P�rr��R<�\ d`�H�A��$�	��AR��#SW2 ��-��@�Oz�%qA7p�yRE�U�U�01�,�HK�2]g0�qP�� N� �EAM0GW�OR���MRC]V3�^ ���O�0M�C�s	���|�REF_���x (�+T� ������p���3_RCH 4(a�P�І�hrj�NA8�5��0�_ ��2�����L@��n�@@OU ~7w6���Z��a2[��RE�p�@;0�\�c�a'2K�@S+UL��]��C��0�3^��� NT��L� 3��(6I�(6q�(3� L��Q5��Q5I�]7q��}�Tg`4D`�0|.`0�AP_HUCv�5SA��CMPz��F�6�5�5�0_�aR ��a�1I\!X�9���GFS��ad ���M��0p�UF�_x��B� �ʼ,RO`��Q��'����UR�3#GR�`.�3IDp���)�D�;��A��~�IN��H{D��V@AJ���S͓UW mi=�����TYLO*�5�����bt +�cPA�� �cCACH �vR�UvQ��Y��pj�#CF�I0sFR�XqT���Vn+$HO����P!A3�XBf`�(1 ���$�`VPy<� ^b_SZ313he6K3he12J�eh �chG�chWA�UMP\�j��IMG9uP�AD�iiIMRE��$�b_SIZ�$P���0 ��ASYN�BUF��VRTD�)u5tqΓOLE_C2DJ�Qu5R��C���U��vPQuEC;CUlVEMV �U<�r�WVIRC�aIuVTPG���rv1s��5qMPLAqa��v��V0�c��� C/KLAS�	�Q�"��d  �ѧ%ӑӠ�@}¾�$�Q���Ue� |�0!�rSr�T@�#0! �r�iI���m�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f � >֦3�@Sp��SLOW>�ROBACCE���!� 9�VR�#���p:���cAD�����PAV��j�� D����M_qB"���^�JMPG ��g:�#E$SS�C��F�vPq��h$ݲvQS�`qVN��wLEXc�i T`��sӂ��Q�FLD6 �DEsFI�3��02���:��VP2>�Vj� �A���V�4[`MV_PI s��t���A�@��FI��|�Z��Ȥ������A���A��~�GA�ߥ1 LOO��1 JCB���Xc��^`�#PLANE��R��1�F�c�����pr�M � [`�噴��S���� f����Af��R�Aw�״rtU��pRKE��d�VANC�A��.�� k���ϲ��BR_AA� l ��2� ��p�#����Gm h���O K�$�������kЍ0OU�&A�"A�
p�pSuK�TM@FVIEM 2l ��P=��҇n <<��dK�U�MMYK1P���`D��ACU���#AU��o $��TIT�$�PR����OP��?�VSHIF�r�p`J�Qsԙ�lfOxE$� _R�`U�#����s��q�������G�"G�޵'�T��$�SCO{D7�CNTQ i�l�>a�-� a�;�a�H�a�V���T1�+�2u1��D��ܲ��  � SMEO�Uq��a�JQЖ����a_�R[�r4�n�*@LIQ�AA^/`�XVR��s��n�TL�P�ZABC�t�t�c��
AZIP��u,���LVbcLn"����MPCFx�v�:�$�� ���DMY_LN�������@y�w Ђ(a�u�� MCM�@CbcCOART_�DPN�? $J71D��=NGg0Sg0ΛBUXW� ��UXGEUL|By�X���	��|!Z��x 	���m��YH�Db  y� 80���0EIGH&�n�?(� H��9��$z ���|�,����$B� Kd'���_��L3�RVS�F8`���OVC�2@'�$|�>P&��
q�4��5D�TR�@ �9VD��SPHX��!�{ ,� *<��$R�B2 2 ����C!�  �@ V+| b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/ ?�/�/V(7%3@/R/ d/v/�/6?�/�/�?�?@�?O4OOION;4]? o?�?�?�?SO�?�?�O�_�O0_Q_8_f_N;5 zO�O�O�O�Op_�O_ o8o�_MonoUo�oN;6�_�_�_�_�_�oo %o4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8����� Ǐ=�_�n���R���şx��ڟN;G � џ�
�� ����W�i�{����� ��ï�.�������A��dW�<�N�|� ������Ŀֿ�ޯ� ��0�B�_�R�d�� �϶������������ �*�L�^��rτ�
� �����������&�p8�J�l�~� `ҟ @�з��������-����&�,� ��9�{�����a��� ������������A 'Y����� ����a#�1�
��N;_MO�DE  ��S ��[�Y�AB���
/\/*	|/��/R4CWORK_{AD�	�T1/R  ���� ��/� _INTVA�L�+$��R_O�PTION6 ��q@V_DAT�A_GRP 2,7���D��P�/~? �/�?�9��?�?�?�? OO;O)OKOMO_O�O �O�O�O�O�O_�O_ 7_%_[_I__m_�_�_ �_�_�_�_�_!ooEo 3oioWoyo�o�o�o�o �o�o�o/e S�w����� ��+��O�=�s�a� ������͏���ߏ� �9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_T�IM����� SC�R ��Ƙ_��5�;#U!P"�Z���� �?E�W�i�{����� .�ïկ�����'(+~�T"2F��"�dR�I�Y��2�o+@a얿����)�u�� k0ϴ��_; ��  T� �� �2�D�)�T D��Q�zόϞϰ��� ������
��.�@�R߀d�v߈ߚ�/V凷�����߽���R�;�o ��W�p��
�t���Diz$� �0 � �T"%!�� ����������� ����*�<�N�`�r� �������������� &8J\n�� ������"4FX ��࿁� ������/` 4�=/O/a/s/�/�/�/@�/�/�/�!!/ �0޲ k�ݵu�0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ ok$o6oHo Zolo~o�o�o�o�o1/ �o�o 2DVh z�/5?����� ���&�8�J�\�n� ��������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	���-�?�Q�c�u��� ���`Ò�ϯ��� �)�;�M�_�q�����@����˿ݿ� �����3� ���&2�,��	1234�5678v�h!�B!��2�C
h���0�ϵ��� �������!�3�9ѻ� \�n߀ߒߤ߶����� �����"�4�F�X�j� |�h�K߰��������� 
��.�@�R�d�v��� ����������� *<N`r��� ����&�� J\n����� ���/"/4/F/X/ j/|/;�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�/�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ �?L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o=_�o�o�o�o �o�o 2DVh�z�����h� �����u�o.�@�R����Cz  B���   ���2�&� � _�
~���  	�_��2�Տ����_�%p������ďi� {�������ß՟��� ��/�A�S�e�w��� ������N������ +�=�O�a�s������� ��Ϳ߿���'�9�DK�_������<v��_��$SCR_G�RP 1
�� �� t{ ��� ���	 �����������������_������)�a�����&�DE� �DW8���l�&�G��CR-35iA� 9012345�67890��M�-20��8��C�R35 ��:�
������������� ��:֦�Ӧ�G���&������	��]�o������:���#H���>�����������&���ݯ:� �j����g������B�t����������9A����  @�`���@� ( ?��=��Ht�P
��F?@ F�`z� y������ � $H��Gs^p��B��7� �/�0//-/f/Q/ �/u/�/�/�/8���P�� 7%?����"?W?x-2?<���]?� H�1�?t�ȭ7��������?-4A , �&E@�<�@G�	B-1 3OZOlO-:�HA�H�O�O|O P�B(�B�O�O_���EL_DEFAU�LT  �����`SHOTSTR#]A7R�MIPOWERFOL  i�/UYToWFDO$V /U�RRVENT 1�����NU �L!DUM_E�IP_-8�j!?AF_INE#P�_�-4!FT�_->��_;o!��`o ��*o�o!RPC_OMAIN�ojh�vo��o�cVIS�oii���o!TPpP�U�Ydk!
�PMON_PROXYl�VeZ�2r��]f��!R?DM_SRV��Y9g�O�!R��k���Xh>���!
�`M���\i���!R�LSYNC�-9�8֏3�!ROS̽_-<�4"��!
�CE4pMTCOMd���Vkn�˟!	��OCONS̟�Wl����!��WASR�C��Vm�c�!N��USBd��XnR� ��Noӯ�������!���E��i�0���WR�VICE_KL �?%�[ (%SVCPRG1��D-:Ƶ2ܿ�˰3�D	�˰4,�1�˰5T�DY�˰6|ρ�˰7�� ��˰�����9����ȴf�!�˱οI�˱ ��q�˱ϙ�˱F��� ˱n���˱���˱�� 9�˱��a�˱߉�� 7߱��_������ ��)����Q���� y��'���O���� w������� ��˰��İd�c�� ����=( as^����� �/�/9/$/]/H/ �/l/�/�/�/�/�/�/ �/#??G?2?k?V?}? �?�?�?�?�?�?O�? 1OCO.OgORO�OvO�O �O�O�O�O	_�O-_��_DEV �Y��MC:5X��`GTGRP �2SVK ��bx 	� 
 ,�PK 5_�_�T�_�_ �_o�_'o9o o]oDo �ohozo�o�o�o�o�o �o5{�_g� �������� �?�&�c�u�\����� ��Ϗ���J\)��� M�4�q���j�����˟ ݟğ��%���[� B��f������ٯ�� �����3��W�i�P� ��t���ÿ���ο� ��A�(�e�L�ί�� RϿ��ϸ������ � �O�6�s�Zߗߩߐ� �ߴ������'�~ϐ� ]���h������ �������5��Y�@� R���v���������@� 	��?&cu\ ������� �;M4qX�� �����/�%// I/[/B//f/�/�/�/ �/�/�/�/�/3??W? �L?�?D?�?�?�?�? �?O�?/OAO(OeOLO �O�O�O�O�O�O�O�O�_"Ud �NLy�6 * 		S=>��+c"_�VU@Tn_Y_B����B�2�J�j�~Q´~_g_�_�Q%�JOGGING��_�^7T(?VjZ��Rf��Y��A�/e�_%o7e�Tt�] /o�o{m�_�o�m?Qi �o�o;)Kq%��o�}os�� ����9�{`�� )���%���ɏ���ۏ �S�8�w��k�Y��� }���ş���+��O� ٟC�1�g�U���y��� ����'����	�?� -�c�Q���ɯ����w� ��s����;�)�_� ����ſOϹϧ����� ����7�y�^ߝ�'� ��ߵߣ�������� Q�6�u���i�W��{� ������=��M��� A�/�e�S���w����� �������=+ aO������u� ��9']� ��M����� �/5/w\/�%/�/ }/�/�/�/�/�/=/"? 4?�/?�/U?�?y?�? �?�??�?9?�?-OO =O?OQO�OuO�O�?�O O�O_�O)__9_;_ M_�_�O�_�Os_�_�_ o�_%oo5o�_�_�o �_[o�o�o�o�o�o�o !coH�o{� �����; �_ �S�A�w�e������� я���7���+��O� =�s�a������П� ����'��K�9�o� ������_���[�ɯ�� �#��G���n���7� ��������ſ���� a�Fυ��y�gϝϋ� �ϯ�����9��]��� Q�?�u�cߙ߇ߩ��� %���5���)��M�;� q�_���߼��߅��� ����%��I�7�m��� ����]����������� !E��l��5� ������_ D�we��� ��%
//��� =/s/a/�/�/�/��/ !/�/??%?'?9?o? ]?�?�/�?�/�?�?�? O�?!O#O5OkO�?�O �?[O�O�O�O�O_�O _sO�Oj_�OC_�_�_ �_�_�_�_	oK_0oo_ �_co�_so�o�o�o�o �o#oGo�o;)_ Mo����o� ���7�%�[�I�k� ���������ُ� ��3�!�W���~���G� i�C����՟���/� q�V������w����� ���ѯ�I�.�m��� a�O���s�������߿ !��E�Ͽ9�'�]�K� ��oϑ�����Ϸ� ���5�#�Y�G�}߿� ����m���i������ 1��U��|��E�� ��������	���-�o� T������u������� ����G�,k���_ M�q���� ���%[I m���	��� //!/W/E/{/��/ �k/�/�/�/�/	?? ?S?�/z?�/C?�?�? �?�?�?�?O[?�?RO �?+O�OsO�O�O�O�O �O3O_WO�OK_�O[_ �_o_�_�_�__�_/_ �_#ooGo5oWo}oko �o�_�oo�o�o�o C1Sy�o��o i�����	�?� �f�x�/�Q�+���Ϗ �����Y�>�}�� q�_�������˟��� 1��U�ߟI�7�m�[� }����ǯ	��-��� !��E�3�i�W�y�ϯ ��ƿ�������� A�/�eϧ���˿UϿ� Q���������=�� dߣ�-ߗ߅߻ߩ��� �����W�<�{��o� ]���������/� �S���G�5�k�Y��� }��������������� C1gU���� ��{����	? -c���S�� ����/;/}b/ �+/�/�/�/�/�/�/ �/C/i/:?y/?m?[? �??�?�?�?? O?? �?3O�?COiOWO�O{O �O�?�OO�O_�O/_ _?_e_S_�_�O�_�O y_�_�_o�_+oo;o ao�_�o�_Qo�o�o�o �o�o'ioN` 9������ A&�e�Y�G�i�k� }�����׏���=�Ǐ 1��U�C�e�g�y��� �֟���	���-�� Q�?�a���ݟ��퟇� �ϯ��)��M��� t���=���9���ݿ˿ ��%�g�Lϋ��� mϣϑϳ�������?� $�c���W�E�{�iߟ� �߯������;���/� �S�A�w�e������ �������+��O� =�s������c����� ������'K��r ��;������ �#eJ�}k �����+Q"/ a�U/C/y/g/�/�/ �//�/'/�/?�/+? Q???u?c?�?�/�?�/ �?�?�?OO'OMO;O qO�?�O�?aO�O�O�O �O__#_I_�Op_�O 9_�_�_�_�_�_�_o Q_6oHo�_!o�_io�o �o�o�o�o)oMo�o A/QSe�����%{,p�$S�ERV_MAILW  +u!��+q~�OUTPUT��$�@�RV� 2�v  $�� (�q�}��SA�VE7�(�TOP1�0 2W� d? 6 *_�π(_������#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u����������Ͽݷ��Y�P��'�FZN_C�FG �u�$�~����GR�P 2�D� ?,B   A[�+q�D;� B\���  B4~�R�B21��HELL���u��j�k��2�����%RSR �������
�C�.�g� Rߋ�v߈��߬������	���-�?�Q��  �_�%Q���(_���,p��⦼�ޖ�g�2,pd�����HK 1�� ��E�@�R� d��������������� ��*<e`r����OMM ������FTOV_�ENB�_���HO�W_REG_UI��(�IMIOFW�DL� �^�)WAIT���$V�1�^�NTIMn���VA�|_)_UNIT����LCTRY�B�
�MB_H�DDN 2W� 2�:%0 �pQ/ �qL/^/�/�/�/�/�/��/�/�"!ON_ALIAS ?e�	f�he�A?S?e? w?�:/?�?�?�?�?�? OO&O8OJO�?nO�O �O�O�OaO�O�O�O_ "_�OF_X_j_|_'_�_ �_�_�_�_�_oo0o BoTo�_xo�o�o�o�o ko�o�o,�oP bt�1���� ���(�:�L�^�	� ��������ʏu�� � �$�Ϗ5�Z�l�~��� ;���Ɵ؟����� � 2�D�V�h�������� ¯ԯ���
��.�ٯ R�d�v�����E���п ���ϱ�*�<�N�`� r�ϖϨϺ���w��� ��&�8���\�n߀� �ߤ�O���������� ��4�F�X�j�|�'�� �����������0� B���f�x�������Y� ��������>P bt����� �(:L�p ����c�� / /$/�H/Z/l/~/)/ �/�/�/�/�/�/? ?�2?D?V?]3�$SM�ON_DEFPR�O ����1 �*SYSTEM*�0m6RECAL�L ?}9 (� �}8copy� virt:\o�utput\tc�pserv3.p�c md: ov�er =>370�27840:35�7235  .8�7.149.�015172]?O+M�4�frs:orde�rfil.dat��4tmpback�\=>147�89�308�?+O�O-N/��2mdb:*.*�TOfOoO�O_$_7D3x?D:\�OIP�O�@��O_�_�_;@4?Ua G_Y_�Et_�_o)o<O NO�O�Oo�o�o�OUo �Opo�o%8_�_�_ n_ ���_GY�_ ~�!�4oFo�ojo� �����o�o_��oz�� �0B�f������ ��Q��v�������
xyzrate 61 ʟܟ� �ȑ���6�?�_�17516 _�q�����&�9�tpdisc 0ɯۡݯ�������7�tpconn 0 H�Z�l�~��!�4�9?�Q�G� ۡ���Ϝ�/�0��Z� Ҫpς��%߸�ȟZ��֦��ߗߩ� }5���P�b�u߇��*�}}<�?test_�1�er�<16279�1424:263469 �ߍ��2� D���̿z������� ���������.�@��� d�v����������� ������������a w�-�?��c�� ����P]��� /(/;��q/�/ �/9�K/]/o/�/?$?|��߽27168޾ �/?�?�?��RS9 y?
OO/A�?T8�?�O�O�O8�6�?�8e�mpY7680 �vO�O_�O.�F*.d�O�N�O _�_�_�/1 J_\_n_�_o#o 6?ȯ�R�_�_o�o�o �?�?TO�Hzo0O BO�o�G�o��8���$SNPX_A�SG 2�����q� �P 0 '%�R[1]@1.Y1��y?��s%� !��E�(�:�{�^��� ����Տ��ʏ��� A�$�e�H�Z���~��� џ����؟�+��5� a�D���h�z�����ů �ԯ���
�K�.�U� ��d�������ۿ��� ���5��*�k�N�u� �τ��ϨϺ������ 1��U�8�Jߋ�nߕ� �ߤ����������%� Q�4�u�X�j���� ���������;��E� q�T���x��������� ��%[>e �t������ !E(:{^� �����/�/ A/$/e/H/Z/�/~/�/ �/�/�/�/�/+??5? a?D?�?h?z?�?�?�? �?�?O�?
OKO.OUO �OdO�O�O�O�O�O�O _�O5__*_k_N_u_ �_�_�_�_�_�_�_o 1ooUo8oJo�ono�o��o�d�tPARAM� �u�q ��	��jP�d�9p�ht��pO�FT_KB_CF�G  �c�u�sO�PIN_SIM  �{vn���p�pRVQSTP/_DSBW~r"t|�HtSR Zy� � &!pOB�195_SERV� M���vTO�P_ON_ERR�  uCy8�PT�N Zuk��A4�RING�_PR�D��`V�CNT_GP 2�Zuq�!px 	 r��ɍ���׏��w�VD��RP 1�i p�y��K�]� o���������ɟ۟� ���#�5�G�Y���}� ������ůׯ���� �F�C�U�g�y����� ����ӿ��	��-� ?�Q�c�uχϙϫ��� ��������)�;�M� _�qߘߕߧ߹����� ����%�7�^�[�m� ������������ $�!�3�E�W�i�{��� ������������ /ASew��� ����+= Ovs����� ��//</9/K/]/ o/�/�/�/�/�/�/? �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O�O)�PRG_CO7UNT8v�k�GuNKBENB��FEMpC�:t}O_UPD 1}�{T  
4O r�O�O�O__!_3_ \_W_i_{_�_�_�_�_ �_�_�_o4o/oAoSo |owo�o�o�o�o�o�o +TOas �������� ,�'�9�K�t�o����� ����ɏۏ����#� L�G�Y�k��������� ܟן���$��1�C� l�g�y���������ӯ ����	��D�?�Q�c� ��������ԿϿ�� ��)�;�d�_�q�=L�_INFO 1޵E�@ �2@���������� ��ٽ`y*�d��h'��¬߾�=`y;MYS�DEBUGU@�@���d�If�SP_PwASSUEB?xۿLOG  ��ʠC��*ؑ�  ���A��UD1�:\�ԘΥ�_MPAC�ݵE&�8�A���V� �A�SAV �!�������X����SVZ�TEM�_TIME 1"����@ 0  fX���������$T1SVGU�NS�@VE'�E���ASK_OPT�IONU@�E�A�A�+�_DI��qOG�B�C2_GRP 2�#�I�����@� � C���<Ko�CF�G %z��� 8�����`��	� .>dO�s� ������* N9r]���� ���/�8/#/\/n/v$Y,�/Z/�/�/ H/�/?�/'??K?]� k?=�@0s?�?�?�?�? �?�?O�?OO)O_O MO�OqO�O�O�O�O�O _�O%__I_7_m_[_ }__�_�_�X� �_�_ oo/o�_SoAoco�o wo�o�o�o�o�o�o =+MOa�� �������9� '�]�K���o������� ��ɏ���#��_;�M� k�}��������ß� ן��1���U�C�y� g�������������� �	�?�-�c�Q�s��� �������Ͽ��� �)�_�Mσ�9��ϭ� ������m���#�I� 7�m�ߑ�_ߵߣ��� ��������!�W�E� {�i���������� ����A�/�e�S�u� w������������� +=O��sa�� �����9 ']Kmo��� ����#//3/Y/ G/}/k/�/�/�/�/�/ �/�/??C?��[?m? �?�?�?-?�?�?�?	O �?-O?OQOOuOcO�O �O�O�O�O�O�O__ ;_)___M_�_q_�_�_ �_�_�_o�_%oo5o 7oIoomo�oY?�o�o �o�o�o3!Ci W������ ���-�/�A�w�e� ���������я�� �=�+�a�O���s��� ����ߟ͟��o�-� K�]�o�ퟓ�����ɯ��צ��$TB�CSG_GRP �2&ץ��  �� 
 ?�  6�H�2� l�V���z���ƿ��������(�d׊E+�?�	 �HC���>���G����C�  �A�.�e�q�C��N>ǳ33��S�/]���Y��=Ȑ� C\�  Bȹ��B���>����P���KB�Y�z��L�H�0�$����J�\�n�����@�Ҿ����� ����=�Z�%�7��鈴�?3�����	�V3.00.�	�cr35��	*����
�������Ƈ� 3��4�  7 {�CT�v�,}��J2�)��������CFG +�ץ'� *�������I����.<
�<b M�q����� ��(L7p[ ������/ �6/!/Z/E/W/�/{/ �/�/�/�/.�H��/? ?�/L?7?\?�?m?�? �?�?�?�? OO$O�? HO3OlOWO|O�O��� �Oӯ�O�O�O!__E_ 3_i_W_�_{_�_�_�_ �_�_o�_/oo?oAo So�owo�o�o�o�o�o �o+O=s� E���Y���� �9�'�]�K�m����� ��u�Ǐɏۏ���5� G�Y�k�%���}����� ßşן���1��U� C�y�g�������ӯ�� ����	�+�-�?�u� c����������Ͽ� ��/�A�S�����q� �ϕϧ��������%� 7�I�[���mߣߑ� �������߷��3�!� W�E�{�i����� ��������A�/�e� S�u������������� ��+aO� s��e����� 'K9o]� ������#// G/5/k/}/�/�/[/�/ �/�/�/�/??C?1? g?U?�?y?�?�?�?�? �?	O�?-OOQO?OaO �OuO�O�O�O�O�O�O ___M_�e_w_�_ 3_�_�_�_�_�_oo 7o%o[omoo�oOo�o �o�o�o�o!3�o �oiW�{��� ����/��S�A� w�e�������я���� ���=�+�M�s�a� ��������ߟ�_	� ��_ן]�K���o��� ����ۯɯ���#�� �Y�G�}�k�����ſ ׿��������U� C�y�gϝϋ��ϯ��� �����	�?�-�c�Q� s�u߇߽߫������ ��)��9�_�M���� /����i������%� �I�7�m�[������� ������������E Wi{5���� ����A/e S�w����� /�+//O/=/_/a/ s/�/�/�/�/�/�/? '?��??Q?c??�?�? �?�?�?�?�?O�?5O GOYOkO)O�O}O�O�O��O�N  �@S� V_R�$T�BJOP_GRP� 2,�E�  ?�Vi	-R4S.;\��@�|u0{SPU �>��UT� @�@LR	 ��C� �Vf  �C���ULQLQ>�33�U�R�����U�Y?�@=�Z�C��P��ͥR�>�P  B��W$o�/gC��@g�d�Db�^����eeao�P&ff�e=��7LC/kaB� o�o�P��P�ef�b-C�p��^�g`�d�o�PL�Pt<�eVC\  �Q�@�'p�`�  �A�oL`�_wC�BrD�S�^��]�_�S�`<P�B��P�anaa`C�;�`L�w�aQo�xp�x�p:���XB$'tMP@�PCAHS��n���=�P𥅡�trd<M�g E�2pb����X�	� �1��)�W���c�� ����������󟭟�7�Q�;�I�w���;d��Vɡ�U	V3�.00RScr35QT*�QT�A��� E�'�E�i�FV#�F"wqF>���FZ� Fv�R�F�~MF����F���F��=�F���F�ъ�F��3F����F�{G
�GdG��G#
�D���E'
EMK�E���E����E�ۘE����E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F���vF�u�<#�_
<t���ٵ�=�_��V� �R�p�V9� ]E_STPARtp�H�FP*SHR\�ABL/E 1/;[%�S�G�� �W�G�BG�G� WQG�	G�E
G�GȖ�QG��G�G�ܱv�RD	I~�EQ�ϧϹ�������W�O_�q�{ߍߐ�߱���w�S]�CS  !ڄ���������� ��&�8�J�\�n��� ���������� ]\�`� ��	��(�:������
��.�@�w�NUoM  �EEQ�P	P ۰ܰw�_CFG 0���)r-PIMEBF_TTb��CSo�,GVERڳ-B,�R 11;[ 8I��R�@� �@&  ����� ��//)/;/M/_/ q/�/�/�/�/�/?�/ ?J?%?7?M?[?m?> �@�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_l�_�Y@cY�M�I_CHAN8 �c cDBGLVĂ�:cX�	`ET�HERAD ?*f�\`��?�_�uo�oQ�	`ROUT6V!	
!�d�o~�lSNMASKQh|cba255.u�ߣ'9ߣY�OOLOFS_DIb���U;iORQCT�RL 2		�Ϸ~T����� #�5�G�Y�k�}����� ��ŏ׏�����.���R�V�PE_DE�TAI/h|zPGL�_CONFIG �8�	���/�cell/$CID$/grp1V�@̟ޟ����Ӏ�o ?�Q�c�u�����(��� ϯ������;�M� _�q�����$�6�˿ݿ ���%ϴ�I�[�m� ϑϣ�2��������� �!߰���W�i�{ߍ��߱�%}F�������/�A�C�i�H� Eߞ����������?� �.�@�R�d�v���� ������������* <N`r��� ����&8J \n��!��� ��/�4/F/X/j/ |/�//�/�/�/�/�/ ??�/B?T?f?x?�? �?+?�?�?�?�?OO �?>OPObOtO�O�O�O����User� View ��}�}1234567890�O�O�O_#_`5_=T�P��]_���I2�I:O�_�_�_�_�_�_X_j_�B3�_GoYo�ko}o�o�o o�op^4 6o�o1CU�ovp^5�o���� �	�h*�p^6�c� u����������ޏp^7R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3� �OM�_�q��������y  e��Yz���	�� -�?�Q���uχϙ�俀����������>�� e�5i��c�u߇ߙ߫� ��d������P�)�;� M�_�q��*�<��i� ��������)���M� _�q������������ ����<�û��=Oa s��>����* '9K]f� Q�������/ �%/7/I/�m//�/ �/�/�/n<��^/? %?7?I?[?m?/�?�? �? ?�?�?�?O!O3O �/<׹��?O�O�O�O �O�O�?�O_!_lOE_�W_i_{_�_�_FOXG9 +_�_�_oo(o:o�O Kopo�o)_�o�o�o�oP�o ��	g�0�o M_q���No� ���o�%�7�I�[� m�&l�n��Ə؏ ���� ��D�V�h� ��������ԟ柍� g�ڻ}�2�D�V�h�z� ��3���¯ԯ���
� �.�@�R���3uF�� ����¿Կ������ .�@ϋ�d�vψϚϬ� ��e�w���U�
��.� @�R�d�ψߚ߬��� ��������*���w� ��v������� w�����c�<�N�`� r�����=�w��-��� ��*<��`r ����������  ��1C Ugy�����<��    -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_��  
��(  }�%( 	 y_ �_�_�_�_�_�_o	o +o-o?ouoco�o�o�o:�Z* �Q &�J\n�� ����o���9� (�:�L�^�p������ ���܏� ��$�6� }�Z�l�~�ŏ����Ɵ ؟���C�U�2�D�V� ��z�������¯ԯ� ��
��c�@�R�d�v� ����᯾�п�)�� �*�<�N�`ϧ����� �Ϻ��������&� 8��\�n߀��Ϥ߶� ��������E�"�4�F� ��j�|������� �����e�B�T�f� x�������������+� ,>Pb��� ������� (o�^p��� ���� /G$/6/ H/�l/~/�/�/�/�/ /�/�/?U/2?D?V?�h?z?�?�/�`@  �2�?�?�?�3�7�P���!frh:\�tpgl\rob�ots\m20i�a\cr35ia.xml�?;OMO_O qO�O�O�O�O�O�O�O ���O_(_:_L_ ^_p_�_�_�_�_�_�_ �O�_o$o6oHoZolo ~o�o�o�o�o�o�_�o  2DVhz� �����o�
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ �ݟ��&�8�J�\� n���������ȯߟٯ ���"�4�F�X�j�|�@������Ŀ־�8.1� �?@88�?�ֻ�ֿ� 3�5�G�iϓ�}ϟ��� ���������5��A��k�U�wߡ߿��$T�PGL_OUTP�UT ;�!�!/ ������ ��,�>�P�b�t�� ������������ (�:�L�^�p�������������2345678901������ ���"��BT fx��4�����
}$L^ p��,>���  //$/�2/Z/l/~/ �/�/:/�/�/�/�/?  ?�/�/V?h?z?�?�? �?H?�?�?�?
OO.O �?<OdOvO�O�O�ODO VO�O�O__*_<_�O J_r_�_�_�_�_R_�_ �_oo&o8o�_�_no �o�o�o�o�o`o�o�o "4F�oT|� ���\��}���@��0�B�T�e�@�������� ( 	 ��Џ����� �<�*�L�N�`����� ����ޟ̟���8� &�\�J���n�������@��ȯ���"������ �*�X�j�F�����|� ¿Կ��C���ϱ�3� E�#�i�{�忇ϱ�S� ���������/ߙ�S� e�߉ߛ�y߿���;� ������=�O�-�s� ���ߩ��]������� �'����]�o���� ��������E����� 5G%W}����� �g���1� Ug	w�{�� =O	//�?/Q/// u/�/��/�/_/�/�/ �/�/)?;?�/_?q?? �?�?�?�?�?G?�?O �?OIO[O9OO�O�? �O�OiO�O�O�O!_3_ �O_i_{__�_�_�_��_�_�R�$TPOFF_LIM >�|op:��mq�bN_SV`  �l�jP_MOoN <6�d�opop2l�aST�RTCHK =�6�f� bVTCOMPAT-h�af�VWVAR >rMm�h1d �o� �oop`ba_�DEFPROG �%|j%ROB�195_SERV�	�j_DISPL�AY`|n"rINST_MSK  t|w ^zINUGp��odtLCK�|}{QUICKMEN��dtSCRE�p�6��btpsc@dt�q��b*�_.��ST�jiRACE_CFG ?Mi��d`	�d
?��u�HNL 2@"|i����k r͏ ߏ���'�9�K�]��w�ITEM 2A��� �%$12�34567890<����  =<��П<��  !���p��=��c��^� ���������.���R� �v�"�H�ί��Я� �����*�ֿ���r� 2ϖ�����4�޿�ϰ� ��&���J�\�n���@� ��d�v��ς������ 4���X��*��@�� ���ߨ������� T���x������l� �������,�>�P��� ����FX��d���� ��:�p" ��o����� F6HZt~�� N/t/�/��// /2/ �/V/?(?:?�/F?�/ �/�/j?�??�?�?R? �?v?�?QO�?lO�?�O �OO�O*O|O_`O _ �O0_V_h_�Ot_�O_ _�_8_�_
oo�_@o �_�_�_Lodo�_�o�o 4o�oXojo3�oN�o r��o��s��S�B���z� 3 h��z ��C�:y
 P�v�]���~�UD1:\������qR_GRP� 1C��� 	 @Cp���@$��H�6�l�Z��|� ����f���˟���ڕ?�  
���<� *�`�N���r������� ޯ̯��&��J�8�Z���	�u�����s�SCB 2D� �����(�:��L�^�pς��|V_C�ONFIG E����@����ϖ�OUTPUT F�������6�H� Z�l�~ߐߢߴ����� �������#�6�H�Z� l�~���������� ����2�D�V�h�z� ��������������
 �.@Rdv�� �����) <N`r���� ���//%8/J/ \/n/�/�/�/�/�/�/ �/�/?!/4?F?X?j? |?�?�?�?�?�?�?�? OO/?BOTOfOxO�O �O�O�O�O�O�O__ +O>_P_b_t_�_�_�_ �_�_�_�_oo'_:o Lo^opo�o�o�o�o�o �o�o $����!� bt������ ���(�:�-o^�p� ��������ʏ܏� � �$�6�G�Z�l�~��� ����Ɵ؟���� � 2�D�U�h�z������� ¯ԯ���
��.�@� Q�d�v���������п �����*�<�M�`� rτϖϨϺ������� ��&�8�J�[�n߀� �ߤ߶���������� "�4�F�W�j�|��� ������������0� B�S�f�x��������� ������,>P a�t��������(:L/x���k}gV �K���//&/ 8/J/\/n/�/�/�/W �/�/�/�/?"?4?F? X?j?|?�?�?�?�/�? �?�?OO0OBOTOfO xO�O�O�O�?�O�O�O __,_>_P_b_t_�_ �_�_�O�_�_�_oo (o:oLo^opo�o�o�o �o�_�o�o $6 HZl~����o ���� �2�D�V� h�z��������ԏ� ��
��.�@�R�d�v� ��������Ϗ���� �*�<�N�`�r����� ����˟ޯ���&� 8�J�\�n����������Ż�$TX_SCREEN 1G�g�}�ipnl/��g?en.htmſ��*�<�N�`ϽP�anel setupd�}�dϥϷ����������ω�6� H�Z�l�~ߐ�ߴ�+� ������� �2�߻� h�z������9�g� ]�
��.�@�R�d��� ������������� }���<N`r�� ;1��& 8�\��������QȾUALR�M_MSG ?��� �Ȫ-/ ?/p/c/�/�/�/�/�/ �/�/??6?)?Z?%�SEV  -��6"ECFG �I��  }ȥ@�  A�1�   B�Ȥ
 [?ϣ��?OO%O 7OIO[OmOO�O�O�G~�1GRP 2J�;w 0Ȧ	 �?��O I_BBL_NOTE K�:�T��l�Ϣ�ѡ�0RDE�FPRO %+ (%N?u_Ѡc_�_ �_�_�_�_�_o�_o�>o)oboMo�o\INUSER  R]��O�oI_MENH�IST 1L�9 � ( _P���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1�oCUgy�)
13/������p� �}936�I�[�m��� ������̏ޏ����� &�8�J�\�n������ ��ȟڟ�����"�4� F�X�j�|������į ֯�����f9Rq�� B�T�f�x��������� ҿ����ϩ�>�P� b�tφϘ�'�9����� ����(߷�L�^�p� �ߔߦ�5������� � �$����Z�l�~�� ���C�������� � 2��/�h�z������� ��������
.@ ��dv����� _�*<N� r�����[� //&/8/J/\/��/ �/�/�/�/�/i/�/? "?4?F?X?C�U��?�? �?�?�?�?�/OO0O BOTOfO�?�O�O�O�O �O�O�O�O_,_>_P_ b_t__�_�_�_�_�_ �_�_o(o:oLo^opo �oo�o�o�o�o�o  �o$6HZl~i? {?������ 2�D�V�h�z����-� ԏ���
����@� R�d�v�����)���П ���������N�`� r�������7�̯ޯ� ��&���J�\�n�����������$UI�_PANEDAT�A 1N����ڱ  	�}�����!�3�E�W� )Y�}�7�� �Ϻ��������i�&� �J�\�C߀�gߤߋ� ����������"�4��\X�7�� �q}� �ϕ���������B� ���%�I�[�m���� ��
�����������! E,i{b�� ����l�ܳ 7�<N`r��� �-���//&/8/ �\/n/U/�/y/�/�/ �/�/�/?�/4?F?-? j?Q?�?�?%�?�? �?OO0O�?TO�xO �O�O�O�O�O�OKO_ �O,__P_b_I_�_m_ �_�_�_�_�_oo�_ :o�?�?po�o�o�o�o �oo�o sO$6H Zl~�o���� ��� �2��V�=� z���s�����ԏGoYo �.�@�R�d�v�ɏ ����П����� �<�N�5�r�Y����� ��̯���ׯ�&�� J�1�n�������ȿ ڿ����c�4ϧ�X� j�|ώϠϲ���+��� �����0�B�)�f�M� �ߜ߃��ߧ������� ��P�b�t��� ��������S���(� :�L�^����i����� ������ ��6 ZlS�w�'�9�}���"4FX)�}��l�� ���/j'//K/ 2/D/�/h/�/�/�/�/ �/�/�/#?5??Y?���C�=��$UI_P�OSTYPE  �C�� �	 e?�?�2QU�ICKMEN  ��;�?�?�0RE�STORE 1O�C�  '�L?��6OCC1O��maO�O�O�O�O �OuO�O__,_>_�O b_t_�_�_�_UO�_�_ �_M_o(o:oLo^oo �o�o�o�o�o�oo  $6H�_Ugy �o������ � 2�D�V�h�������� ԏ����w�)� R�d�v�����=���П ������*�<�N�`� r��������ޯ� ��&�ɯJ�\�n��� ����G�ȿڿ������7SCRE�0?��=u1sc�+@u2K�3K�4�K�5K�6K�7K�8<K��2USER-�2ϦD�ksMì�3��4���5��6��7��8����0NDO_CFG P�;� ��0PDATE ����None��2��_INFO �1QC�@��10% �[���Iߊ�m߮��� �����������>�P�3�t��i���<-�O�FFSET T�=�ﲳ$@����� �1�^�U�g������� ���������$-�ZQcu���?�
�����UFRAM/E  ����*��RTOL_ABRqT	(�!ENB*~GRP 1UI��1Cz  A� �~��~����B����0UJ��9MSK  hM@�;N%8��%��/�2VCCMf��V�ͣ#RG�#EY�9���/����-D�BH�p71�C���3711?�lC0�$MRf2_�*PS�Ҵ�	����~XC56 *ȋ?�6���1$�5ڴ��A@3C�N�. ��8�? ��OOKOx1FOsO�5�51��_O�O�� B����A 2�DWO�O7O_�O8_ #_\_G_�_k_}_�__ �_�_�_�_"o�OFoXo.�%TCC�#`mI1��i������ G�FS��2aZ; ��| 2345678901�o�b��� ��o��!5a�4�BwB�`56 311:�o=L�Br5v1 �1~1�2��}/��o�a ��#�GYk} �p�������ُ �1�C�U�6�H���5� ~���ߏ���	���4>�dSELEC)M!�v1b3�VIRToSYNC�� ����%�SIONTM�OU�������F��#b������(u F�R:\H�\�A\��� �� M�C��LOG��  � UD1��EX�����' B@ ����̡m���̡  OBCL�1��H� �  �=	 1- n6  -�������[�,S�A�`=�S�͗��ˢ��TRAIN⯞b�a1l�
0d�$j�T2cZ; (aE2� ��i��;�)�_�M�g� qσϕϧ���������	��F�STAT dm~2@�zߌ��*j$i߾��_GE��#eZ;�`0��
� 02��HOM�IN� f����� ~�����Б�C�g�X���JMP�ERR 2gZ;
  ��*jl�V�7� �������������
���2�@�q�d�v�B�_�ߠRE� hWޠ$L�EX��iZ;�a1-�e��VMPHASOE  5��c&���!OFF/�F�PU2n�j�0��
��E1@��0ϒE1!1?s33�����ak/�kxk䜣!
W�m[�䦲�[�����o3;�  [i{�� ��/�O�?/ M/_/q/��/��// �/'/9/�/=?7?I?s? �/�?�/�/�?�??O m?O%O3OEO�?�?�O �?�O�O�?�O�O�O_ _gO\_�OE_�O�_�O �O/_�_�_�_oQ_Fo u_�_|o�o�_�oo�o �o�o�o;oMo?qof -�oI���� �7�[P��� ������ˏ��!�3� (�:�i�[�ŏg�}�������TD_FIL�TEW�n�� �ֲ:���@���+� =�O�a�s�������� �֯�����0�B��T�f�x���SHIF�TMENU 1o[�<��%��ֿ�� ��ڿ����I� �2� �V�hώ��Ϟϰ��������3�
�	LIVE/SNAP'�vsfliv���E����ION� * Ub�h�menu~߃�����ߣ�6��p���	����LE�.�50�s�P��@� ��AɠB8
z�z��}��x�9�~�P�� ����MEb���<�Z0���MO��q����z�WAITD_INEND�������OK1�OU�T���SD��TI]M����o�G� ��#���C���b�������RELEASE�������TM����=���_ACT[������_DATA r��%L�����xRDISb�E_�$XVR�s����$ZABC_G_RP 1t�Q��,#�0�2���ZIP�u'�&�����[MPCF_OG 1v�Q�0��/� w�ɤ�� 	�Z/  85�/�/H/�/l$?��+�/�/�/?�/��/???r?�?  �D0�?�?�?�?�?�;���x�]h_YLIND֑y�� ��� ,(  *VOgM.�SO�OwO�O�M i?�O�O ^PO1_�OU_<_N_�_ �O�_�_�__�_�_x_ -ooQo8o�_�o�oY�&#2z� � ��oC�e?a?>N|h�oq����qA�$D�SPHERE 2{6M��_�;o�� �!�io|W�i��_�� ,��Ï���Ώ@�� /�v���e�؏��p�����������ZZ�� �N