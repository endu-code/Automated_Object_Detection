��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CESS0s!_81s!J3�> �! � �$SOFT�T_�IDk2TOTAL7_EQs $�0�0�NO�2U SPI_OINDE]�5Xk2SCREEN_(4�_2SIGE0�_?q;�0PK_FI�� 	$THK�YGPANE�4 �� DUMMY1"dDDd!OE4LA!�R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Dc@�D5�F6�F7*�F8�F9�G0�G�G@JA�E�GbA�E�G1�G!1�G �F�G2�B!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HO30IO�0� }%�SMACRO�ROREPR�X� D+��0��R{�T UT�OBACKU��0 �)DE7VIC�CTI*0�A� �0�#�`B�S�$INTERVA�LO#ISP_UN9I�O`_DO>f7�uiFR_F�0AI�N�1���1c�C�_WAkda�jOF�F_O0N�DEL��hL� ?aA�a1bc?9a�`C?��P��1E��#sATB��d��MO� �cE' D [M�c���^qREV�BI�Lrw!XI� QrR�  � OD��P�q$NO�^PM�Wp�t�r/ "�w� �u�q�r�0�D`S p �E RD_E�pCq�$FSSBn&$CHKBD_SE^e�AG G�"$SLOT_��2=�� 	V�d�%��3 a�_EDIm  O � �"��PyS�`(4%$EP�1��1$OP�0�2��a�p_OK�UST1P_C� ��d���U �PLACI4!��Q�4�( raCOM9M� ,0$D�����0�`��EOWBn�IG�ALLOW� �(K�"(2�0VAARa��@�2ao�L�0;OUy� ,Kva�y��PS�`�0M_O�]����CCFOS_UT~p0 "@�1�3�#�ؗ`X"��}R0  4F IMCM�`O#S�`��Hupi �_�p�BA�!���M/ �h�pIMPEE_F�N��N���@O���r�D_�~�n�Dry�F� dCC_��r0  T� '��'�DI�n0"��pu�P�$I�������F�t XF� GRP0��M=q�NFLI�7��0U�IRE��$g"� S�WITCH5�AX�_N�PSs"CF_�LIM� �; �0EED��!���qP�t�`PJ_dVЦMODEh�.Z`��PӺ�ELBOF � ������p� ���3���� FB/���0�>�G� �>� WARNM�`/���qP��n�NST�� COR-0bF�LTRh�TRAT�PT1�� $AC�C1a��N ��r$�ORI�o"V�RT��P_S� CHG*�0I��rT2��1
�I��T�I1��>� x i#�Q\��HDRBJ; TCQ�2L�3L�4L�U5L�6L�7L�8L��9s!��O`S <F +�=�O��#92^��LLECy�"MULTI�b�"N���1�!���0T�� �STY�"�R`�=l�)2`����*�`T  |� �&$��۱m��P�̱�UT�O���E��EXT�����ÁB���"2Q� (䈴![0�������<�b+�� "D"���ŽQ��<煰kc!(�9�#���1���ÂM�ԽP��" q'�3�$ L� �E���P<��`A�$�JOBn�T���l�TwRIG3�% dK� ������<���\��+��Y�p�_M��&� t�pFLܐBN9G AgTBA� �� �M��
�!��p� �q��0�P[`��O�'[���0tna*4���"J��_R���ECDJ��IdJk�D�%C�`�Z���0���P_�P��@ ( @F RO.��&�t�sIT�c�NOMࠀ
����S� �`T)"w@���Z�P�d���RA�0��2b"�����
$T����MD%3�T��`U31��ʩp(5!HGb�T1�*E�7�c�KAb�pWAb�cA4#YNT��>�PDBGD�� *(��PUt@X���W���AX��a��ewTAI^cBUF���0!+ � l7n�PIW�*5 P�7M�8M�9
0�6}F�7SIMQS@�>KEE�3PAT�n�^�a" 2`#�"�L�64FIX!, !���!d��D�2Bus�=CCI�:FPCH�P:BAD�aHCEhAOGhA]HW�_�0>�0_h@�f�Ak���F�q@\'M`#�"�DE3�- l�p3G��@FSOES]FgHBSU�I�BS9WC��. ` =��MARG쀳β�FACLp�SLEWxQe�ӿ�6�MC�/�\pSM_JBM����Q�YC	g�e#�0� ā�CHN-�MP�$G� Jg��_� #��1_FP$�!TCuf!õ#�� ���d�#a��V&��r��a;�fJR���rSoEGFR�PIO�^ STRT��N���cPV5���!41 �r��
r>İ�b�B�~O�2` +� [���,qE`&�,q`y��Ԣ}t��yaSIZ%���t�vT�s� �z|�y,qRSINF} Oбc���k��`��`��`L�ĸ T`7�CRCf�ԣCC/�9��`�a�uah�ub'�MIN@��uaDs�#�G�D�YC��C�����e�q0���� �EV�q�F*�_�eF��N3�s�Pah��Xa+p,5!��#1�!VSCA$?� A��s1�"!3 ��`F/k��_�U ��g��]��C�� a�s���R�4� �����N����5a�R��HANC��$L�G��P�f1$+@NYDP�t�AR5@N^�`�a�q���c��ME�108���}0��RAө�CAZ 𨵰�%O��FCTK��s`"��S�PFADIJ�O J�ʠ�ʠ���<����Ր��GI�p�B�MP�d�p�Dba��AcES�@	�K�W_���BAS�� �G�5 � M�I�T�C�SX[@@�!62�	-$X���T9�{s�C��N�`�a~P_H�EIGHs1;�WI�D�0�aVT ACϰ�1A�Pl�<����EXPg���|��C}U�0MMENU���7�TIT,AE�%)�a2��a��g8 P� a�ED�E� ��PDT��R�EM.��AUTH?_KEY  ����R�� �b�O	���}1ERRLH� �9c \� �q-�OR�D�B�_ID�@l �PU�N_O��Y�$SCYS0��4g�-�I��E�EV�#q'�P�XWO�� �: �$SK7!f2 &�T�d�TRL��; ��'AC�`��ĠINMD9DJ.D��_��bf1��f���PL�A��RWAj���SD��A��!+r|��U�MMY9d�F�10�d�&���J�<��}1P�R� 
3�PO9S��J�= ��$V$�q�PLB~�>���SܠK�?�����CJ�@����EN5E�@T��A���S�_�RECOR��B�H 5 O�@7=$LA�>$~�r2��R��`�q�b`�_DLu��0RO�@�aT[� Q��b������! }О��PAUS���dE�TURN��MR�U�  CRp�E�WM�b�AGNAL:s2$LA�!�?$PX�@$P�y A �Ax�1C0 #ܠDO�`X��k�W�v�q�GO_A7WAY��MO�ae����]�CSS_C�CSCB C �8'N��CERI����J`u�QA0�}���@�GAG� R �0�`��{`��{`OF�q�5��#+MA��X��І�LL�D� �$���sU�D)E%!`|���OVR10W��,�OR|�'�$E�SC_$`�eDSB#IOQ��l ��B.�VIB&� �c,������f�=pSSW����f!VL��PL|���ARMLO
���`����d7%SC� �bALspH�MPCh �Ch �#h �#
h 5�UU���C�'��C�'�#�$'�d�#C \4�$�pH��Ou��!Y��!�SB���` k$4�C�P3Wұ46�$VOLT37$$`�*�^1���$`O1*�$o��0R�QY��2b4�0DH_THE����0S�<�4�7ALPH�4�`����7�@ �0�qb7
�rR�5�88� ×@���"��Fn�	MӁVHBPFUAF�LQ"D�s�`�THR��i2dB�����G
(��PVP�����������1�J2�B�E�C�E�CPSu�Y@��F b3���H�(V�H:U�G��
X0��FkQw�[�N�a�'B���C INH=BcFILT��� $��W�2�T1�[ @��$���H YАAF�sDO��Y�R p� fg�Q�+�c5h`�Q�iSh�QPL��x�Wqi�QTMOU�# c�i�Q\��X�gmb��Hvi�h�bAi�fI�aCHIG��ca	xO��hܰ��W�"vAN-uX!��	#AV�H!Pa8$P�ד#p�RE_:�A�a��B�qN0�X�MCN�0��f1[1�qVE�p��Z2;&f�I�QO�u�r�x�wGldDN{G|d��aF>!�9��a9M:�U�FWA�:�Ml���X�Lu��$!����!l�ZO����0%�O�lF�s�13�DI�W�@��Q����_��!CURVAL԰0rCR41ͰZ�C <�r�H�v���<�`��<�(�f�CH�QR3��S���t���Xp�VS!_�`�ד�F��ژ������N�STCY_ E L����1�t�1�T�U��24�2B�NI �O7������DEV�I|� F��$�5�RBTxSPI2B�P���BYX�����T��HNDG>��G H tn���L��Q�C���t5��Lo0 H���閻�FBP�{tF�E{�5�t��T��I��DO���uPMC�S�v>�f>�t�"HOOTSW�`s�?wELE��J T��@�e�2��25�� O� ��HA7�E��344�0q?��A�K �� �MDL� 2J~PE��	A��s��t��È�s�JÆG!��r�D"�ó�����\�TO���W�	��/��SL{AV�L  �0INPڐ���`%ن�_CFd�M� $��ENU��O�G��b�ϑ]զP�0�`ҕ�]�IDMA0�Sa��\�WR�#���"]�VE�$a�SK�I�STs��sk$��2u���J�������	��Q���_SVh�E�XCLUMqJ2M!ONL��D�Y��|�P�E ղI_V�A�PPLYZP��HI�D-@Y�r�_M�2��VRFY�0��r�<1�cIOC_f��"� 1������O��u��LS���R$DU/MMY3�!���S=� L_TP/Bv��"���AӞ�ّ Ns ���RT_u^�� �G&r�[�O D��P_B�A�`�3x�!IF ��_5���H������� �� P� $4 KwARGI���� q�2O ��_SGNZ�Q q�~P/�/PIGNs�l�$�^ sQ>ANNUN�@�T`<�U/�ߴ�LAzp�]	Z�d~�E�FwPI�@ R �@�F?IT�	$TOTA%��d����!�M�NIY�S+���E�yA[�
DAYS\ԃADx�@��	� ��EFF_AXIb?�TI��0zCOJ�A �ADJ_RWTRQ��Up��H<P�1D �r5̀Ll�T�0? ]P�"p���mtpd��V 0@w�G���������SK�SU� ��C�TRL_CA�� �W�TRANS��6PIDLE_PAW���!��A�V���V_�l�V ��DIAGS���X� /$2�_SE�#TAC���t!�!00z*@��RR��vP�A���p ; SW��!�!�  ��ol�U���oOH��PP̱ ��IR�r��BR1K'#��"A_Ak��� x 2x�9ϐZs2���%l�W�0t*�x%R7QDW�%MSx�t5�AX�'�"��LIF�ECAL���10��N�1{"�5Z�3{"�dp5�ZU`}�MOT�N°Y$@FLA��cZOVC@p�5H�E	��SUPPOQ�ݑAq� Lj (C��1_X6�IEYRJZRJWRJ�0TH�!UC��>6�XZ_AR�p�Y2�HCOQ��S�f6AN��w$�I{CTE�Y `��CACHE�C9øM�PLAN��U7FFIQ@�Ф0P<�1	��6
�	�wMSW�EZ 8w �KEYIM�p��TM~�SwQq�wQ#�|���OCVIE� ��[ A�BGL8��/�}�?� TR?�j�D\p�ذST��!�R� �T� �T� x�T	��PEMAIf��ҁ��_FAU%L�]�Rц�1�qU�� �TRE�^< $Rc��uS�% IT��BCUFW}�W��N_�N� SUB~d��C|�p�Sb�q�bSAV�e �bu �B��� �gX�^AP�d�u+p�$�_~`8�e�p%yOTT���
�sP��M��OtT�Lw#AX � ��X~`9#��c_G�3
�YN)_1�_�D��1� �2M���T��F��H@ g�`� 0p��Gbn-sC_R�AIK���r�t�RoQ�u7hN�qDSPq��rP��A�IM�c6�\����sB2�U�@�A�sM*`#IP���s�!DҐ6�CTH�@n�)�OT�!�6�HSDI3�AB#SC���@ Vy���� �_D�CONVI�G���@3�~`F�!�pd��psq�SCZ"���sMERk��qFB��k��p�ET���aeRFU&:@DUr`����x�CD,���@p;cHR�A!��bp�Ք�Ք+PSԕC��r�C��p��Е|Sp�cH *�LX�:cd�Rqa�| �� ��W��U��U��U�P	�U�OQU�7R�8R��9R��0T�^�1k�1�x�1��1��1��1���1��1ƪ2Ԫ2T^�k�2x�2��2��U2��2��2��2ƪ�3Ԫ3^�3k�x�3P���o���3��3���3ƪ4Ԣ�EX9Tk!0�d <� 7h �p�6�pO��p����Na�FDRZ$eT^`V�Gr����䂴2�REM� Fj��BO�VM��A�TR�OV�DT�`-�MX<�IN��0,�W!'INDKЗ
w�׀�p$DG~q36���P�5�!D�6�RI�V���2�BGEAR��IO�%K�¾DN �p��J�82�PB@�CZ_MCM�@�1��r@U��1�f ,⑞�a? ���P\I�!?I�E��BQ����`m���g� j_0Pfqg RI9e�j�k!UP2_ 3h � �cTD�p�〪�! a�����bB;AC�ri T�P�b��`�) OG��%p���p��IFI�!`�pm�>��	�PT�"���MR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4�@��Uk��� �T�FS#p�Tl �P���e�qP�p$GEX_���1M�2��2� 3�5��9G ���m ��Ѝ��SW�eOe6DEBcUG���%GR���pU�#BKU_�O�1'� �@PO��I5�5MSf��OOfswSM���E�b?��0�0_E �n �p��p�/TERM�o�ƐO�ORI+�p�HOZ�SM_���b�q�P�TA��r�! �U}P�Rs� -�1��2n$�' o$�SEG,*> ELT}O��$USE�pNFIAU"4�e1����#$p$UFR����0ؐO!�0����OT�'�TAƀU�#wNST�PAT��<P�"PTHJ�����E�P rF�V"ART��``%B`�abU!REyL:�aSHFT���V!�!�(_SH+@M�$���� ��@N8r�����OVRq��rSSHI%0��UN� �a�AYLO����qI�l����!�@��@ERV]��1�?:�¦'��2��%��5�%�RC<q��EASYM�q�EFV!WJi'��}�E���!I�2��U@D��q�%Ba��
5Po��0��p6OR�MY� `G	R��t2b5n� �� ��UPa�Uu �t�")���TOCO!1S�1POP ��`P�pC�������Oі�`REPR3��aOX�P�b�"ePR�%�WU.X1��e$PW�R��IMIU�2R_	S�$VIS��#(A�UD���Dv" vΥ�$H���P_AWDDR��H�G�"�Q�Q�QБR~pDp1�w H� SZ�a���e�ex�e��SE؄�r��HS��MN~vx �0��%Ŕ��OL���p�<P��-��ACROxlP_!QND_C���ג�1�T �ROUP$T��B_�VpQ�A1Q�v��c_��i���i ��hx��i���i��v�ACk�IOU��D��gfsu^d�y $|�P_D��VB�`bPRM_�b^�ATTP_אHa�z (��OBJE�r��P��$��LE�#�s`{ � ���u�AB_x�T�~�S�@�DBG�LV��KRL�YH�ITCOU�BG�Y LO a�TE�M��e�>�+P'�,PS�S|�P�JQUER�Y_FLA�b�HQW��\!a|`u@f�PU�b�PIO�� "�]�ӂ/dԁ=dԁ���L�IOLN��}ꖐ��CXa$S�LZ�$INPU�T_g�$IP#�P4��'� ��SLvpa~��!�\�W�C-�Bx�0���pF_ASv��$L ��w �DF1G�U�B0m!���0HY��ڑ��UOPs� ` ������[�ʔ[�і"�[PP�SIP�<�іI��2���IP_MEsMB��i`� X��cIP�P�b{�_N�`����R�����bSP��p$FO�CUSBG�a~�U=J�Ƃ �  � �o7JOG�'�DI�S[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A���APHIb�Qt�]�D� J7J\����� _KEYt�� �KՀLMO�Na���$XR���ɀ��WATCHa_��3���EL��b}Sy~���s� ���!V�g� �CTR�3򲓥��LG�D�� �R��I�
LG_SIZ���J�q XIƖ�I�FDT�IH� _�jV�GȴI�F�%S O���q �Ɩ���v������K�S����w�kR�N����E�@�\���'�*�U�s�5��@L>�4�DAUZ�EA�pՀ�Dp�f��GH�B#�OGB�OO��� C���PIT���� ���REC��SCRNě���D_p�aMARGf�`��:���TH�L���S�s��W�Ը��Iԭ�JGMO�MgNCH�c��FN���R�Kx�PRGv�UqF��p0��FWD��HL��STP��V`��+���Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*� a28����Gh�0CPO��������M8��Ģ��EX��TUIv�I��(�4� @�t�x�J0J�~�P���J0��N�a�#ANqA��O"�0VAIA���dCLEAR�6DCS_HI"�/cj�O�O�SI�r�S��IGN_��vpq�uᛀT�d� DEV-�LLA �°SBUW`��x0mT<$U�EM���Ł����0�A�R���x0�σ�a�@O�S1�2�3�8a�`� �ࠜh��AN%-���-�IDX�DP�2MRO��Գ!V�ST��Rq�Y{b~! �$E&C+��p.&A&���`� L��ȟ%Pݘ��T\Q�UE�`�Ua~��_ � �@�(��`�����# �M�B_PN@ R`r��<R�w�TRIN��P���BASS�a	6I�RQ6_�M�C(�� ��C�LDP�� ETRQ�LI��!D�O9=4FALʡh2�Aq3zD᱌q7��LDq5[4q5ORG�)�2�8P�R ��4/c�4=b� 01�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?0�?RIAtaMID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCESH?RΡ�BMhPa�͠��BD4�E�q`�`�F_A�J�C[��O�H� K��� \ȶ��bTf$� ��LI��q�SREQUIR�E�#MO�\�a�XD�EBU���AL� M䵔 �p���P�c�AA�AN��
Q�qa�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N�i�PST9� � �4��LOC�RI쀀�EX�fANGx��A�AODAQ䵍��@$��9�ZMF�����f��"��%8u#ЖVSUP�%��FX�@IGGo�� �rq�"��1��#B��$���p%#by���rx���vbPDAT	AK�pE;���R���M��*� t�`MD�qI��)�v� �tĀA�wH�`��tDIyAE��sANSW�P�th���uD��)�b�ԣ(@$`� PC�U_�V6�ʠ�d�PL�Or�$`�R���BD���B�p������A�RR2�E� � ��V�A/A d�$CALI�@��G�~�2��!V��<;$R�SW0^D"��ABC�hD_J�2SE�Q�@�q_Ju3M�
G�1SP�$,��@PG�n�3m�u�3p�@��JkC���2�'AO)IMk@{BCSKP^:ܔ9�wܔ	Jy�{BQܜ�����`_AZ.B��?��EL��YAOCMaP�c|A)��RTьj���1�ﰈ��@1ќ������Z��SMaG��pԕ� ER!����AINҠACk�p����b�n _�������D��/R��DIU��CD�H�@
�#a�q$�V�Fc�$x��$���`@���b���̂�E�H �$�BELP����!ACCEL���kA°�IRC_R�pG0��T!�$PS�@B2L  ����W3��ط9� ٶPAT!H��.�γ.�3���p�A_��_�e�-B�`�C���_MG��$DD��ٰ��$FW�@�p����γ�����DE��PPAB�N�ROTSPE�Eu��O0��D�EF>Q����$U�SE_��JPQPCD��JY����-A 6qYN�@A�L�̐�nL�MOU�NG���|�OL�y�INC U��a�¢ĻB��ӑ�AENCS���q�B��X���D�IN�I��0���pzC�VE�����23_U ��b�/LOWL���:�O0��0�Di�B�PҠȠ ��PRC����MOS� gTMOpp�@-GPERCH  M�OVӤ �����! 3�yD!e�]�6�<�� ʓA����LIʓdW�ɗ��:p3�.�I�TRKӥ�AY����?Q ^���m�b��`p�CQ�� MOM�B?R�0u��D���y�0Â擰DUҐZ�S_BCKLSH_C�� ��o�n��TӀ���x
c��CLALJ���A��/PKCHKtO0�Su�RTY� B�q��M�1�q_
#Nc�_UMCP�	C�΂�SCL���LMTj�_L�0X����E�� �� ����m�h���6��P	C����H� �P�Ş�CN@�"XT����C�N_��N^C�kCS	F����V6����ϡpj���nCAT�SHs�����ָ1����֙���������PAL���_P���_P0�� e���O1u�$xJaG� P{#�OG�>��TORQU(�p� a�~����Ry������"_W��^�����4t��
5z�
5I;I ;Iz�F�`�!��_8�1���VC��0�D�B�21��>	P�?�B�5JRK��<�2�6i�DBL_�SM�Q&BMD`_D9Lt�&BGRV4
D0t�
Dz��1H_���31�8JCOSEKr�EHLN�0hK�5oDt�jI���jI<1�J�LZ1�5Zc@y��1MYqA�HQB�THWMYTHET=09�NK23z�/Rln�r@CB4VCBn�CqPASfaYR<4gQt�gQ4VSBt��R?U'GTS���Cq��a���P#���Z�C$DUu ��R䂥э2�V�ӑ��Q�r�f$NE��+pIs@�|� �$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b�FP�c�j�FR�VrhVghTd��lV�jV�kV�kUV�kV�kV�kV�iHrh�f�r�m!�x�kUH�kH�kH�kH�kUH�iOclOrhO���nO�jO�kO�kO��kO�kO�kO�FF�.bTQ���E��egSPBALANCE���RLE�PH_'US�P衅F��F��FPFULC�3��3��E��1�l�UTOy_p �%T1T2t���2NW�����ǡ@��5�`�擳�T��OU���� INSE9G��R�REV��R����DIFH��1�l��F�1�;�OB��;C��2� �b�4?LCHWAR��;��ABW!��$ME�CH]Q�@k�q��AXk�P��IgU�i��� 
���!����ROB��CR��ͥ�8*�C��_s"T �� x $W�EIGHh�9�$�cc�� Ih�.�IF� ќ�LAGK�8S�K��K�BIL?�O1D��U��STŰ�P�; �����������
�Ы�L�� � 2�`�"�DEB�U.�L&�n��PM'MY9��NA#δ�9�$D&���$���� Q �D�O_�A��� <@	���~��L�BX�P�N��+�_7�L�t��OH  �� E%��T���ѼT��<���TICK/�C��T1��%������N��c�Ã�R L�S���S�����PROM�Ph�E� $IR� X�~ ���!҇MAI�0��j���_�9����t�l�Rn�0COD��FU`�+�ID_" =����~�G_SUFF<0G 3�O����DO��ِ��R��Ǔـ��S����!{�������	�H)�_FI���9��ORDX� ����36��X������GR9�S��Z�DTD��v�ŧ�4 *�L_N�A4���K��DEF_I[�K���g��_����i��Ɠ�š���IS`i �萚����e����4�0i��Dg����D� O|��LOCKEA!�uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ�{� ���}��v�Ա�� g������^���K‒Փ����!w�N�P@'���^���,`�W\�l[R�7�TEF�Ĩ �OULOOMB_u�0�wVISPITY��A�!OY�A_FR1Id��(�SI��B�R������3��
�W�W��0��09_,�EAS%��@�!�& "���4p�}G;� h ���7ƵCOEFF_AOm���m�/�G!2%�S.�߲CA5�����u�GR` � � $R� �X]�TME�$R�s�XZ�/,)�ER�T;��:䗰�  ]�LLt��S�_SV�&�($~����@�� "SETU��MEA��Z�x0��u������ � �� �� ȰID@�"���!*��&P���$*�F�'����)3��#���"�5;`:*��REC���!�7�SK_���� P	�1_USER��,��4���D�0��VEL,2�0���2�5S�I��0�MT�N�CFG}1� � ���Oy�NO�RE��3��2�0SI����� ��\�UX�-�ܑPDE�A $KEY_��}��$JOG<EנSVIA�WC�� 1�DSWy���
��CM7ULT�GI�@@�C��2� 4 p�#t�+�z�XYZ���쑡���z� �@_ERR��� ��S L��-���@��s0BB/$BUF-@X17�MOR�� H	�CU�A3�z�1Q��
��3���$��FV��2z��b�G�� � $cSI�@ G�0VO B<`נOBJE&�!F�ADJU�#EEL�AY' ���SD�WO�U�мE1PY���=0QT i�0�W�DIR$ba�pے�ʠDYN�HeT��@��R�^�X�����OPWORK}1��,�SYSBU@p 1SOP�aR�!�jU�k�PR��2�e�PA�0�!�cu� 1OP��UJ��a'�D��QIMAG�A�	��`i�IMACrI�N,�bsRGOVCRD=a�b�0�aP�`�sʠ� �^uz�L�P�B�@��!PMC�_E,�Q��N@�M��rǱ��1Ų7�=qS�L&�~0���$OVSL\G*E��*E2y�Ȑ�_=p�w�� >p�s���s	�����B8�t�#}1� @�@;����OE�RI#A��
 N��X�s�f�{�*�PL}1�,RTv�m��ATUSRBTRC#_T(qR��B ������$ �Ʊ��,�~0�C D��`-CSALl`��SA���]1gqXE@���%���C��J��
���UP(4����P!X��؆�q��3�w�� �PG�5�? $SUB�������t�JMPWAcITO��s��LOyCqFt�!D=�CVF	ш��y���R`�0��CC_CTR�Q�	�IGNR_PLt�/DBTBm�P��z�#BW)����0U@����IG�a��Iy�TNLN��Z�R]aK� !N��B�0�PE�s����r��f�SPD}1� L	�A�`gఠ�S���UN�{���]�R!�BDLY�2����7�PH_PK��E��2RETRI1Et��2�b���;FI�B� �����8� 2��0DB�GLV�LOGS�IZ$C�KTؑUdy#u�D7�_�_T1@�EM�@C\1A��ℽR��D�FCHE3CKK�R�P�0��e��@&�(bLEc�" PA9�T���P�C�߰PN�����A�Rh�0���Ӯ�PO��BORMATT naF�f1h���2�S���UXy`	�6�PL|B��4�  rE/ITCH��7�9�PL)�AL_ G� $��XPB�q�� C,2D�!��+2�wJ3D��� T�pPDCKyp��oC� �_ALPH���BaEWQo���� ��|I�wp � �b@?PAYLOA��m��_1t�2t���J3AR��؀դ֏�la�TIA4��5��6,2MOMCP������h�����0BϐAD��p������PUBk`AR��;���;������z4�` I$PI\Ds�oӓ1yՕ�w�T2�w�Z��I��I��I���p����n���y�e`�9S)bT�S/PEED� G��(� Е��/���Е�`/��e�>��M��ЕSAMP�6V��/���Е#MO�@ 2@�A�� QP���C��n������� ����LRf`kb�ІE9h�EIN09��7 S.В9
yPy�/GAMM%S���D$GET)bP�ciD]��2
�IB�:q�I�G$HI(0;�A��LREXPA8)LWVM�8z)��g���C�5�CHKKp]�0�I_��h`eT��n� q��eT,����� �$�� �1�iPI� RCH�_D�313\��30L�E�1�1\�o(Y�7 ¾t�MSWFL �M.��SCRc�7�@�&���%n�f�SV���PB``�'�!�B�sS_SAV&0ct5B3NO]�C\�C2^� 0�mߗ�uٍa��u� ��u:e;��1���8��D�P��������� )��b9��e�GE��3��V�e�Ml��o � �YL��QNQSRlbfq XG�P�RR#dCQpH� �S:AW70�B�B�[�CgR:AMxP�KCAL�H���W�r�(1n�rg�M�!o�� �F�P@}t$WP�u�P  r��P5�R<�RC� R��%�6�`��� �Ôqsr X��OD�qZp�Ug�ڐ>D� ��OM#w�J?\?n?@�?�?��9�b"�e�:]�_��� |��X 0��bf��qf��q`��ȏgzf��Eڐ� )	Ag�"�5���Fd�PB��PM�QU��� � 8L�Q�COU!h QTH�I�HOQBpHYSfY�ES��qUE�`t�"�O���  �1P�@\�UN���C�f�O�� P���Vu��!����OGSRAƁcB2�O�t�VuITe �q:pINFO�����{�qcB��e�OI�r� (�@SLEQS��q���p�vgqS����{ 4L�ENABDR>Z�PTIONt���p��Q���)�GCF��G�$J�q^r�� R���U�g��B�n�_ED����ѓ �F��PK���E'NU߇وA�UT$1܅COPY������n�00MNx���PRUT8R� �Nx�OU���$G[rf�e�RG�ADJ���*�X_:@բ$�����P��W��P��} ��)󂐶}�EX�YCDR[ ~�NS.��F@�r�LGO�#�NY�Q_FREQR�W`� �#�h�TsLAe#�����ӄ �CRE�� s�IF��sNmA��%a�_Ge#STATUI`e#MAIL�����q �t�������ELE�M�� �/0<�FEASI?�B��n��ڢ�vA�]� � I �p��Y!q]�t#A��ABM���E�p<�VΡY�BASR�Z���S�UZ��0$�q���RMS_TR ;�qb ���SY�	�ǡ���$���>C�Q`	~� 2� _ �TM������̲�@ ��A��)ǅ�i$DOUd�s]$Nj���PR+@z3���rGRID�q�M�BARS �TY�@�|�OTO�p��� Hp_}�!����d��O�P/�� � �p�`POR�s��}�.��SRV��)����DI&0T����� �#�	�#�4!�5!�6J!�7!�8�e�F��2��Ep$VAL�Ut��%��ֱ��/��� ;�1�q��1���(_�AN�#��ⓡRɀ(���TOTcAL��S��PW��Il��REGEN�1�cX��ks(��a����`TR��R��_!S� ��1ଃV�����⹂Z�E��p�q���Vr���V_H��DqA�S����S_Y,1��R4�S� AR�P2�� ^�IG_S!E	s����å_Zp���C_�Ƃ�ENHA�NC�a� T �;�������IN�T�.��@FPsİ_OVRsP�`p�`��Lv��o��7�}���Z�@�SLG�AA�~�25�	��D��YS�BĤDE�U�̦���TE�P���G� !Y��
�J��<$2�IL_MC�x r#_��`TQ�`��q����'�BV�C�P�_� 0�M�	V1V�
V1�2�2�U3�3�4�4�
 �!���� � m�A�2;IN~VIBP����1�2�2�3*�3�4�4�A@p-�C2���p� �MC_Fp+0B�0L	11d���M501Id�%"E� S`�R�/�@KEEP__HNADD!!`$$^�j)C�Q���$��"	��#O�a_$A�!pK��#i��#REM�"��$��½%�!�(U�}�e�$HPWD � `#SBMSUK|)G�qU2:��P	�COLLAB � �!K5�B�� ��g��pITI1{9p#n>D� ,�@FLAP>��$SYN �<�M�`C6���UP�_DLYAA�ErDGELA�0ᐢY�`�AD�Q��QSwKIP=E� ���XpOfPNTv�A�0P_Xp�rG�p�RU@ ,G��:I+�:IB1:IG� 9JT�9Ja�9Jn�9J{к9J9<��RA=s� X���4�%1�Q}B� NFLIC�s��@J�U�H�LwNO�_H�0�"?��RIT�g��@_PA�pG��Q� �K�^�U�W��LV�d�NGRLT�0_q��O�  p" ��OS��T_JvA� V	�APPR_W�EIGH�sJ4CH?pvTOR��vT���LOO��]�+�tVJ�е�ғA�Q�U�S�X�OB'�'���J2TP���7�X�T� <a43DP=`Ԡ\"<a�q�\!��RDC��L�+ �рR��R�`� ��RV��jr�b�R�GE��*��cN�FL�G�a�Z���SPC��s�UM_<`^2�TH2NH��P.a �1� m`EFv11��� lQ `�!#� <�p3AT�  g�S�&�Vr�p�tMq�Lr���HOME(wr�t2'r�-?�Qcu��w3'r逪������w4'r�'�9�K�]�o���
�w5'r뤏��ȏڏ(����w6'r�!�3��E�W�i�{��w7'r퀞���ԟ����w8'r��-�?�Q�c�u�R�uS$0�q�p�� sF��`la�!`P�����`/���-�IO[M�I֠��q�POWE�� ���0Za*��� ��5��$DSB� GNAL���0C�pm�S2323�� �~`��� / I3CEQP��PEp���5PIT����OPB�x0��FLOW�@T�RvP��!U���CU:�M��UXT�A��>w�ERFAC�� �U����ʱC�H��� tQ  _���>�Q$����O)M��A�`T�P#�UPD7 A�ct�T��UEX@�ȟ�U �EFA: X"�1RS9PT�����T ���PPA�0o񩩕`EXP�IOS���)Ԃ��_���%��C�WR�A��ѩD�ag֕`~ԦFRIENDsa�C2UF7P����TO;OL��MYH C2�LENGTH_V�TE��I��Ӆ�$SE����UFI�NV_���RsGI�{QITI5Bb��Xv��-�G2-�G17�w�SG�X��_��UQQD=#���AS��d~C�`��qᾭ� �$$C/�S�`����� )`|����VERSI� ���)`�5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����� ����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT��C��  ��DI�N�O�A�Dq�EXE��HPV_��AT�Qz
��LARM�RECOV ��RgLMDG �*�5�OLM?_IF *��`d�O�_�_�_�_j�_�'o9oKo]onm, 
��odb��o�o�o0�o^��$� z, �A   2D{�P�PINFO u[ �Vw��������`����� ��*��&�`�J���n�����DQ���� 
��.�@�R�d�v���𚟬���a
PPLI7CAT��?�P���`Ha�ndlingTo�ol 
� 
V�8.30P/40�Cpɔ_LI
8�83��ɕ$ME�
F0G�4�-
?
398�ɘ��%�z�
7�DC3�ɜ
�No+neɘVr���ɞ_@6d� ~Vq_ACTIVU���C죴�MOD�P���C�I��HGA�PON���O�UP�1*�� Ai�m����Қ_��6��1*�  �@��������Q����Կ�@�
���=�� ���5��Hʵl�K�HTTHKY_��/�M� SϹ���������%� 7ߑ�[�m�ߝߣߵ� ���������!�3�� W�i�{�������� ������/���S�e� w��������������� +�Oas� ������ '�K]o��� �����/#/}/ G/Y/k/�/�/�/�/�/ �/�/�/??y?C?U? g?�?�?�?�?�?�?�? �?	OOuO?OQOcO�O �O�O�O�O�O�O�O_ _q_;_M___}_�_�_��_�_�_�_kŭ�TO�p��
�DO_CL�EAN9��pcNM  !{衮o�o��o�o�o��DSP�DRYRwo��HI��m@�or��� ������&�8�J���MAXݐWdak�H�h�XWd�d��>�PLUGGW�Xg\d��PRC)pB�`E�kaS�Oǂ�2DtSEGF0�K � �+��o�or�����p�����%�LAPO b�x�� �2�D�V�h� z�������¯ԯ�+�TOTAL����+�_USENUO�\�� e�A�k­�RGD�ISPMMC.�2��C6�z�@@Dr\��OMpo�:�X�_S�TRING 1	~(�
�M!��S�
��_ITwEM1Ƕ  n� �����+�=�O�a� sυϗϩϻ����������'�9�I/�O SIGNAL���Tryou�t Modeȵ�Inpy�Simu�lateḏO�ut��OVE�RRLp = 10�0˲In cy�cl�̱Pro?g Abor��̱�u�Status�ʳ	Heartb�eatƷMH �Faul	��Aler�L�:�L�^�p����������� ScûSaտ��-�?� Q�c�u����������� ����);M_q��WOR.�û� �����+ =Oas��������//'.PO����M �6/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�?8�?�?H"DEVP.�0 d/�?O*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8_J_\_n_PALT	��Q�o_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o8�o�_GRIm�û 9q�_as��� ������'�9� K�]�o�������'�R	�݁Q����)� ;�M�_�q��������� ˟ݟ���%�7�I�ˏPREG�^���� [�����ͯ߯��� '�9�K�]�o�������෿ɿۿ�O��$A�RG_� D ?	����0���  	]$O�	[D�]D���O�e�#�SBN_�CONFIG �
0˃���}�C�II_SAVE � O�����#�T�CELLSETU�P 0�%  ?OME_IOO�O�%MOV_H������REP��J��UTOBACK�����FRwA:\o� Q�,o���'`��o����� ��  f�o�����*�!�3�`��Ԉ��f���� ������o�{��&�8� J�\�n���������� ��������"4FX j|�������끁  ��_�i�_\ATBCK�CTL.TMP �6.VD GIF? .TP D_xq��N.E#��.f�INI�P�Օ��c�MESSAG�����8��ODEC_D����z��O�0��c�PAUSM!!��0� ((O 3�U/g+Q/�/u/�/�/ �/�/�/�/�/)??M?�;?q?70$: TSK�  @-��T�f�UgPDT��d�0�
&XWZD_ENqB����6STA��0��5"�XIS��U�NT 20Ž�� � 	�? ,"�>UO��oO�O�O�O��O�O_�O&_�7AM[ET߀2CMP_  ?��Od_�_0E�SCRDCFG }1�6��	��Ź��_�_oo (o:oLo��o�Q���_ �o�o�o�o�o�o]o �o>Pbt���o9�i�GR<@M/��s/NA�/�	�i��v_ED�1��Y� 
 �%{-5EDT-��'�GETDAT�AU�o�9��
�-(i�H�o�f�\�ּA��  ���2 �&�ȏE�D���~� ŏ׏m����3��&� �J�\�ߟJ�����9�ǟ�4���ϯ�\�����]�o�����5 N������\�w��)�;�ѿ_��6ϊ�g� ��\�CϮ���ϝ�+��7��V�3�z�\��@z�����i����8������]���F� �ߟ�5����9~������]����Y�k�����CR�!ߖ� ��W�q���#�5���Y���p$�NO_DEL���rGE_UNU�SE��tIGAL�LOW 1���(*SYS�TEM*}S	$SERV_GR��}V� : REG�q$�}\� NUM�
<��PMUB }U�LAYNP}\PMPAL�>CYC10#6� $\ULSU`�8:!�Lr~�BOXORI��CUR_��PoMCNV��10L�T4DL!I�0��	����B N/`/r/�/�/�/�/�/����pLAL_OU�T �;���qW?D_ABOR=f��q;0ITR_RT�N�7�o	;0NON�S�0�6 
HCC�FS_UTIL s#<�5CC_@�6A 2#; h� ?�?�?O#O�]CE�_OPTIOc8�qF@RIA_IIc f5Y@�2�0�F�Q�={]2qނA_LIM�2�.� ��P��]B���K}X�P
�P�,2O�Q��B�r�qF�PQ5T1)TR�H�_:JF_PA�RAMGP 1�<g^&S�_�_�_��_�VC�  C��d�`�o!o`��`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?���2HE ONFI�� E?�aG_P�1#; ���o 1CUgy�a�KPAUS�1�yC ,���� �����	�C�-� g�Q�w���������я4���rO�A�O�H~�LLECT_�B1�IPV6�EN. QF܍3�NDE>� ��G�71234567890���sB�TR����%
 	H�/%)����� ��W���0�B���f�x� ��㯮���ү+���� �s�>�P�b������� ���ο��K��(Ϡ:ϓ�^�|��B!F�� �I|�IO #��<U%e6�'��9�K���TR�P2$���(9X�t�Y޼`�%�̓ڥH��_MO-R�3&�=��i� �A�$��H�6�l�Z���~S��'�=�r_A? �a�a`��@K��RʭdP��)F�haÃ-�_�'�9�%
@�k��G� ��%Z�^%��`�@c.��PDB��+���cpmidbg��X	3 :�`@`@�QU��p��N�  �����)X���]�`@sX<�^��@�s�g�$� �sf�l�q��ud�1:��:J��DE�F *ۈ��)��c�buf.t�xt����_L�64FIX , ������l/[Y/�/}/ �/�/�/�/
?�/.?@? ?d?v?U?�?�?�?�?��?�?,/>#_E -���<2ODOVOhOXzO�O6&IM��.o�=YU>���d�
�6IMC��2/���ñdU�C��20�M��QT:Uw�Cz  B��i�74<�8���7@@�7(�8�CG�7�0�w�i�9;���9��9;�
>�PD�%�Qs]�=7[3=e3D�=7Y=7X��E\=7Wްw��D4'��22o��D|����� �𺪢�C�C���e�
�xObi�D4cdv`D��`/�`v`s]�E�D D�` �E4�F*� ?Ec��FC��u[�F���E��f�E��fFކ3�FY�F�P3��Z��@�33 ;?��>L���Aw��n,a@��@e�5!Y���a���`A��w�]=�`<#ךW�?��oyJRSMOFST (�,bI+T1��D @3��
�e�rQ
�a��;��b�w?���<��M�NTESTR�1O�CR@�4�4�>VC5`A�w�Ia�+a�aORI`CTPB͖U�C�`4����r��:d����qIj?�5��qT_�?PROG ��
��%$/ˏ�t��NUSER  k��������KEY_TBL'  ����#a��	
��� !"�#$%&'()*�+,-./��:;�<=>?@ABC��GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?�����������LCK�
����S�TAT/��s_AU�TO_DO ��	�c�INDT_ENBP���Rpqn�`�sT2����STOr`쓯�XC�� 26����8
SONY XC-56��"b����@��F(� А�H�R50w���>�P�7<b�t�Aff����ֿ� Ŀ����C� U�0�yϋ�fϯ��Ϝ���������-ߜ�TR�L��LETEͦ ���T_SCRE�EN ���kcs���U�MMENU 17�� <ܹ���w� ��������K�"� 4��X�j������ ������5���k�B� T�z������������� ��.g>P� t������ Q(:�^p� ���/��;// $/J/�/Z/l/�/�/�/ �/�/�/�/7?? ?m? D?V?�?z?�?�?�?�? �?!O�?
OWO.O@OfO��OvO�O�O(y��RE�G 8�y�����`�M�ߎ�_MAN�UAL�k�DBC�O��RIGY�9�DBG_ERRL��9�ۉq��_�_��_ ^QNUML�I�pϡ�pd
�
�^QPXWORK 1:���_5oGoYo�ko}oӍDBTB_NN� ;������ADB_A�WAYfS�qGC�P 
�=�p�f_A!L�pR��bbRY�[�t
�WX_�P 1<{y�n�,�%oc�Pl��h_M��ISO���k@L��sONTImMX��
���v�y
��2sMOTN�END�1tREC�ORD 1B��� ���sG�O� ]�K��{�b�������� V�Ǐ�]����6�H� Z���������#�؟ ������2���V�ş z��������ԯC��� g��.�@�R���v�� ��	���п���c�� ��#ϫ�`�rτϖ�� ��)ϳ�M���&�8� ��\�G�Uߒ�߶��߀��I������4��  �p7�n���ߤ��� ������"���F�1� ��|��������[��� ��i���BTf����bTOLERE�NC�dB�'r�`L���^PCSS_CCSCB 3C>y�`IP�t}�~� <�_`r�K������/�{� �5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O��O_�~�LL� D���&qET�c�ao C[C��P�ZP^r_ A� p� �sp��QGPt[	 A�p�Q�_�[A? �_�[oU�pc�P�pSB�V �c�(a�PWoio{h+
�o�h�o�oY���[	r�hLU�tNH��8*��3J72ܘߊ�c��aD�@VB��|�G����+��K� �otGhXGrcso����e�B   =���2�a>�tYB�� �pQC�p�q�aA"�H�S �Q-��q���ud�v������AfP ` 0����D^P��p@5�a
_�XTHQH����a aW>� �a9P��b�e:�L�^� h�Hc�́PQ�RFQ �PU�z�֟�o\^� �-�?��c�u���zCz�ů�b2x�Щ�RD��r��y�G����S̡0� �]�0�.��@���EQ�p��F�X�ѿUҁ�п�VSȺNST�CY 1E��]�ڿ��K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߒ���DEVICE ;1F5� MZ�� �a��	� ��?�6�c���	{䰟���_HNDGD G5��VP���R�LS 2H�ݠ��/�A�S�e��w����� ZPARA�M I�FgHe~�RBT 2K�܋8р<��WPpCU�C��,`¢P�Z��z��%{�C*  �2�jMTLU,`"nPB, s� �M� }�gT�g��
#B��!�bcy� [2Dchz�����/��/gT#�I%D��C�` �b!�R��A��A�,��Bd��A5��P��_C4kP�!�2�C��$Ɓ�]�f�fA�À��B�� �| ���/�/�T (��54a5�} %/7/d?/M?_?q? �?�?�?�?�?O�?O O%O7OIO�OmOO�O �O�O�O�O�O�OJ_!_ 3_�_�_3�_�_�_�_ �_o�_(ooLo^oЁ =?k_IoS_�o�o�o�o �o�o�o#5G �k}����� ��H��1�~�U�g� y�ƏAo�Տ���2� D�/�h�S���go���� ԟ����ϟ���R� )�;���_�q������� ���ݯ�<��%�7� I�[�m��������� }�&��J�5�n�Yϒ� �Ϗ��ϣ�ѿ���� ��F��/�Aߎ�e�w� �ߛ߭���������B� �+�x�O�a���� ��������,���%�b� M���q����������� ����L#5� Yk}��� � �61CUg �������� 	//h/���/w/�/�/ �/�/�/
?�/.?@? I/[/1/_?q?�?�?�? �?�?�?�?OO%OrO IO[O�OO�O�O�O�O �O&_�O_\_3_E_W_ �_?�_�_�_�_�_"o oFo1ojoE?s_�_�o m_�o�o�o�o�o0 f=Oa��� �������b� 9�K���o���Ώ��[o ��(��L�7�I����m������$DCS�S_SLAVE �L���ё���_4D�  љ��CFoG Mѕ��������FR�A:\ĐL-�%0�4d.CSV�� � }�� ���A Vi�CHq�z����p��|�����  ������Ρޯ̩ˡҐ-矩*����_CR�C_OUT N�������_FS�I ?њ ����k�}����� ��ſ׿ �����H� C�U�gϐϋϝϯ��� ������ ��-�?�h� c�u߇߽߰߫����� ����@�;�M�_�� ������������� �%�7�`�[�m���� ������������8 3EW�{��� ���/X Sew����� ��/0/+/=/O/x/ s/�/�/�/�/�/�/? ??'?P?K?]?o?�? �?�?�?�?�?�?�?(O #O5OGOpOkO}O�O�O �O�O�O _�O__H_ C_U_g_�_�_�_�_�_ �_�_�_ oo-o?oho couo�o�o�o�o�o�o �o@;M_� �������� �%�7�`�[�m���� ����Ǐ������8� 3�E�W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿� ��'�P�K�]�oϘ� �ϥϷ���������(� #�5�G�p�k�}ߏ߸� ������ �����H� C�U�g������� ������ ��-�?�h� c�u������������� ��@;M_� ������� %7`[m� ������/8/ 3/E/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO�sO�O�O�O�O�C�$�DCS_C_FS�O ?�����A P �O�O_?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo ~o�o�o�o�o�o�o�o 72DVz� ������
�� .�W�R�d�v������� ������/�*�<� N�w�r���������̟ ޟ���&�O�J�\� n���������߯گ� ��'�"�4�F�o�j�|� ������Ŀֿ�������G�B�T��OC_RPI�N_jϳ��� �ς��O����1�Z�U��NSL��@&�h߱� ��������"��/�A� j�e�w������� ������B�=�O�a� ���������������� '9b]o� ������� :5GY�}�� ����///1/ Z/U/g/y/�/�/�/�/ �/�/�/	?2?-???Q? z?u?��ߤ߆?�?�? �?OO@O;OMO_O�O �O�O�O�O�O�O�O_ _%_7_`_[_m__�_ �_�_�_�_�_�_o8o 3oEoWo�o{o�o�o�o �o�o�o/X Sew����� ���0�+�=�O�x� s���������͏ߏ� ��'�P�K�]�o������ �PRE_CH�K P۫�A ~��,8�2x��� 	 8�9�K���+�q���a� ������ݯ�ͯ�%� �I�[�9����o��� ǿ��׿���)�3�E� �i�{�YϟϱϏ��� ��������-�S�1� c߉�g�y߿��߯��� �!�+�=���a�s�Q� ����������� ���K�]�;�����q� ������������#5 �Ak{�� ����CU 3y�i���� ��/-/G/c/u/ S/�/�/�/�/�/�/? ?�/;?M?+?q?�?a? �?�?�?�?�?�?�?%O ?/Q/[OmOO�O�O�O �O�O�O�O_�O3_E_ #_U_{_Y_�_�_�_�_ �_�_�_o/ooSoeo GO�o�o=o�o�o�o�o �o=-s� c������� '��K�]�woi���5� ��ɏ��������5� G�%�k�}�[������� ן�ǟ����C�U� o�A�����{���ӯ�� ��	��-�?��c�u� S�������Ͽ῿�� ���'�M�+�=σϕ� w�����m������%� 7��[�m�K�}ߣ߁� ���߷����!���E� W�5�{��ϱ���e� ������	�/��?�e� C�U������������� ��=O-s� ���]���� '9]oM�� �����/�5/ G/%/k/}/[/�/�/� �/�/�/�/?1??U? g?E?�?�?{?�?�?�? �?	O�?O?OOOOuO SOeO�O�O�/�O�O�O _)__M___=_�_�_ s_�_�_�_�_o�_�_ 7oIo'omoo]o�o�o �O�o�o�o!�o1 W5g�k}�� ����/�A��e� w�U�������я��o ����	�O�a�?��� ��u���͟����� '�9��]�o�M����� ����ۯ��ǯ�#�ů G�Y�7�}���m���ſ �����ٿ�1��A� g�E�wϝ�{ύ����� ��	�߽�?�Q�/�u� ��e߽߫ߛ������� �)���_�q�O�� ������������ 7�I���Y��]����� ����������!3 WiG��}�� ��%�A�1 w�g����� �/+/	/O/a/?/�/ �/u/�/�/�/�/? �/9?K?�/o?�?_?�? �?�?�?�?�?O#OO GOYO7OiO�OmO�O�O �O�O�O_�O1_C_%? g_y__�_�_�_�_�_ �_�_o�_+oQo/oAo �o�owo�o�o�o�o �o);U__q� �������%� �I�[�9����o��� Ǐ�����ۏ!�3�M ?�i��Y�������՟ �ş����A�S�1� w���g�����������ӯ�+�=��$DC�S_SGN Q�K�c��7m� �14-JAN�-19 08:3O8   O�l� ����� N.D�Ѥ���������h��x,rWf*σ��^M��  O�V�ERSION �[�V3.5�.13�EFLO�GIC 1RK���  	���P�?�P�N�!��PROG_ENB  ��6Ù�o�ULSE  T����!�_ACCL{IM���������WRSTJN�T��c��K�EM�Ox̘��� ���INIT S.�G�Z����OPT_SL �?	,��
 	�R575��Y�7�4^�6_�7_�50
��1��2_�@ȭ��><�TO  Hݷ�t��V�DEX���dc����PAT�H A[�A\��g�y��HCP_�CLNTID ?<��6� @ȸ�����IAG_GR�P 2XK�? ,`��� � �9�$�]�H������123456�7890����S�� |�������!�� ��H���;� dC�S���6� ����.�R v�f��H� �//�</N/�"/ p/�/t/�/�/V/h/�/ ?&??J?\?�/l?B? �?�?�?�?�?v?O�? 4OFO$OjO|OOE� �Oy��O�O_�O2_��@_T_y_d_�_,
�B^ 4�_�_~_`Oo �O&oLo^oI��Tjo�o .o�o�o�o�o �O' �_K6H�l�� �����#��G��2�k�V���B]�?��  �~�x6�븊������2޽�*�iƁD|��8���DR��8�Ƈ����(���L�B\ډ�4  �?}��dI�C� ���������ϟ����ICT_CONF_IG Y���>��egU����STBF_TTS��
��b����Û�u�O�MAU��|�MSW_CF6�Z���  �OCV7IEW��[ɭ������-�?�Q�c� u�G�	�����¿Կ� �����.�@�R�d�v� ϚϬϾ�������� ��*�<�N�`�r߄�� �ߺ���������&� 8�J�\�n���!�� �����������4�F�`X�j�|����RC£	\�e��!*�B^�������C2g{�S�BL_FAULT� ]��ި�GP�MSKk��*�TD?IAG ^:�ա�I��UD1�: 6789012345�G�BSP�-?Qcu� ������//�)/;/M/tJ��
@�q��/$�TREC	P��

��/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO�0OBOi/{/xO�/UM�P_OPTIONk���ATR¢l��	��EPMEj��OY�_TEMP  ?È�3B�J�Ps�AP�DUNI���m�Q��YN_BR�K _ɩ�EMGDI_STA"U��aQSUNC_S1`ɫ �FO�_�_�^
�^dpOoo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{�E�����y �Q��� �2�D�V� h�z�������ԏ� ��
��.�@�R�d��z �������˟��� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i��������� ÿݟ�����/�A� S�e�wωϛϭϿ��� ������+�=�O�a� {�iߗߩ߻�տ���� ��'�9�K�]�o�� ������������� #�5�G�Y�s߅ߏ��� ��i�������1 CUgy���� ���	-?Q k�}�������� �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?u?�? �?�?��?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_m?w_�_�_�_�?�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9Ke_W� ���_�_���� #�5�G�Y�k�}����� ��ŏ׏�����1� C�]oy�������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;���g�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�_�i�{ߍߟ߹� ����������/�A� S�e�w������� ������+�=�W�E� s������ߧ������� '9K]o� ������� #5O�a�k}�E ������//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-?GY c?u?�?�?��?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_Q?[_m__�_ �?�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/I_ Sew��_��� ����+�=�O�a� s���������͏ߏ� ��'�A3�]�o��� ����ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����9� K�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ���ߑ�C�M�_�q� �ߝ��߹�������� �%�7�I�[�m��� ������������!� ;�E�W�i�{��ߟ��� ��������/A Sew����� ��3�!Oa s�������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? +=G?Y?k?!?��? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	_#?5??_Q_ c_u_�?�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o -_7I[m�_� �������!� 3�E�W�i�{������� ÏՏ����%/�A� S�e�q�������џ �����+�=�O�a� s���������ͯ߯� ���9�K�]�w��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����������'�1� C�U�g߁��ߝ߯��� ������	��-�?�Q� c�u��������� ��m��)�;�M�_�y� �������������� %7I[m� �������! 3EWq�{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/�/+?=?O?i _?�?�?�?�?�?�?�? OO'O9OKO]OoO�O��O�O�O�O�O�O? ��$ENETMO�DE 1aj5�  0�054_F[PR�ROR_PROG %#Z%6�_�Y�dUTABLE  #[t?�_�_�_g�dRSEV_NUM� 2R  ��-Q)`dQ_AUT�O_ENB  �PU+SaT_NO>a �b#[EQ(b W *��`��`��`	��`4`+�`�o�o�oZdHIS%c1+PSk_ALM 1c#[� �4�l0+�o;M_q��r�o_b``  #[�aFR�zPTCP_VER !#Z�!�_�$EXTL�OG_REQ�f9�Qi,�SIZ5�'��STKR�oe�~)�TOL  1{Dz�b�A '�_BWD�p��Hf���D�_DI�� dj5SdDT1KRņSTEPя�P���OP_DOt�QF�ACTORY_T�UN�gd<�DR_?GRP 1e#YNa�d 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ�ԟ ���1��U�@�y�d��v�����ӯ����LW
? I�kn�,��tۯ�j�U���y��B�  B୰�>��$  A@��s�@UUUӾ����Ͼ��E�� E�`F@ F�5U/��,��L���M���Jk�Lz�p�JP��Fg{�f�?�  s���9�Y9}��9��8j
��6��6�;���l����z �!� �� Q�)������[FEATUROE fj5��JQ�Handl�ingTool �� "
P�English �Dictiona�ry�def.�4D St�a�rd�  
! �hAnalo�g I/OI�  �!
IX�gle� ShiftI�d��X�uto So�ftware U�pdate  r�t sѓ�mati�c Backup~�3\st���ground E�dit��fd�
Camer�a`�Fd�e��Cn?rRndIm����3�Common� calib U}I�� Ethe��n��"�Monit{or�LOAD8��tr�Relia�by�O�ENS�Da�ta Acquiys>��m.fdp�?iagnos��]��i�Document VieweJ���870p�ua�l Check �Safety*� �cy� �hanceod Us��Fr�����C �xt. oDIO :�fi��s m8���end��ErrI�L��S�������s  t P%a�r[�� ����J944FCTN Menu��ve�M� J9l�T�P InT�fac�{�  744��G���p Mask �Exc��g�� R�85�T��Pro�xy Sv��  �15 J�igh�-Spe��Ski>
� R738Г�~�mmunic���ons�S R7���urr�T�d�02�2��aю�conn�ect 2� J�5��Incr��s�tru,Қ�2 R�KAREL �Cmd. L��u�a��R860hR�un-Ti��En�vL�oa��KU�e�l +��s��S/�Wѹ�7�Lice�nse���rod�u� ogBook�(System)��AD pM�ACROs,��/�Offs��2�NDFs�MH�� �����MMRC�?��O�RDE� echS�top��t? � 84fMi$�|� 13dx��]е��܏���Modz�witchI�VP��?�:��. sv��2Optm�8�2���fil��I ��2g� 4 !+ulti-T�����;��PCM funY�Po|���4$��b&Regi� r\ �Pri��FK+�7���g Num �SelW  F|�#�� Adju����60.��%|� �fe���&tatuď!$6���%��  �9 J6RDM Robot)��scove2� 5;61��RemU�=n@� 8 (S�F3Servo�����)SNPX� b�I�\dcs<�0}�Libr1��OH� �5� fl�0��58��So� =tr�ssag4%G /91�p ���&0���p/I�� � (ig TMIL�IB(MӋ�Firm����gd7���s�'Acc����0�XAsTX�Heln���*LR"1��Sp�ac�Arquz�iOmulaH��� Q�n��Tou�Pa�D�I��T��c��&���ev. f.sv�USB po���"�iP�a�� � r"1Unexcept��`0i$/���n�H59� VC&�r��[6���P{�<�RcJPRIN�V�;� d T@�TSP� CSUI�� r��[XC��#Web� Pl6�%d -c�1R�@4d������I�R66?0FV�L��!FVGridK1play C�lh@X����5RiR�R.@�~��R-35iA|���Ascii��8�"��� 51f�c�Upl� � (T�����S��@rit�yAvoidM l�`��CE��rkδCol%�@�Gu"F� 5P��j}P�����
 B�L�t� 120C C� o�І!J�D�P��y��� o=qz�b @DCS b ./��c��O��q��D`�; ���qckpgaboE4�DH@��OTШ�main �N��1.�H��an�.��A> aB!FR�LM���!i ���M�I Dev�  (�1� h8j��spiJP��� �@��Ae1�/�r���!hP� M-2� i��߂^0ii�p6�PC���  iA/'�Pa�sswo�qT�RGOS 4����qedav�SN��Cli����G6x Ar�� �47�!���5s�DsER��Tsup>Ryt�I�7 (M�aΪT2DV�
�3D Tri-���&���_8;�
�A�@D�ef?����Ba�: deRe p 4�t0��e�+�V�s�t64MB DR;AM�h86΢�FRO֫0�Arc�� visI�ԙ�n<��7| ), �b��Heal�wJ�\h���Cell`��p� �sh[��� Kq:w�c� - �v�b��p	VCv�tyy�ys�"Ѐ6�u�t��v�m���xs ���TD_0��J�m㖙` 2��a[�>R �tsi�MAILYk�/F2�h��ࠛ 90 H��F02�]�q�P5'���T10C��5����FC��Uz�F9�GigEH��S�t�0/A� if��!2��boF�dr�i=c �OL�F�S����" H5�k�OPT ��4�9f8���croP6��@��l�ApA��Syn.(RSSG) 1L�\1y�rH�L� (2x5�5�d�p�CVx9����estb�$SР��> \pϐ�SSF�e$�tex�D o���A�	� �BP���a�(R00��Qirt��:���2@)�D��1�e�VKb@_l Bui, n��WAPLf��0��1Va�kT�XCGM��D���L����[CRG�&a�YBU��YK�fL��pf��k�\sm�ZTAf�@�О�Bf2�и��V#�s�d��� r���CB��@�
f���WE��!!��
���T�p��DDT�&4 Y�V�`��EH����
�#61Z��
�R=2�
&�E (Np��F�V�P K�B���#��Gf1`?G���H�р?eI�e ����LD�4L��N��7\s@����`���M��deSla<,��2�M�� "L[P��`?@��_�%�����S��M-F�TSO�W�wJ57��VGF��|�VP2֥ 5\ b�`0&�cV:���T;�T� �<�ce,�?VPD��$
eT;F��DI)�<�I�a\so<��a-�6Jc6s6�4L�M�bV9R�h���Tri� � ���5�` �f�@�������P
� ����`>��Img PH�[�l��I/A  DVP�S��U�Ow���!%S�Skastdp�n)ǲt�� SWI�MEST�BFe�00��-Q� �_�PB�_�Rued�_�T��!�_�S ��_bH573o2c2��-oNbCJ5N�Iojb)�Cdo�cxE��o�_�lp��o �TdP�o�c�B�or�2 .rٱ(Jsp�Efr�SEo�f1�}�r3s RGoeELS��sL����s������B	��S\ $�F�ryLz�ftl�o~�g�o ���������?������P  �n�&�"�l  ��T�@<�^��Y��e��u8Z���alib��Γ��ɟ3����f��\v ��e\c��6�Z�f�T�v�R �VW���8S��UJ9�1����i�ů[c91�+o�w8���847�:��A4�j��Q���t6�m���vrc.�����HR���ot8�0ݿ��  ���8ޯ�460�>eS0L�97���U���Ϧ�60.� g�н�@+��'�ܠ�Ϻ�8co&��DM߱U"����d�ߕpi�߲T! �&�na;�� ���u%��ⅰI��lo`R�d��1a59gϘ�ŭ���95�ϔ�R����1��?��o�#� �1A�/���vt{�U�Weǟ���ￇ73�[���7�ρ�C WL��62K�=fR���8��������d����2�ڔ����@��@" "http�����t7 ��� v R7��78�����4�� ��TT�PT�#	��eP#CV4/v߀�j�Q�Fa7��$N�0�/2��rIO�)/;/M/6.sv3�64i�oS�l? torah?*�|`�?��AM/�?
??p.?0�k/��1 JO0��� ,O�tro���0[P��OB4c.K?�g�'�)�24g?�� (1B�Od�\iOA5csb�?U_�?vi�/i��/�/Wn��`�o%�Fo�4l�$of���oXF I)xo�cm3p\7��mp���d�uC��lh����o(AA�_Bt� �o]6P���m�I?�w�@���na$O��4*O0wi�8%P�?"�bsg?�]7��YEM���8woVJ̇/ե11?o��DMLs�BC��7J��\���(�52�XFa AP�ڟ<�v�`/ş�aqs����/OIf��1�9��VRK���ph�քH�5+�=�IN/¤SckiW�/�IF�0�_�%��fs�I�O�l����"<𜿚$�`����\jԿz5bON�vrouς�3(�ΤH (DϮ��?sG ��|��F�Ou������ �D)O��*�3P$� FӅ�k��ϻ���럴�� �PL��ʿ��pb3ox�ߦebo����Sh �>�R.�0wT{����fx6��P���D��3��#_I\Im;YEe�OԆM�8hxW�=Ete,���dGct\���O$kR�������Xm*���r�o3��D�l�j9���V'�  FAC���|@�ք f?6KARE0�_�~� (Kh��.cf���WpoO�_K�up��a���H/j#�- Eqd/�84���$qu�o��/ o2o?Vo<�7C�)�s��NJԆ�|?�3l\�sy�?�40�?Τwaio�u]?�w58�?�,F�$OJ�
?Ԇ"Iio�!�V��u&A�f�PR�ߩ5, s���v1\  �H552B�Q2�1p0R78�P510.R0 � nel J�614Ҡ/WATUP��d8PW545*�H8R6��9VCAM�q97PCRImP\1tP�UIF�C8Q28  ingsQy0��4P� P63P @P PS�CH��DOCqVڀD �PCSU���08Q0=PqpV�EIOCr��� P5�4Pupd�PR6q9aP���PSET�p�t\hPQ`Qt�8P7�`Q�!MASK���(PPRXY䞓�R7B#POCO�  \pppb3 6���PR�Q��b1Pdy60Q$cJ539.e�Hsb��vLC�H-`(�OPL-Gq\bPQ0]`��P(`HCR��4`�S�aund�PMCISIP`e0aPle5=P9s�p(`DSW� � � qPb0`�aPa��(`P�RQ`Tq�RE`(Poa6901P<cPCM�PHc{R0@q\j23b��V�`E`�S`UPvisP`E` c�`UPc�PRS	a�bJ69�E`sFRDmPsRwMCN:eH931P�HcSNBARa�rHLB�USM�qc�Pvg52�fHTCIP0cTMIL�e"P�`�eJ �PA�PdST�PTX6p967PTEL�p��P�`�`
Q8P8$Q48>a"PP�X�8P95�P`[�9�5qqbUEC-`F;
PUFRmPfa�hQCmP90ZQVCqO�`@PVIP%�w537sQSUIzVsSX�P�SWEBIP��SHTTIPthrFQ62aP�!tPG����cIG؁�`c�P;GS�eIRC%��c'H76�P�e Q�Qr|�Ror��R51P0 s:P�P,t53=P8u)8=Py�C�Q6]`0�b�PI��q52]`sJ56E`s���PDs�CL�qPt5�\r�d�q75UP cR8䀑�u5P sR55 ]`,s� P8s��P�`pCP�PP�SJ77P0\o�6��cRP,P�cR6�ap�`�Q�taT�79P`�64̑Pd87]`�d90�P0c��=P,���5�9,ta�T91P� ��p1P(S���Qpai�P�06=P- C�PF��T	���!aLP PT�S�pL�CAB%�I БIQ` ;�H�UPoPaintPMS�P�a��D�IP|�STY�%�t\patPTO��b�P�PLSR76č`�5�Q��WaNNn�Paic�qNNE`��ORS�`�cR6�81Pint'�FC�B�P(�6x�-W`M��r��!(`OBQ`p�lug�`L�aot �`OPI-���P�SPZ�PPG�Q7v�`73ΒPRQ�ad�RL��(Sp�PS��n�@�E`o�� �PTS-�ǈ W��P�`ap�w�`��P`cFVR��PlcV3D%�l�PsBVI�SAPL�Pwcyc+PAPV1��pa_�CCGIP �- U��L�Prog+PCCR�`�ԁ�B�P �PԁK=�"!L�P��p��(h�<�AP��h�̱�@g�Bـ�
TX�%���CTC�ptp��2��P927"0ҝPs2��Qb��TC-�rmtl;�	`#1ΒTC9`nHcCTE�Perj�]EIPp.p/�E�P��c��I�use��F�ـvrv�F%���T�G�P� CP��%�d u-h�H-�Tra�PgCTI�p��TL� TRS���p�@נ���IP�PTh�M%�l�exsQTMQ`ve#r, �p�SC:���F��Pv\e�PF�IPSV"+�H�$cj�ـ;tr�aCTW-����CPVGF-��SVP=2mPv\fx���pac�b��e��bVP4яfx_m��-��SVsPD-��SVPF�P�_mo�`V� cV֣�t\��LmPov�e4��-�sVPR��\|�tPV�Qe5.W`V6�*u"��P}�po`���`��CVK��2N�IIP��CV�����IPN9�Gene ���D��D�R�D�����  ��f谔�po{s.��inal��n��DeR���`���d�P��omB���o�n,���R�D�R��\���TXf��D$b��o;mp�� "N��P2��m���! ��=�C-f����=FXqU�����g F��<(��Dt II��r4�D��u�� "����Cx_ui X������f2��h	C�rl2��D,r9ui��Ԣ� it2cl�0co��e"�����ا(.)�� ���� ��{� IQnQ ��I[ ��_�= wo��,b{D� ��|�GG� �����4 �e�� vʷ� ���&� 2��Z� uz������� ��TW&q�~q 5�׷&��o? ;0���  �2� ㉻y� ���W&����� ?�3�� A��e�/�> �\�3&T�{�� 77߸ ����� ���ݵ ֵ��&��{8 �l1���S�) ���d� *J� F'{s ~��� 6w:0� ��,���s�- Q�v�� ��� ��,�T �ZBLnx6���6 ��6w���Par ���s>�E��j�6d;sq��F  ����8���ЁDhel���x��ti-S�0� �Ob��Dbcf�OX�����t OFT��P<A�_�V�ZI� �D��V\�qWS��=� dtle�Ean�(bzd��tit)v�Z�z�Ez XWO H6�6����5 H�6H691b�E4܀TofkstF\� Y682�4�`n�f804�E91�g�`30oBkmon_��E��eݱ�� ql]m��0 J�fh��}B�_  ZDTf�L0�f(P7�Ec�klKV� �6|��D8q5��ّ�m\b��p��xo�k�ktq���g2.g���yLbmkLVts��IF��bk������Id #I/f��GR� �han�L��Vy��%��%ere������io�� ac�-� A�n�h���c�uACl�_�^ir���)�g��	.�@�& yG��R630�� �p v�p�&H�f��3un��R57v�O�JavG�`Y��o;wc��-ASF��`O��7���SM������
af��rSafLa�vl�\F c�w a���?V�XpoV �30��NT; "L�FFM��=�@���yh	a�G-�w�� �m2.�,�t�<�̹�6ԯ��sd_�MC'V����qD���fslm��isc.  ?H5522���21&dc.pGR78����0��708J61�4Vip A�TUu�@�OL�54]5ҴINTL�6�t�8 (VCA����sseCcRI��ȑ��UI��n�rt\rL�28gn��NRE��.f,��63!��,�SCH��d Ek�DOCV����p��C,�<�L�0�Q�isp��EIO��xE,�54���ѽ9��2\sl,�S�ET���lр�lt�2�J7�Ռ�MASK��̀OPRXY҇��7��n�OCO��J6l��3�l�� (SV�l�A�H�L�@Օ��5�39Rsv���#�1��LCH���OwPLGf�outl�q0��D��HCR
svg��S@�h��cCSa�!�{�50���D�l�5!�lQ��DS�W��S����̀��OiP����7��PR����L�ұ�(Sgd����PCM���R-0 \s��5P՝��0���n�q� A�J�1��N�q�2��P�RSa���69�� �(AuFRDx�Խ��RMCN����93A�ɐC�SNBA�F9� HLB��� M��4����h�2A�95z�H�TCaԈ�TMIL�6�j95,��85�7.,PA1�it�o��TPTXҴ �JK�TEL��pi�L�� XpL�80�I�)��.�!��P;�J9=5��s "N����H�UEC��7\c�s�FR��<Q��C��57\{VCOXa�,���IP1jH��SUI�	CSX|1�AWEBa���HTTa�8�R6%2��m`��GP%��IG %tutKIgPGSj�| RC1w_me�H76��:7P�ws_+�?�x�R51�\iw0�N���H�53!���wL�8!�h�R66 ��H���Ԡ���@;J56��1���N0���9�j��L���RQ5`%�A|�5q�r�`b,�8 5��{165!�d�@�"5��H84!�C29��0��PJ����n B[�J77!Ԩ�R6�5h3n���2y36P��3R6��-`�;о Ԩ@��ex�eKJ87��#J;90!�stu+�~@n!䬵�k90�kop�B����@!�p�@|BA�g*�n@!Ԍ�Q��06!�@[�F��FaP�6��́,�T�S� NC[�CA�B$iͰl1I��R�7��@q�y�CM]S1�rog+QM��� �� TY$x�CTOa�nv\+��1�t(�,�6�con��~0��15��JNN��%e:��P��9OR�S%x���8A�81]5[�FCBaUnZQ��P!��p{��CMOmB��"G��OL���x�OPI�$\lr"[�SŠ�T	D7�U��oCPRQR9RL���S�V�~`���K�ETS�$1��0��p�3�Ԩ�FVR1�LZQV3D$ ���sBVa�SAPL1�7CLN[�PV��	r�CCGaԙ��CL��3CCRA�n �"W!B�H�CSKQn\0�p��)��0CTPn�ЌQe���p!$bCt�aT80U�pCTC�y�:�RC1�1 (�s���trl,�r��
T�X��TCaerrm�r�MC"�s��#wCTE��nrr�R�Ea�XPj�^��r#mc�^�a"�P�Q�F!$���$p "��rG1�tTG$c�8��QH�$SCTI��! s��CTLqdACK�Rp)��r]La�R82��M��0YPk�.���OF��.���e�{�CN���^�1�"M�^�a�С�Q�`US��!$��M�QW��$m�VGF�$R� MH��P2�� H5� ΐq��ΐ�$�(MH[�VP�uo�Y����$)��D��h�g��VPF��"MCHG̑`e!�+�V/vpcm�N��ՙ�N��$�VPRqd)��CV�x�V� "�X��,�1�($TIa�t\�mh��K��etpK�A%Y�VP%ɠ�!�PN���GeneB�rip����<8��extt���Y�m�"�(�� HB���)��x��������Ȣ�reCs.�yA�ɠn� ���*���p�@M�<_�NĀ6L���8�Ș�yAvL�Xr��Ȉ2��"R;�Ƚ\�ra��	P�� h86��Gu+ʸ�Ͽ��SeLɨm�9�69 �P�Ȩr�Ȩ2�ɹ1��n2�h� �0L�XR}�RI{�e� L�x����c�Ș���N�vpx�L��"��2\r� ]�N�82�d���b@�ɉa��y1��/�k�@8���A��ruk�ʘ �L�sop��H�}�t!s{�����s��9���j965��Scx��h��5 J9��{�
�PL�J	ee�n��t I[
x�c�om��Fh�L�4 �J��fo��D�IF+�6�Q����rGati|��p��1�0&�
R8l߾�M�����P��8� �j�mK�X�HZ����IN�oڠ��3�qf��vi���80�~�l Sl�yQ��#tpk�xb�j�.� @�R�d������,/n(�8�8�0���
:�aO8�<�Q}�CO�ں�PT��O (��.��Xp|�~H���?�7v �wv��8��22�pm���722��j7�^�@ƙ�f��cf�=Yvr���vcu���O�O@�O�O_#_5_7�3Y_΋�wv4{_�_w<�ʈ�ust_�_�cus�_�Z��oo�,o>oPo�io��ngqe��(pLy747�j�WelʨHM47ZKEq {���[m�gMFH�?�(wsK� 8J�n���o���fhl;��wmfD���? :�}(4	<�g J{��II)�̏މw��X�774�kﭏ/7ntˏ݊e�+���se�/�aw���8�ɐ��EX \�!b+: �p��~�00��nh�,:Mo+�xO���1 "K�O��\a��#0��.8���{h�pL?�j+�mon�:2��t�/�st�?-�w�:���)�;��(8=h�;
d Pۻ��{:  ��� X�J0��re�����STD�!treLANG��x�81�\tqd��������rch.�������htw�v�WWָ� R�79��"Lo�51 (�I�W�h�՜��4�aww� r�vy �623c�wh a?�cti�֐�!�X�iؠ�t ��n,�։�����j��"AJP�@�3p�vr{�H�6z��!��- SeT�� E3�) G�J93�4��LoW�4 (�S������ <���9c1 ��8!4�j9�搉�+���y�
��	�b]tN�ite{�R  ��I@Ո�����P��������	 ����Z�vol��X ��9�<�I�Lp���ld*���FՇ864{��?��K��	�k扐�֘1�wmsk��M�q�Xa�e�����p��0RBT�1k�s.OPTNЦqf�U$ RTCamT��y��U��y��U��UlU6 L�T�1Tx����SFq�Ue�6T��U�SP W�b DT�qT2h�T�!/�&+��TX�U\j6�&�U U�UsfdO&�&ȁT����662DP�N�bi��%�Q�%62V��$���%�� �#�(�(6To6e St�%��#5y�$�.)5(To�%tT0�%�5�W6T���%�#�#orc��#I���#���%cct�6ؑ?�{4\W6965"p6}"�#\j536��8�4�"�?kruO O�,Im?Np�C �?tx�0<O�;�e �%����?
;gcJ7 "�AV�?�;avsf`�O__&_8WtpD_DV_0GT�F|_:UcK6�_�_r�O�3e\s��O2^y`O:�mig:xGvgW! m�%��q!�%T�$E A{60�po6��#37N�)5CR5_2E���$0��.�$Ada�Vd���V��?;Tz7�_�e7DD!TF9���#8�`�%���4y�ted� Z@�A}�@�}�04�N�}�}���}�dcH& }����u 6�vp��v1�u1\b�u�$2}���}� R83��u�"}��"}�val!g���Nrh�&��8�J�Y�o�ue��� �j70�v=1��MI=G�uerfa��{�q���E�N�ء��E{YE�ce A�� �񁏯pV�e�A!���2�Յ�Q�%��u1�e�i �@��H�e����J0�� '��b��T��E In�B�  W�|���537g����(KMI�t�Ԇr��ݟ�am���nеvi!g�U -�v J߆�8⹖F���P�y�ac����2���Rɏ jox��2�� djd�<8r}� og\k�0r��g��wmf�wFro/� Eq'�<4"}�3 J8��oni[��ᅩ}���� o� ��ʛ��Im@�R�e��{n�Є��V�o������ w ����裆"POS\����ͯ� menϖ�⑥O�Mo�43��� �(;Coc� An[�t���"e�a\�vp�ֽ.��cflx$�l�e��8�hr�tr�N�T� CF+�x �E/�t	qi�M�ӓx1c��p�f�lx����Z�cx��
0 h�כh8��mo��=� �H���)� (�vSER,���g�0߆0\r�vX�= ��I n� - �ti���H��VC�828b�5��L"�RC��Gn G/���w�P�vy�\v�vm "oƀlϚ�x`��=e�ߠ-�R-3?������v<M [�AX/2�)�.S�rxl�v#�0���h8߷=� RAXB�A�����9�H�GE/Rצ����h߶'"RXk��F�˦;85��2L/�xB�885_�q�Ro�0siA��5\rO�@9�K��v����8���.�n "�v��88��8s�i ?�9 ƀ�/�$�y O�M�S"���&�9R �H74&�`�745��	p��p��ycrI0C�c�hP0� j��-�a%?o��6D950�R7trl��ctlO�APC���j��ui"�L���  �.���^棆!�A�ѪqH��&-^7��� ��6s16C�q�794h����� M�ƔI���99��(���$FEAT_AD�D ?	����Q%P  	�H._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�`�r������� ��������&8 J\n���������TDEM�O fY   WM_� �������/ /%/R/I/[/�//�/ �/�/�/�/�/�/?!? N?E?W?�?{?�?�?�? �?�?�?�?OOJOAO SO�OwO�O�O�O�O�O �O�O__F_=_O_|_ s_�_�_�_�_�_�_�_ ooBo9oKoxooo�o �o�o�o�o�o�o >5Gtk}�� ������:�1� C�p�g�y�������܏ ӏ���	�6�-�?�l� c�u�������؟ϟ� ���2�)�;�h�_�q� ������ԯ˯ݯ��� .�%�7�d�[�m����� ��пǿٿ���*�!� 3�`�W�iϖύϟ��� ��������&��/�\� S�eߒ߉ߛ��߿��� ����"��+�X�O�a� ������������� ��'�T�K�]����� ������������ #PGY�}�� ����L CU�y���� ��/	//H/?/Q/ ~/u/�/�/�/�/�/�/ ???D?;?M?z?q? �?�?�?�?�?�?
OO O@O7OIOvOmOO�O �O�O�O�O_�O_<_ 3_E_r_i_{_�_�_�_ �_�_o�_o8o/oAo noeowo�o�o�o�o�o �o�o4+=ja s������� �0�'�9�f�]�o��� ������ɏ�����,� #�5�b�Y�k������� ��ş����(��1� ^�U�g����������� ����$��-�Z�Q� c������������� � ��)�V�M�_ό� �ϕϯϹ�������� �%�R�I�[߈�ߑ� �ߵ���������!� N�E�W��{���� ���������J�A� S���w����������� ��F=O| s������ B9Kxo� �����/�/ >/5/G/t/k/}/�/�/ �/�/�/?�/?:?1? C?p?g?y?�?�?�?�? �? O�?	O6O-O?OlO cOuO�O�O�O�O�O�O �O_2_)_;_h___q_ �_�_�_�_�_�_�_o .o%o7odo[omo�o�o �o�o�o�o�o�o*! 3`Wi���� ����&��/�\� S�e����������� ���"��+�X�O�a� {����������ߟ� ��'�T�K�]�w��� �������ۯ��� #�P�G�Y�s�}����� ���׿����L� C�U�o�yϦϝϯ��� �����	��H�?�Q� k�uߢߙ߫������� ���D�;�M�g�q� ����������
�� �@�7�I�c�m����� ����������< 3E_i���� ���8/A [e������ ��/4/+/=/W/a/ �/�/�/�/�/�/�/�/ ?0?'?9?S?]?�?�? �?�?�?�?�?�?�?,O #O5OOOYO�O}O�O�O �O�O�O�O�O(__1_ K_U_�_y_�_�_�_�_ �_�_�_$oo-oGoQo ~ouo�o�o�o�o�o�o �o )CMzq �������� �%�?�I�v�m���� �����ُ���;�  2�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ������������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ��������'9   :>Ugy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/� A�S�e�w��������� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/
=C6Yk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ������/�A��$FEAT�_DEMOIN [ E��q��>�}Y�INDEXf��u��Y�ILEC�OMP g�;����t�T����SETUP2 �h������  N ܑ��_A�P2BCK 1i~��  �)B�D��%�C�>��� 1�n�E����)���M� ˯�������<�N�ݯ r������7�̿[�� ϑ�&ϵ�J�ٿWπ� Ϥ�3�����i��ύ� "�4���X���|ߎ�� ��A���e�����0� ��T�f��ߊ����� O���s�����>��� b���o���'���K��� ������:L��p ����5�Y�} �$�H�l~ �1��g�� / 2/�V/�z/	/�/�/ ?/�/c/�/
?�/.?�/ R?d?�/�??�?�?M? �?q?O�?O<O����P� 2�*�.VRCO�O�0*��O�O�3�O�O�5w@P�C�O_�0FR6�:�O=^�Oa_�KT ���_�_&U�_�\h�R_<�_�6*.FzOo"�1	(SoEl�_io�[STM �b�o�^�+P�o�m�0iP�endant POanel�o�[H�o� �g�oYor�ZGIF|��e�Oa��ZJPG �*��e`���z��JJS��ĭ��0@���X�%
�JavaScri3ptُ�CSʏ1���f�ۏ %Ca�scading �Style Sh�eets]��0
A�RGNAME.D)T���<�`\��^����Д៍�АDISP*ן���`$�d���V�e��CLL�B.ZI��=�/`:�\��\�����C?ollabo鯕�	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V����zό�!ߘ�TPEI?NS.XML(�@��:\<����Cus�tom Tool�bar}��PAS�SWORD���>�FRS:\��� �%Passwo�rd Config��?J���C��"O ��3�����i����"� 4���X���|����� A���e�����0�� Tf�����O �s��>�b �[�'�K�� �/�:/L/�p/� �/#/5/�/Y/�/}/�/ $?�/H?�/l?~??�? 1?�?�?g?�?�? O�? �?VO�?zO	OsO�O?O �OcO�O
_�O._�OR_ d_�O�__�_;_M_�_ q_o�_�_<o�_`o�_ �o�o%o�oIo�o�oo �o8�o�on�o� !��W�{�"� �F��j�|����/� ďS�e��������� T��x������=�ҟ a������,���P�ߟ 񟆯���9����o� ���(�:�ɯ^��� ��#���G�ܿk�}�� ��6�ſ/�l������ ����U���y�� ߯� D���h���	ߞ�-����Q߻��߇��,��$�FILE_DGB�CK 1i������� ( �)
SU�MMARY.DG<,���MD:`�����Diag Summary�����
CONSLO�G��y����$����Console �log%���	TPOACCN��%g������TP AccountinF����FR6:IP�KDMP.ZIP�����
��)����E�xception�-����MEMCH�ECK������8�Memory �Data��L�N�)�RIPE����0�%�� Packets LE���$Sn�STAT*#�� %LS�tatus�i	FTP�/�/��:�mment �TBD=/� >�)ETHERN�E�/o�/�/��?EthernU<�?figuraL��~'!DCSVRF1/�/)/B?�0 v�erify alylE?�M(5DIFF:? ?2?�?<F\8diff�?}7|o0CHGD1�?8�?�?LO �?sO~3&�
I2BO)O;O��O bO�O�OG�D3�O�O�OT_ ��O{_
VUPDATES.�P�_��?FRS:\�_�]���Update?s List�_���PSRBWLD.CMo���Ro�_�9�PS_ROBO�WEL^/�/:GI�G��o>_�o�G�igE ��nos�ticW�N�>��)�aHADO�W�o�o�ob�S�hadow Ch�ange��{8+"rNOTI?�=O��Not�ific�"��O��A�PMIO �o��h��f/��o�^7U�*�UI3�E��W��{�UI���� ��B���f��_����� ��O���������>� P�ߟt������9�ί ]�򯁯�(���L�ۯ p������5�ʿܿk�  Ϗ�$�6�ſZ��~� �wϴ�C���g���� ��2���V�h��ό�� ����Q���u�
��� @���d��߈��)�� M���������<�N� ��r����%�����[� ���&��J��n ��3��i� �"�X�| ��A�e�/� 0/�T/f/��//�/�=/�/�/�$�$FI�LE_�PPR�P���� �����(MDON�LY 1i5�  
 �z/Q?�/ u?�/�?�?t/�?^?�? O�?)O�?MO_O�?�O O�O�OHO�OlO_�O _7_�O[_�O_�_ _ �_D_�_�_z_o�_3o Eo�_io�_�oo�o�o Ro�ovo�oA�o ew�*��`�����&�O��*VISBCK,81;3*.VDV�����FR:\o�ION\DATA\���/��Visi�on VD filȅ��&�<�J� 4�n������3�ȟW� �����"���F�՟� |������m�֯e��� ���0���T��x��� ���=�ҿa�s�ϗ� ,�>���b���ϗ� ��K���o��ߥ�:����^����ϔ��*MR�2_GRP 1j�;�C4  ;B�}�	 71�������E�� E��  F@ F��5U������L����M��Jk��Lzp�JP���Fg�f�?ǀ  S����9��Y9}�9���8j
�6̿�6�;��Ag�  ���BH��[B���B���$�������������@UUU#�����Y� D�}�h����������������
C��_C�FG k;T �M���]�N�O :
F�0� � \�RM_�CHKTYP  �0�}�000���OM_MIN�	x���50]X� SSBdl5:0��bx��Y���%TP_D�EF_OW0x�|9�IRCOM���$GENOV_RD_DO*62n�THR* d%�d�_ENB� ��RAVC��mK�� ��՚�/�3�/��/�/�� [�M!OUW s�܋}��ؾ��8�g�;?�/7?Y?�[?  C��0�����(7�?�<B�?B�����2��*9�N SMTT#t[)��X�4�$HOSTCd{1ux���?k 	zHzKzO2x��O�Ie�O�O 	__-_;Z�O^_p_�_�_�O�_KP	ano?nymous�_�_�_oo1o yO�O�O zo�_�OM_�o�o�o�o ?_.@Rd�o�_ �_�����;oMo _oqos`��o������ ��̏����&�8� [�����������ȟ �!�3��G�4�{�X� j�|���Տ��į֯� ����e�B�T�f�x� ��џ����	��=� �,�>�P�bϩ��Ϙ� �ϼ����'�9��(� :�L�^ߥ���ɿw��� ����� ��$�6��� Z�l�~��ߴ����� ����� �g�yߋߝ� z����߰��������� ?�.@Rd���� ������;�M� _�q�s`����� ���//&/I 7/�n/�/�/�/�/#O~\AENT 1v
;� P!J/?  ��/3?"?W?? {?>?�?b?�?�?�?�? �?O�?AOOeO(O�O LO^O�O�O�O�O_�O +_�O _a_$_�_H_�_ l_�_�_�_o�_'o�_ Koooo2o{oVo�o�o �o�o�o�o5�oY .�R�v��zQUICC0���3��t14��"�����t2��`�r�ӏ!ROUTERԏ���#�!PCJ�OG$���!1�92.168.0�.10��sCAMgPRTt�P�!d�11m�����RT폟������$NAME �!�*!ROB�O���S_CFG� 1u�) ��Auto-started/FTP&��= ?/֯s����0�B� �f�x���������S� �����,������ ���ϼ�ޯ�������� �ʿ'�9�K�]�oߒ� ߥ߷��������� (:~�k�Ϗ�� �����������1� C�f���y��������� ���,�>�R�?�� cu��`���� �(�$M_q ������ / H%/7/I/[/m/4�/ �/�/�/�/�~/?!? 3?E?W?i?����? �/�?/�?OO/O�/ �?eOwO�O�O�?�ORO �O�O__+_r?�?�? �?�O|_�?�_�_�_�_ o�O'o9oKo]ooo�_ o�o�o�o�o�o�oF_ X_j_~ok�_�� ����o���1� TU��y����������U�)�_ERR �w3�я�PDUS_IZ  g�^�p����>�WRD� ?r�Cq� � guestb�Q�c�u��������"�SCDMNGR�P 2xr����Cqg�\�b��K� 	P01�.00 8(q /  �5p�5pz��5pB  ��{ ���H�W��L��L��L�����O8�����Xl�����a4� x���Ȥ�x��8����\���)�`�;F�������d��.�@�R�ɛ_GROUUېy������	ӑ���QUPD'  ?u����İ�TYg����T�TP_AUTH �1z�� <!iPendan���-�l���!K?AREL:*-�6�H�KC]�m��U��VISION SET���ϴ�g�G� U������R�0��H� Bߏ�f�x��ߜ߮���CTRL {�����g�
S�F�FF9E3��At�FRS:DEFA�ULT;�FA�NUC Web ?Server;�)� ���9�K��ܭ����������߄WR_C�ONFIG |�ߛ ;��ID�L_CPU_PC�Z�g�B�Dpy� ;BH_�MINj�)�~}�GNR_IO���g���a�NPT_�SIM_D_������STAL_SC�RN�� ���TPMODNTOL������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMASTE���ɾeSLAVE� ~��c�O_�CFGٱBUO��O@CYCLE�n>T�_ASG s1ߗ+�
 � ���//+/=/O/ a/s/�/�/�/�/��WNUM��
@�IPCH�^RTRY_CNZ���@�������� @kI�+E�z?�E�a�P_MEMB?ERS 2�ߙ�k $���2�����7�?�9a�SDT_ISOLC  �����$J23_�DSM+�3JO�BPROCN��J�OG��1�+��d8�?���+�O�/?
�LQ �O__/_�OS_e_w_�_`�O Hm@��E|#?&BPOSREQO~��KANJI_����a[�MON #����b�yN_go�yo�o�o�o�Y�`3��<� ��e�_ִ��_�L���"?`EYL_OGGINLE��������$LA�NGUAGE ,��<T� {q��LGa2�	�b���zg�xP��  ���g�'��b����>�MC:\�RSCH\00\�<�XpN_DISP �+G�J��O�O�߃LOCp�Dz����AsOGBOOK ������0󑧱����X��� ��Ϗ����a�*��	p�����!��m��!���=p_BU�FF 1�p��2F幟���՟D�� Collab?orativǖ� ��F�=�O�a�s����� ��֯ͯ߯���B��9�K���DCS }�z� =���'� f��?ɿۿ���H@{��IO 1�� ~?9ü��9�I�[� mρϑϣϵ������� ���!�3�E�Y�i�{߀�ߡ߱��������E��TMNd�_B�T� f�x���������� ����,�>�P�b�t��������L��SEVtD0��TYPN�1�$6���QR�S"0&��<2FL 31�"�J0���������GT�P:pOF�NG�NAM1D�mr�tUPS�GI"5�aO5}�_LOADN@�G %�%O�LPTE^��*MAXUALRM�'p���(��_PR"4�F0d��1�B_P{NP� V 2�C�	MDR07�71ߕ�BL"8�063%�@ ��_#?�ߒ|/�C�A�z�6��/���/Po@�P 2��+ ��ɖ	T 	t  ��/�%W?B? {?�k?�?g?�?�?�? O�?*OONO`OCO�O oO�O�O�O�O�O_�O &_8__\_G_�_�_u_ �_�_�_�_�_o�_4o oXojoMo�oyo�o�o �o�o�o�o0B% fQ�u���� ����>�)�b�M� ����{��������Տ ��:�%�^�p�S��������D_LDX�DISApB�M�EMO_APjE� ?C
  �,�(�:�L�^�p�������ISC 1�C ����4��������4��X���C�_MSTR ����w�SCD 1���L�ƿH��տ� ��2��/�h�Sό�w� �ϛ��Ͽ���
���.� �R�=�v�aߚ߅ߗ� �߻�������<�'� L�r�]������� �������8�#�\�G� ��k������������� ��"F1jUg ������� B-fQ�u����h�MKCFG� ����/�#LT�ARM_��7"0�0N/V$� �METPUᐒ3�ퟎ�ND� ADC�OLp%� {.CMN�T�/ �%� ����.E#>!�/4�%_POSCF�'�.�PRPM�/9ST�� 1��� 4@��<#�
1�5 �?�7{?�?�?�?�?�? �?)OOO_OAOSO�O wO�O�O�O�O_�A�!�SING_CHK�  �/$MODAQ,#����.;U�DEV 	��	�MC:o\HSI�ZEᝢ��;UTA�SK %��%$�12345678�9 �_�U9WTRI�G 1���l3%% ��9o��"ocoFo5#�V�YP�QNe��:SE�M_INF 1��3' `�)AT&FV0�E0po�m)�aE�0V1&A3&B�1&D2&S0&�C1S0=�m)GATZ�o;"tH? g�a[o�xA�� z���� �o>� �o'��K��� ����я:�L�3� p�#�5���Y�k�}�� ����$�[�H���~� 9�����Ưد������ ��ӟ�V�	�z����� ��c�Կ����
��.� ��d��)�;��Ͼ� q�������˿<��� `�G߄ߖ�IϺ�m�� �ϣ����8�J��n� !ߒ�M�������h_�NITOR� G �?�[   	�EXEC1�/�2*5�35�45�55��P�7�75�85�9� 0�Қ�4��@��L� ��X��d��p��|�������2��2���2��2��2��2���2��2��22*3��3��3@�;Q�R_GRP_SVw 1��k (�A�3�3:5E}��3�����ܴ �{j]�Q_�D��^�PL_N�AME !3%�,�!Defa�ult Pers�onality �(from FD�) �RR2� �1�L6(L�?�,0	l d �������� //(/:/L/^/p/�/��/�/�/�/�/�/ZX2 u?0?B?T?f?x?�?�?�?�?\R<?�?�? O O2ODOVOhOzO�O��O�OZZ`\RD�?�N
�O_\TP�O :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo _)_~o�o�o�o�o�o �o�o 2DVh z�[omo���� 
��.�@�R�d�v����������Џ� �Ef  Fb� �F7���   ��!��d��@� R�6�t������l�๟ʝ�����  ݘ����"�@�F�d����� "𩯹�ݐAG�  ϩU[�$�n�B�E� �� � @oD�  �?��� �?�@��A@�;�f��FH� ;�	}l,�	 |���j�s�d�>�� ��� K(���Kd$2K ���J7w�KY/J˷�ϜJ�	�xܿ�� @I���_f�@�z���f�γ�N�������	Xl��������S��ĽÔ��X������5���  �����A?oi#��;���� � �l� �Ϫ�-����ܛG�G�Ѳ���@n�@a   �  ���ܟ*�͵	'� �� H�I� ��  �Рn�:��Èl�È=�s�̈́�в@��@�Е����/������̷NP�  '�,���-�@
��@���?=�@�A���B�  C�j�a�Be�Ci���@#�Bи�N� L 2������bbdʷBР��P����0̠�����ADz՟� n�3��C�i�@�R�RиYщ��  �@�w ���  ��?�ff������n� ɠ#ѱy9�G
(���I�(�@uP@~����t�t���>�����;�Cd;���.<߈<�g�<F+<L�������,�d�,�̠�?fff?��?&�&��@��@x���@�N�@�?��@T�H�� ��!-�ȹ�|�� 
`�������/ /</'/`/r/]/�/��eF���/�/�/�/@m?��/J?�(E���G�#�� F Y�T?�?P?�?�?�?�? �?O�?/OO?OeOk� �O�IQOG�?�O1?��OmO_0_B_T_������A_�_	_�_P�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�ol�o���W�����o;C�E� q�H�d��؜a@q��e��F�BµWB]��NB2�(A����@�u\?��D�������b�0��|�uR�����
x~�ؽ���Bu*C���$�)`�$ ����GC#����rAU�����1�eG��D�I�mH��� I:�I��6[F���C��I��J�:�\IT�H
~�QF�y��p���*J�/ I8�Y�I��KFjʻCe�o��s��� ��Џ���ߏ�*�� N�9�r�]��������� ���۟���8�#�\� G�����}�����گů ���"���X�C�|� g�����Ŀ������ �	�B�-�f�Qϊ�u� ���ϫ��������,� �P�b�M߆�qߪߕ� �߹�������(��L� 7�p�[����������s(4��3:�����$���3���d�,�4��x@�R�wa����l�<~�wa���e����wa4 �{����@��(L:ueP�	P~�A�O�������	���� G2W}h� �����/�� �O�O7/m/[(d=�s/ U/�/�/�/�/�/?�/�1??U?C?y?�=  �2 Ef9gFb-��77�9fB)aa�)`C9A`�&`w`@ -o�?9de�O-OOQOpn�?�?�O�O�O�O�9c?�0�A7ht4Rw`w`!w`xn
 �O9_K_]_o_ �_�_�_�_�_�_�_�_po#ozzQ ��h���G���$MR�_CABLE 2}�h �a:�T� @@�0�A�e��a�a�a��`���0�`C�`�aO8�CtB�m�m�o�f�#���0��0�DO����al?��o�h8�  ���C�07�d4
.�d��`�`�aC�p�bHCE�hm�gҠ`��0�q�p�b0��B���,����5C����y��c -���H� �2���V��� ��������'�"��� D������o<�\ ��������������w*,�** \c�OM �ii����ŋ��%�% 234567O8901i�{� f�H����������1�����
��`��not sent� 5���;��TESTFECS�ALGR  eg�`��1d.�š
:�� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.xsml��ֿ  Z��DEFAU�LT�mi4\bGRPw 2�M�  =���7�E  �%F�orce�sor� check  �����z��p����h5-��ϻ���������%!1st c�leaning �of cont.� v�ilatiCon��}�Rߗ+��@[�ߔߦ߸����mech�cal,`������0��h5k�@�R�d�v������(�rolle _Ƶ����/����(�:�L��Ba�sic quarterly��������,����������F�M��:(�"GpBP(�X_h5��@�����#C���M"��{Pb�t���Sup�pq�grease���?/&/�8/J/\/��C+ ge���. batn�y`/��/h5	/�/�/��/? ?_�ѷenB'�v��/�/��/����?�?�?�?�?�GX=?O(�Dp"CrB1O��0�/`OrO�O�O`�O�t$��Lf��C!-(��A�O:�OO$_�6_H_Z_l_�t*cgabl�O(���S!<(��Q�_:�
_�_ �_oo0oo)(Ӂ/�_�_���_�o�o�o�o��o�O@haul1�l�2r x(�<qC:��op�������Repla�W�fUȼ2�:�.�_4�F�X�j�|�(�$ %���ߟ����#���
� �.�@���d���ŏ׏ ����П����U�*� y�����r��������� 	�q��?�߯c�8�J� \�n���ϯ�����ڿ )����"�4�Fϕ�j� ��˿����������� �[�0�ϑ�fߵϊ� �߮�����!���E�W� ,�{�P�b�t����� ������A��(�:� L�^���������� ���� $s�H�� ����q����� 9]o�Vhz ���U�#�G /./@/R/d/��/�/ ��//�/�/??*? y/N?�/�/�?�/�?�? �?�?�???Oc?u?JO �?nO�O�O�O�O+Jkb	 H�O�O__6M 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<ND@� �bA?�  @!Q _����Fw�� �H;* �** @A>F �pRT�f�x�:�������ҏ��eO^C7� Տ#�5�G�	�k�}��� ُ���c�����W� �C�U�g���ß)��� ��ӯ���	��-�w� ����9�������m�Ͽ���=�O�E!Q��$MR_HIST� 2�>EN�� �
 \
B$ 23�45678901P^�f�#��]�9O ���φϸ�O�)�;� ���q߃ߕ�L�^߬� ���ߦ����7�I� � m�$���Z���~��� ���!���E�W��{��2�����h�����:�S�KCFMAP  ]>EQ��r�5�!P����ON�REL  .��3���EXCFENB8
��Q�FNCXJJOG_OVLIM8dN�\� ��KEY8�=�_PAN7�\���RUN�����SFSPDT�YPxC��SIG�N8JT1MOT��G��_CE_�GRP 1�>EV��@���� �/Ⱥ��/�/ U//y/0/n/�/f/�/ �/�/	?�/???�/c? ?\?�?P?�?�?�?�?��?O)OOMO,���Q?Z_EDIT5 �)TCOM_CF/G 1���[�O�O�O 
�ASI �y3�
__B+[_O_��>O��_bHT_ARC_�U.Ń	T_MN�_MODE5���	UAP_CPL��_gNOCHEC�K ?�� �� o.o@oRodo vo�o�o�o�o�o�o�o�*!NO_WAIT_L4~GiNT�A���EUw�T_ERRs2���3��ƱJ���b��>_)��|MO�se��}x:O��´4�?8�?������ �~�rPARAuM�r������j���5�5�G� = ��d�v�~�X����� �������֟�0����b�t�����S�UM_RSPAC�E�����Aѯۤ�$?ODRDSP�S7�cOFFSET_�CARt@�_�DI�S��PEN_FILE:�7�AF��PTION_IO���q�M_PRGw %��%$*�����M�WORK ��yf ���춍���   � ������	 ч�����It���RG_DSBL'  ��C�{u���RIENTTOJ7 �C~�A���UT_SIM_EDy���V�?LCT ��}{Bx �٭��_PEX�P�=��RAT�W d�c��UP )���`���e�w�X]ߛߩ��$�2r��L6(L?}���	l d�� ����&�8�J�\�n� �������������@�"�4�F�X���2�� ��������������*�<w�Tfx �������J`[ˣG ���Tz��Pg� �����/"/4/ F/X/j/|/�/�/�/� ��/�/??0?B?T? f?x?�?�?�?�?�?�? �?�/�/,O>OPObOtO �O�O�O�O�O�O�O_�_(_:_��O��y_�]2ӆ��_�^�_ �_�W^]^]��/ooSog��Hgrohozo�o �o�o�o�oF`�#|>`�A�  9y�����OK�1�k_�����<��EA�~nq @D�  �qh����nq?��C��s��q1� ;�	l>��	 |�Q�sy�r�q>��u� �sF`H<zH�~�H3k7G�L�zHpG�99l7�k_B�T��F`C4��k�H���Rt��-�Ae���k������s���  �ሏ����Ee�BVT���dZ>=���ڏ ���q-�Fk�yԵ{FbU�= n�@6�  ����z�Fo��Be	'�� � ��I�� �  �<:p܋=���ڟ���@���B��,���B���g�AgN���  '|���g�V�B��p�BӀ�C׏����@  #��Bu�&����� �bbd�B:p2��>�`m�6p�Z�=Dz?o }�܏������׿�������Ǒ��� f�  O� �M���*�?�ff�_8�J�ܿC 3pϑ�ñ8=  �ϵʖq.·�(= �ŁP���'��s�tL�>���/�;�Cd;���.<߈<��g�<F+<L  ��^oiΚrd@��r�6p?fff?�?�&�п�@��@�x��@�N�@���@T싶� Z���ћtމ�u�߈w 	�x��ti�>�)�b�M� ��q���������� ���:�%�^��������W���S�E�  G��=F�� F k���������1U @yd����� �q��	��{�A���h�����a��ird��A{/w/PJ/5/n/vAG�A���":t�/ C^/�/Z/< ލ?���/�/X1??���W����:g��pE� ~1�?�04�0
1�1@I�Ӏ��BµWB�]�NB2�(A���@�u\?����������b��0�|�uR�Ｃ�
�>������Bu*�C��$�)`���? ���GC�#���rA�U����1��eG���I�m�H�� I:��I�6[F����C4OI��J��:\IT�H
~QF�y�O�l@�*J�/ �I8Y�I��KFjʻC��-?�O �O__>_)_b_M_�_ �_�_�_�_�_�_o�_ (oo%o^oIo�omo�o �o�o�o�o �o$ H3lW�{�� �����2��V� h�S���w�����ԏ�� �����.��R�=�v� a�������П����ߟ ��<�'�`�K�]��� ������ޯɯ��&��8�#�\��3(J���33:a������J��3��c4�����������������ڿ�n����ex��n�4 �{2� 2�r�`ϖτϺϨ��%%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ����� �����3��W�B�{�f�4���������d �A����!��1�3�E� {�i�������������  2 Ef�7�Fb�7��6BX�!�!� C9� �� n�@�/`r������#x���+=�3?, V�8Jv�n�n��n��.
 D�� ���//%/7/I/�[/m//�/�:� ���ֻ�G���$�PARAM_ME�NU ?2���  �DEFPULS�E�+	WAIT�TMOUT�+R�CV? SH�ELL_WRK.�$CUR_STY�L� 4<OPT�JJ?PTB_?Y2C�/?R_DECSN  0�Ű<�?�?�?�?�? OO?O:OLO^O�O�O�O�O�O�!SSREL_ID  .�����EUSE_P�ROG %�*%8�O0_�CCCR0�B���#CW_HOST7 !�*!HT�_�=ZT��O_�Sh_zQ��S�_<[_TIME�
2�FXU� GDE�BUG�@�+�CGI�NP_FLMSK�o5iTRDo5gPG�Ab` %l�tkCyHCo4hTYPE�,� �O�O�o# 0Bkfx��� ������C�>� P�b���������ӏΏ �����(�:�c�^��p�����7eWORD� ?	�+
 	�RSc`n�PNeS��C4�JOv1΃�TE�P�CCOL�է�2��gLP� 3��n��OjT�RACECTL �1�2��! ��� �Қ�q�DT Q��2�Ǡ��D Ȼ ��:�� 3ܠ�ԯ� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� �������������� &8J\n�� ������Щ *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6 Fl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� N�߮���������� �,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�?��?�9�$PGTR�ACELEN  ��1  ����0��6_U�P ����RA@�1����1_CFG �ES�3�1
@�<D�<DVOaG�0uO$BD�EFSPD ��/L�1�0��0H�_CONFIG s�E�3 �0��0d�D��2 ��1�APpDsA�A�0���AIN'@TRL ��/MOA8pEQP�E�E��G�pA<D�AILID(C��/M	bTGRP �1ýI l��1B  ������1A�33FC�� F8� E�� @eN	�A�AsA��Y�Y�A�@� 	� vO�Fg�_ ��8cokB;`baBo�,o>oxobo�o�1>�?��?B/�o�o�~�o =%<��
C@y d��"����<��  Dz@�I� @A0�q� �������ˏ ���ڏ���7�"�4�@m�X���|���Ú)ґ�
V7.10b�eta1HF �@����Aq���Q  �?M� �BܠP�p ��C��&�B�EQA���Q�P�Q��� ß[�m����<CA ��0�b�A��̯ޯ���1!CeQKNOW_�M  lE7FbTSoV ĽJ�B oC_�b�t��������������1�]aSM�SŮ�K ���	NE���ĿK���>ODbb��A �RP����0�Ŗά�bQMR�S��T��iN���d���V]S�T�Q1 1�K
 4MU�i��c�kF K�]�oߠߓߥ߷��� ����2��#�h�G�Y� ��}�������
���(���,�27�I��1G�<t�H��P3^�p�����,�4��������,�5(:,�A6Wi{�,�7����,�8�!�3,�MAD�6 �F,�OVLD  �KD�xO.�PARNUM  �|/�T_SCH� E
9'!G)�3Y%UPD/%�E�/P�_CMP_��0@��0'7E�$ER_CHK�%5H�&�/��+RS���bQ_M�O�+?=5_'?O�__RES_G6��:� I�o�?�?�?�?O�? O7O*O[ONOOrO�O �O�{4]��<�?�O z5���O__|3 #_ B_G_|3V b_�_�_|3 � �_�_�_|3� �_�_�o|3Oo>oCo|2V� 1�:�k1!�@�c?�=2THR_�INRc0i!�o5d޲fMASS�o Z��gMN�o�cMON�_QUEUE ��:�"�j0��t4N�� U1Nv�+DpE�NDFqd?`yEXEo`u� BEnpPAsOPTIOMwm;Dp�PROGRAM %$z%Cp}o(/~BrTASK_I���~OCFG ��$/�K�DATA���T���j12 ,ź�̏ޏ�����&� 8�J�\�n���������ȟ{�INFO�����3t��!�3�E�W� i�{�������ïկ� ����/�A�S�e�w�(����Θ� 4�FlJ�a K_N��T��˶ENBg ڽw1���2��GN�2��ڻ P(O��=���]ϸ�@y���v� �u��uɡdƷ_EDIT� �T�����G�W�ERFL�x�c)�RGADJ Ҷ�/A�  $�?j00���a�Dqձӆ5��?��ʨ�<u�j0�%e�������FӨ�2�R��	HJ;pl�G�b_�>�p�Aod�t$��*�/� **:@�j0�$�@�5Y�T���^��q�߈b~� L��\�n����� ����������4�F� t�j�|����������� ��bLBT� x����:�� $,�Pb�� �/����/~/ (/:/h/^/p/�/�/�/ �/�/�/V? ??@?6? H?�?l?~?�?�?�?.O �?�?OO O�ODOVO �OzO�O_�O�O�O�O �Or__._\_R_d_�_@�_�_�_�_�_�f	g� io�pWo�o{d�o��~o�ozoB�PR�EF �Rږp��p
�IORIT�Y�w[���MPDcSP�q��pwUT6�|���ODUCT3������OG��_TG��8��ʯr�TOENT 1���� (!AF�_INE�p,�7��!tcp7�_��!udN���!�icmv��ޯrX�YK�ض���q)�� ,�����p� �&�	��R�9�v�]� o�����П�����ퟐ*��N�`�*�sK���9}�ߢ���Ư B,�/6쒯���������At�,  �Hp��P�b�t����u��w�HANCE C�R��:�wd��连�2s�9Ks���PORT_NUM��s�p���_CARTREP{p|�Ω�SKSTA�w� d�LGS)��ݶ��tӁpUnothing��������{��TEM�P ޾y��'e���_a_seiban�o\��olߒ�}� �ߡ���������"�� �X�C�|�g����� ���������	�B�-� f�Q���u��������� ����,<bM �q��������(L�VER�SIyp�w} �disable�dWSAVE �߾z	2600/H768S?��!ؿ����/ 	�5(�r)og+^/y�e@{/�/�/�/�/�*�,D/? �p���_�p� 1�Ћ� �����Wh?z?��W*pURGE��B��p}vgu,�WF�0DO�vƲ�vW%��4(��C�WRUP_DE?LAY �\κ5�R_HOT %�Nf�q׿GO�5R_NORMAL&H�r6O<�OZGSEMIjO�O|�O(qQSKIPF3	��W3x=_98_ J_\_]�_�_{_�_�_ �_�_�_�_	o/oAoSo owoeo�o�o�o�o�o �o�o+=aO q������� �'��7�]�K��������)E�$RA{����K/�zĀÁ_PoARAM�A3��Kw @.�@`�6�1�2C<��y���C�6$�BÀB�TIF�4`�RCV�TMOUu�c�]�ÀDCRF3��I� �+Q;X�X�D[mD����1=\�2��+�]��^�ޅ��e���k_-_�yS;�C�d;��.<���<�g�<F+<L���Ѱ��d�u�L�������ϯ ����)�;�M�_����RDIO_TYPE  M=U�k��EFPOS1 1��\�
 x4/� ����+�$/<��$� ��pϩ�D���h��ό� �'������o�
ߓ� .ߤ�Rߌ������� 5���Y���i��*�<� v���r��������� U�@�y����8���\� ����������?��c�����2 1�K ԿX�T�x��3 1�����nY�S4 1�'9K�/�'/>�S5 1����/�/�/�/:/S6 1�Q/c/u/�/-?�?Q?�/S7 1� �/�/
?D?�?�?�?d?S8 1�{?�?�?��?WOBO{O�?SMASK 1L��O�D�GXNO���F&�<^��MOTEZ�Ż4��Q_ǁ�%]pA�݂��PL_RAN�G!Q]�_QOWER� �ŵ�P1VS�M_DRYPRG %ź%"O�_�UTART �^��ZUME_PRO�_�_4o��_EXE�C_ENB  <J�e�GSPD`O`8WhՅjbTDBro�j�RM�o�hINGV�ERSION �Ź#o�)I_�AIRPURhP q�O(�MMT_�@�T�P#_ÀOBOT_ISOLC�N�TV@A'qhuNA�ME�l��o�JOB�_ORD_NUM� ?�X#q�H768  �j1Zc@�r
v�rV�s��rw�?�r?�r��pÀPC_TIM�Eu�a�xÀS23�2>R1�� L�TEACH ?PENDANw�:G�X�!O M�aintenance Consj2�����"��No UseB�׏�������1�C�y�V�N�PO�P@�YQz�cS�CH_L`3�%^ �	ő��?!UD1:럒�=R�@VAIL�q@��Ӏ�J�QSPAC�E1 2�ż ��YRs�i�@Ct�YR�Ԁ'{��8�?��˯����"� ��7�2�c�u�����G� ��߯ѿ򿵿�(�� u�AC�c�u������ ��߿���ϵ��(�� =�_�qσϕ�C߹��� ���߱��$��9�[� m�ߑߣ�Q������� ���� ���	�W�i�{� ���M�������5��� .S�e�w����� I�������* ?as��E� ����/&//;/ ]o������/ 2/�/?"?�/7?Y/k/ }/�/�/O?�/�/�?�?��?O0OOKA���*SYPpM*�8.30261 yB�5/21/201?8 A �WPfG�|�H�_TX`�� !$COMME��$USA�p $ENA�BLEDԀ$I9NN`QpIOR�B�@�RY�E_SIGNi_�`�AP�AIT�C��BWRK�BD<�_�TYP�CRIND�XS�@W�@%VFR�I{�_GRPԀ?$UFRAM�rSR�TOOL\VMYH�OL�A$LENGTH_VTEBT�IRST�T  �$SECLP�XU�FINV_POS��@$MARG�I�A$WAIT��`�ZX2�\�VG2�GG1�AI�@�S�Q�	g�`_WR�BNO_?USE_DI�BuQ/_REQ�BC�C]S�$CUR_TC�QP�R"a^f �GP_STATUS�A @ �A3`�B,Lk�H$zc1�h�P�@���@_�FX� �@E_MLT7_CT�CH_�J�`�CO�@OL�E�CGNQQ$W�@w�b�#tDEADLOC�KuDELAY_�CNT�a3qGt�a�$wf 2 JR1[1$X<�2[2�{3[3$Zwy�q %Y�y�q%V�@�c�@�b�$V�`�RV�UV3�oh>b�@ � 8�d�0arMSKJ�Lg�WaZ�C`NRK�PS�_RATE�0$`���S
`�Q�TAC��GPRD���e�S*���a4�A�0�DG�A� 0�P�flp bquS2ppI�#`
`��P 
�S\` � �A�R_E�NBQ �$�RUNNER_A)XI�<`ALPL�Q�R�U�THICQ$�FLIP7��DTF�EREN��R�IF'_CHSU�IW��%V)�G1����$Př�A�Q�Pݖ_JF��PR_P�	�R�V_DATA�A�  $�ET�IM���$VAL�U$�	�OP_ �  �A � 2 �SC�*�	� �$ITP_!�SQ]PNPsOU}�o�TOTL��o�DSP��JOGsLIb��PE_PKpRc�Of�i��PX]P�TAS�$KEPT_MIR��¤"`�M�b�APq�aE �@�y�q�g@١c�q�;PG�BRK6�x�t��L�I��  ?�pSJ�q�P�ADEz��ܠBSOCz�MO�TNv�DUMMY{16Ӂ$SV�`�DE_OP��SFSPD_OVR
����@LD����OmR��TP8�LE���F������OV��S!F��F����bF�d��ƣ&c)�fQc�LCH�DLY��RECOQV���`��W�PM���gŢ�RO������_\F�?� @v�S ��NVER�@�`OFeS�PC,�CSWDٱ�c�ձ���B����TR�G�š�`E_FD}O��MB_CM}���B��BLQ�¢	�dQ�̄Vza�BUP�dg��G
��AM�`��@`KՊ�e�_M!��d�AMf�Q��T$SCA����DF����HBKd�v���IO�U��I'R��PA ����������p��і�?DVC_DB�S!�@x�Q�!�s�d�9�1A���9�3A��ATIEO�0��͠��US����WaAB��R+c��`tá`DؾA��_A�UXw�SUBCP	UP���S�`����3��жc���3�FLA<�B�HW_Cwp"��Ns&�]sAa��$/UNITS�M�F�ATTRIz�Z��CYCL�CNEC�A���FLTR_�2_FI��TARTUPJp����A���LP������_SCmT*cF_F�F_P����b�FS��+�K�CHA/Q��*�d�RSD��Q����Q�v��_TH�PROr���հEMPJ���G�9T� �Q�DI�@y�RAI�LAC/�bMX�L!Of�xS��ځ����X�����PR#�S`a�pp�C� =	��FUNC���RIN`QQP� fԱRA)]R ��pAƠ��AWAR֓F��BLZaWrAkg�ngDAQ�B�rkLD�र&q�dM�K���TI����j��$�@RIoA_SW��AF��Pñ#��%%�p9r�1��MOIQ���D�F_~P(�PD"L�M-�FA�PHRD]Y�DORG�H; �_QP�s%MULS�E~Pz���*�� J⼺Jײ��FAN?_ALMLVG��!�WRN�%HARD�P��UcO�� K2$SHADOW]��kp�a02��� STOdf�+�_^�w�AU{`�R��eP_SBR �z5���:F�� �3_MPINF?�\�8�4��3REGV/1DG�+cVm �C�C�FL(��?�DA`iP���Z`�� ������Z�	 �P(Q]$�A$Z�Q V�|@�[�
� ���EG��o���kAAR���㌵2�axG��wAXE��ROB���RED��W�QD�_�Mh�SYA��AF��FS�GWRI�P~F&��STR����E�˰E"H�)��D�a\2kP�B6P��=V��Dv�O�TO�1)���AR�YL�tR�v�3���F�I&�ͣ$LINQKb!\��Q�_3S���E��QXYZt2�Z5�VOFF��R�R�R�XxPB���ds�G�cF�I�03g�������_J��'�ɲ�S&q�R0LTV[6���aTB�ja�"�bC���DUt�F7�TUR� !X��e�Q�2XP���gFL�E���x@�`��U9Z8���� 1�	)�K��Mw��F9���劂����ORQj��G;W3���#� Ґd ���uz����1�t'OVE�q_�M��ё ?C�uEC�uKB�v'0�x -�wH��t���&  `��qڠ�B�ё�u�q��wh�ECh����ER��K	�EP����AT�K�6e9e0�W���AXs�'� �v�/�R ����! �� ��P��`��` �3p�Yp�1�p� � �� �� (�� 8� � H�� X�� h�� x�� ������DEBU�$%3�I���RAB���ٱ�sV��� 
d�J、 ��@񘧕�������Q ���a���a��3q��Yq�+$�`%"<�cLAB�0b�u�'�GROh���b<��B_s ��"Tҳ*`�0A�u��u8q�p1}�ANDGp��@�����U��p1�� �р�0�Qθuݸ��PN�T0���SERV9E �Z@ $`EmAV�!�PO�� ����nP!�P@�$!Y@  $>�TRQ�b
=��BG�K�%"2\��� ?_  l��5�ND6ERRVb(�I��qV0`;���TOQ:��7�L�@
�R��e G�%�Q�� <�50F�G ,�`�z�>��RA� 2 �d!�����S� � M��pxU ����O�CuG�  >��COUNT6Q��FZN_CFGF�G 4#��6��TG4@�_�=����(���^VC ���M ��"��$6��q ��F!A E� &��X�@� ������A����A9P��P@HEL�0�ҿ 5b`B�_BAS��RSR�6�CSH����1�Ǌ�2��3��4���5��6��7��8��}�ROO����Pf�PNLEA�cAB)�ܫ ��ACKu�IN2O�T��(B$UR0� =�_PU��!0��OU+�Pd�8j���� V��TPFWD�_KAR��� ��R�E(ĉ P�P�>QUE�:RO�p�`r0P1I� x�j�P�8f��6�QSEM��0t��� A��STYL�3SO j�DIX�&p�����S!_TMC�MANRQ��PE�NDIt$KEY?SWITCH����kHE�`BEA�TM83PE{@LEP��>]��U��F���SpDO_HOeM# O�@�EF�p�PRaB�A#PY�C�� O�!���OV_�M|b<0 IOCM��dFQ^�h�HKYA D�Q�7��	UF2��M���p�c�FORC�3WAR�"�OM|@ � @S�#o0U)SP��@1�2&3&4�E���T�O��L�<��8UNLOv�D4�K$EDU1  {�SY�HDDNF�� M�BLOB�  p�SNP�X_AS�� 0�@�0��81$SI=Z�1$VA{��ſMULTIP-��# A� � $��� /4`�B�S��0�C���&FRIFBO�S���3�� NF�ODBU�P߰�%@3;9(űp��S��Z@ x��S�I��TEs�r�cSKGL�1T�Rp&���3B��@�0STMTdq�3Pg@VBW�p��4SHOW�5@��SV��_G�� 3p$PCJ�PИ���kFB�PHSP 1AW�EP@VD�0WC�� ���A00��PB XG XG �XG$ XG5VI6VI7�VI8VI9VIAVIB�VI�XG�YF�0XGFPVH��XbI1oI1|IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1Y1YU2UI2bI2oI2|I2�I2�I�`�X�I2pT�X�I2�I2�I2�I2�I2Y2Y�p�h�bI3oI3|I3�I3��I3�I3�I3�I3��I3�I3�I3�I3��I3Y3Y4�i4�bI4oI4|I4�I4��I4�I4�I4�I4��I4�I4�I4�I4��I4Y4Y5�i5�bI5oI5|I5�I5��I5�I5�I5�I5��I5�I5�I5�I5��I5Y5Y6�i6�bI6oI6|I6�I6��I6�I6�I6�I6��I6�I6�I6�I6��I6Y6Y7�i7�bI7oI7|I7�I7��I7�I7�I7�I7��I7�I7�I7�I7��I7Y7T[�V5P� UD�y"ՠ���
<A62��:t�R��CMD� ���M5�Rv�]��Q_h�R���e����<��YSL���  � �%\2��+4�'�W�BVALU���b��'���FH�IgD_L���HI��9I���LE_���f��$0C�SACѿ! h �V?E_BLCK���|�1%�D_CPU5� � 5ɛ �����C�� ���R " � �PWj��#0��LA�1SBћì���RUN_FLG�� �����ĳ ��������B��H���Х�M��TBC2��# � @ B��e �S�p8=�FTDC�����V���3d�Q�T!HF�����R�L�?ESERVE9��F��3�2�E��Н��X -$��LE�N9��F��f�RA���W"G�W_5�b�14��д2�MO-�T%	S60U�Ik�0�ܱF����[�DEk�21LgACEi0�CCS#0�� _MA� j��z��TCV����z�T�������.Bi�'AH�z�'AJh�#EM5�"��J��@@i�V�z���2Q �0&@o�h�6��JK��VK9��0{���щ�J0�����JJ��JJ��AAAL���������4��5�ӕ N1����딨�.�LD�_�1�* �CF�"% `�GROU���1��AN4�C�#m RE�QUIR��EBqU�#��6�$Tk�2$���zя #��& \�APPR� C� 0�
$OP{EN�CLOS"�St��	i�
��&' �MfЩ����W"-_MG�7C�B@�A���BBR=K@NOLD@�0RTMO_5ӆp1J��P�������������60��1�@ )!�>#�(� ������'��+#PATH''@!6#@!�<#� r� '��1SCA�؆�6IN��UChJ�[1� C0@UM�(Y ��#�"�����*����*��� PAYLO�A~J2LؠR_AN^�3L��91��)1AR_F2L3SHg2B4LO4�!�F7�#T7�#ACRL�_�%�0�'�$��H���.�$HA�2FWLEX��J!�) P�2�D߽߫����0��* : ����z�FG]D����z���%�F1]A�E�G�4�F�X�j�|���BE ������������ (��X�T*�A���@�X I�[�m�\At�T$g�QX<�=��2TX���e mX��������������@����+	�J>+ �-�K]o|��٠AT�F�4�ELPFP���s�J� *� ;JEmCTR�!�A�TN�vzHAN/D_VB.��1��n$, $8`F2Av���SWu	#-� $$M*0 .�]W�lg��PZ����A��� 1�����:AK��]AkA�z��LN�]DkD�zPZ G��C�ST�_K�lK�N}DY ��� A����0��<7 ]A<7W1�'��d�@g`�P��������" 1B$. M�2D%"��H����OASYMj%0�� Bj&-��-W1�/_� {8� �$�����/�/�/�/ 3J<�:9��/�89�D_VI��v����V_UNI�ӛ��cD1J����� ��W<��n5Ŵ�w=4�@�9��?�?<�uc�4��3C�%�H���a/�j��0�DIz�uO��?�k�>S0 �`��I��A� �#���@ģ���@����IPl� 1 � -/�ME.Qp��49�ơT}�PT�;pG �+ Gt� ����'��T�0 $DUMMY1���$PS_�@RF��@  G b�'FLA@ YP(c|��$GLB_TP� ŗ���9 P�q���2 X� z!ST�9�� SBRM M�21_V�T$S/V_ER*0O�p�Ӧ��CL����AGPOl��f�GL~�EW>��3 4H �$Y
rZrW@�x�A1+��A���"	""�U&�4� 8`NZ�"�$�GI�p}$&� �-� �Y�>�5 L�H {��}$F�E^��NEAR(PN�CyF��%PTANC�B�	!JOG�@� �6.@$JOIN�Twa?pd�MSET.>�7  x�E��HQ�tpS{r��up>�8׼ �pU.Q?��� LOCK_FOxV06���BGLV�s�GLt�TEST_sXM� 3�EMP�����_�$U&@%�w`24� Y��5��2�d��3��C�E- ���� $KA�R�QM��TPDRqA)�����VECn@���IU��6��H=Ef�TOOL�C2�V�DRE IS3�ER6��@ACH� 7?Ox �Q��29Z�H I� � @$RAIL_�BOXEwa�R�OBO��?��HOWWAR�1�_�zROLMj��:q�w�jq� �@ O_=Fkp! d�l�>�9�� �R OB8B: �@�c�KOU�;�Һ�3ơ��r�q_�$PIP��N&`H�l�@���#@CORDED�d�p >f�fpO�� �< D ��OB⁴sd���Kӕи��qSYS�A�DR�qf��TCH�t� = ,8`E�No��1Ak�_{��-$Cq,Be�VWVA~��> �  �&��PREV_R�T�$EDIT�r&VSHWRkqP�֑ &R:�v�D���JA�$�a$HECAD�6�� �z#�KE:�E�CPSP]D�&JMP�L~�2�0R*P��?��1�%&I��S�rC�pN�E; �q�wTICK��C��M�1<�3H=N��@ @� 1Gu�!_GPp6��0gSTY'"xLO���:�2l2?�A t 5
m G3%%$R!{�u=��S�`!$�� w`���ճ���Pˠp6�SQU��E��u�T�ERC�Q2�TSUtB ����hw &`gw�Q)�pO���F�@IZ��{��^уPR�kюB1XP9U���E_DO��, �XS�K~�AXI4�@���UR�pGS@�r� ^0�&��p_) �ET�BPm��o�%�0Fo��0A|���CRԍ��a;�{SR�Cl>@ P��b_�yUr��Y��yU ��yS��yS���UЇ�U ���U���U�]��Ul [��Y�bXk�]Cm鯰����YRSC�� oD h�DS~0̕�Q�SP���eAT�ހ���A]0,2N�A_DDRES<B} �SHIF{s��_2+CH�p�I��=qW�TVsrI��E"P���a�CT�
��
;�qVW�A��F \�Ђq��0l|\A@�rC��_B"R{zp�ҩq�TXSCREE��Gv��1TINA���t{����A�b?�H T1�ЂB� ����I��A��BE�y RRO������ B���D��UE4I ��g�!p�S��RSyM]0�GUNEX(@~Ƴ�j�S_S�ӆ�� Á։񇣣�ACY��0� 2H�pUE�;�J�����@GM�T��Lֱ�A��O^	�BBL_| W8�N��K ��0s�OM��LE/r��� TyO!�s�RIGH���BRD
�%qCKG9R8л�TEX�@��>��WIDTH�� ��B[�|�<��I_���Hi� L 8�K���_�!=r���R�:�_��Yґ��O�6q�Mg0紐U䟐h�Rm��LUM8h��FpERVw��P���`�N��^&�GEUR��FP�)�)� LP��(RE%@�a)ק�a�!��Tf �5�6�7�8Ǣ#B�É@���tP�jfW�S@M��USR&�O <�����U�Qs�FO�C)��PRI;Qmx� :���TRIP��m�UN����Pv��0��f%��'���@�0 Q����AG �0T� �a>q&�OS�%�RPo���8�R/�A�H�L�H�4����U¡�SU��g��¢5��OFFT���T�}�O��� 1R�����SN�GUN��6�B_SUB?���,�'SRTN�`TUg2���mCOR| D�RA�UrPE�TZ�#'�VsCC��	3V AC36MFB1f$�c�PG �W (\#��ASTEM������0PE��T3G��X �\ ��MOcVEz�<���AN��� ���M���LIM_X��2��2��7�,�����ı�
��V�F�`E���~��04Y���IB�7���5S���_Rp� 2��� WİGp+@���}СP��3�Zx ���3���A�ݠCZ�DRID����Vy08�90� �De�MY_UBY�d���6��@��!8��X��P_S��3ڶ�L�KBM,�$n+0DEY(#EX`�|����UM_MU� 1X����ȀUS�� ����G0`PACI ���а@��:��:,�:����RE/�3qL�F+C��:[��/TARG��P�r ����R<�\ d�`��A��$�	��ARF��SW2 ��-���@Oz�%qA7p�yREEU�U�01�,�+HK�2]g0�0qP� N� �EAM0G�WOR���MR�CV3�^ ���O*�0M�C�s	���|�REF_��� x(�+T� ����������3_RC H4(a�P�І�hrj�pNA�5��0�_ ��2�����L@��n�@@OAU~7w6���Z�6�a2[��RE�p�@F;0\�c�a'2K�@WSUL��]��C��f0�^��� NT�� L�3��(6I�(6q�(3� L��Q5��Q5I�]7Jq�}�Tg`4D`�0�.`0�AP_HU�C�5SA��CMPBz�F�6�5�5�0_�aAR��a�1I\!X�9��GFS��ad� ��M��0p�U�F_x��B� �ʼ,R�O��Q��'����URF�3GR�`.�3IDp���)�D�;��A,��~�IN��H{D���V@AJ���S͓UWmi=�����TY&LO*�5���󾖄bt +�cP�A� �cCACH�vR�UvQ��Y���p�#CF�I0sFR��XT���Vn+$HO����P!A3�XB�f�(1 ���$�`VPxy� ^b_SZ3132he6K3he12J�eh� chG�chWA�UM�P�j��IMG9�uPAD�iiIMRyE�$�b_SIZ�$�P����0 ��ASY�NBUF��VRT�D)u5tqΓOLE�_2DJ�Qu5R��C���U��vPQuEwCCUlVEMV x�U�r�WVIRC�aIuVTPG���rv01s��5qMPLAqa�R�v�V0�cm� _CKLAS�	�Q�"��d  �ѧ%ӑӠ@}¾�$�Q���Ue |�0!�rSr��T�#0! �r�iI���m�vK�BG��VE�Z�PK= �v�Q��&�_HO�0��f � >֦3�@Sp��SLOW>�R=O��ACCE���!� 9�VR�#���p:����AD�����PA�V�j�� D����M�_B"���^�JMP�G ��g:�#E$SSC��x&�vPq��IhݲvQS�`qVN���LEXc�i T�`�sӂ��Q�FLmD �DEsFI��3�02���:��VP}2�Vj� �A���V�4[`MV_PIs��t���A�@&��FI��|�Z��Ȥ������A���A��~�G9Aߥ1 LOO��1 JCB���Xc��^`�#PLANE��R��1F�c�����pr�AM� [`�噴��S�� ��f����Af��R�Aw��״tU��pRKE<��d�VANC�A\���� k����ܲϡ�R_AA� Al��2� ��p�# Î��m h�@��O K��$������kЍ0O)U&A�"A�
p�p�SK�TM@FVIEM 2l ��P=���n <<��dK�/UMMYK1P���`D�ȡ�C�U��#AU��o �$��TIT�g$PR����OP���VSHIF�r�p`J�Qs�ؙ�fOxE$� _R�`U�#����s��q ������G�"G�޵'�9T�$�SCO{D7�CNTQ i�l�>a� -�a�;�a�H�a�V����1�+�2u1��D�����  � S�MO�Uq��a�J,Q�����a_�R[�ir�n�*@LIQ��AA/`�XVR��s��n�TL���ZABC�t�t�c�]
L�ZIP��u撖��LVbcLn"�^��MPCFx�v:��$�� ���DMY_LN�������@y�w Ђ(a�u� �MCM�@CbcCA�RT_�DPN� �$J71D ��=NGg0Sg0�B�UXW� ��UXE#UL|ByX����	������x 	���m�Y�H�Db  y 8x0���0EIGH�3Fn�?(� H����$z ���|�����K$B� Kd'��_��,L3�RVS�F`���OVC�2'�$|�>P&��
q���5MD�TR�@ �Vc���SPHX��!{ �,� *<�$R��B2 2 ����C!�  ���V+L�Hb*c%g!`+g"�`�V*�,8�?�V+�/V.�/�/?�/�/V(7%3@/R/d/v/ �/6?�/�/�?�?�?O4OOION;4]?o?�? �?�?SO�?�?�O_�O 0_Q_8_f_N;5zO�O �O�O�Op_�O_o8o@�_MonoUo�oN;6�_ �_�_�_�_�oo%o4�Uj�r�N;7 �o�o�o�o�o� B Q�r�5���������N;8�����Ǐ=� _�n���R���ş��ڟ�N;G �) џ�
����?� ��W�i�{�������ï �.�������A��dW�<�N�|����� ��Ŀֿ�ޯ��� 0�B�_�R�d�꿤϶� ������������*� L�^��rτ�
����� �������&�8�J��l�~� `ҟ @�з����ߩ��-����&�,��� 9�{�����a������� ��������A' Y����������a#1�
���N;_MODE�  ��S E��[�Y�B���
/\/*	|/�/R4�CWORK_AD��
<wdT1R  ���� �/� _INTVAL��+$��R_OPT�ION6 ��q@V_DATA_?GRP 27���D��P�/~?�/�? �9��?�?�?�?OO ;O)OKOMO_O�O�O�O �O�O�O_�O_7_%_ [_I__m_�_�_�_�_ �_�_�_!ooEo3oio Woyo�o�o�o�o�o�o �o/eS� w������� +��O�=�s�a����� ��͏���ߏ��9��'�I�o�]�����$�SAF_DO_PULS� �~�������CAN_TIM�����ΑR ��������5�;#U! P"�1!��� �?E� W�i�{�����.�ïկ`�����'(~�ET"2F��Q�dF�"a��2�o+@a얿 ����)�u��� k0ϴ���_ ��  T� � �2�D�)�?T D��Q�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ�x/V凷������߽��R�;��o �W�p��
�t��Diz$�� �0 � � T"1!������� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FX ��࿁����� ��/`4�=/O/a/ s/�/�/�/�/�/�/�!!/ �0޲k�ݵu�0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o k$o6oHoZolo~o�o �o�o�o1/�o�o  2DVhz�/5? ��������&� 8�J�\�n��������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c�u��� ���`Ò� ϯ����)�;�M� _�q���������˿ݿ�� ����3� ����&2,��	�12345678�v�h!B!���2�Ch��� 0�ϵ���������� !�3�9ѻ�\�n߀ߒ� �߶����������"� 4�F�X�j�|�h�K߰� ��������
��.�@� R�d�v����������� ���*<N` r������� &��J\n� �������/ "/4/F/X/j/|/;�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�/�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_�?L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o=_ �o�o�o�o�o�o  2DVhz�����h������u��o.�@�R���Cz�  B��   ����2&� �� _�
���  	�_�2�Տ�X���_�p������ďi�{������� ß՟�����/�A� S�e�w���������N� �����+�=�O�a� s���������Ϳ߿�@��'�9�K�_��丁��<v�_��$S�CR_GRP 1�
� ��� �t ���� ��	 /������� ���������_����8��)�a����&�?DE� DW8����l�&�G�CR-�35iA 901�23456789}0��M-20���8��CR35 ���:�
��������������:֦����G���&������	��]�o����:�?��H���>������������&���ݯ:��j�����g������B�t�Ɛ��������A���� c @�`��@� N( ?�=��Ht��P
��F@ F�`z�y���� �� �$H���Gs^p��B��7��/�0/ /-/f/Q/�/u/�/�/ �/8���P�� 7%?�����"?W?-2?;�-"]? H�1�?t�ȭ7�������?-4A, �&E@��<�@G�B-1  3OZOlO-:HA�H�O\�O|O P�B(�B��O�O_��EL_D�EFAULT  ������`SHOTST�R#]A7RMIPO�WERFL  �i�/UYTWFDO�$V /URRVE�NT 1�����NU L!D?UM_EIP_-8��j!AF_I�NE#P�_-4!FIT�_->�_;o!���`o �*o�o!�RPC_MAINĈojh�vo�o�cVI�S�oii��o!�TPpPU�Yd�k!
PMON?_PROXYl�VAeZ�2r��]f���!RDM_S�RV��Yg�O�!#R��k��Xh>���K!
�`M��\i����!RLSYN�C�-98֏3�!�ROS�_-<�4�"��!
CE4pMOTCOM���Vkn��˟!	��CONSd̟�Wl���!���WASRC��Vm��c�!��USBd��XnR���Noӯ� ������!��E��i��0���WRVICE�_KL ?%�[� (%SVCPGRG1��-:Ƶ2ܿD�˰3�	�˰4,�D1�˰5T�Y�˰6|���˰7�ϩ�˰�����9����ȴf�!� ˱οI�˱��q�˱� ��˱F���˱n���˱ ���˱��9�˱��a� ˱߉��7߱��_� �������)�� ��Q����y��'�� �O����w����� ����˰��İ d�뱭���� =(as^� �����/�/ 9/$/]/H/�/l/�/�/ �/�/�/�/�/#??G? 2?k?V?}?�?�?�?�? �?�?O�?1OCO.OgO RO�OvO�O�O�O�O�O�	_�O-_��_DEV� �Y�M{C:5Xd�GTGRP 2SVK ���bx 	� 
 ,�P5_�_�R �_�_�_�_�_�_3oo Wo>o{o�oto�o�o�o �o�o�o/A�_e ������� �� �=�$�6�s�Z� ��~���͏���H� '�ޏK�2�o���h��� ��ɟ۟���#�5� �Y�@�}�d�v���
� ׯ�Я���1��*� g�N���r�������� ̿	���?�&�c�u� ̯��PϽ��϶����� �)��M�4�q�X�j� �ߎ��߲������%� |��[���f��� �����������3�� W�i�P���t������� ��>�A(e L^������ � =O6sZ �� ���/� '//K/]/D/�/h/�/ �/�/�/�/�/�/#?5? ?Y?�N?�?F?�?�? �?�?�?O�?1OCO*O gONO�O�O�O�O�O�O��O�O_kT �"V	 	_R_=_v_a_�_�_�_��[%��_�_�S���a�Qeo)go Io7omo[o�o�i�_�o i�o�o�o%' 9o�o��o_�� ����!�w�n� �G�����ŏ���׏ �O�4�s���g���w� ���������'��K� ՟?�-�c�Q�s����� �����#�����;� )�_�M�o���ׯ���� ���ݿ��7�%�[� ���ϔ�K�m�Gϵ��� �����3�u�Zߙ�#� ��{ߝߟ߱������ M�2�q���e�S��w� ������%�
�I��� =�+�a�O���s����� ���!���9' ]K������q� m��5#Y� ��I����� /�1/sX/�!/�/ y/�/�/�/�/�/	?K/ 0?o/�/c?Q?�?u?�? �?�??�?O�?�?�? )O_OMO�OqO�O�?�O O�O_�O__%_[_ I__�O�_�Oo_�_�_ �_�_oo!oWo�_~o �_Go�o�o�o�o�o�o 	_o�oV�o/�w �����7�[ �O��_���s����� ͏��3���'��K� 9�[���o����̟� �����#��G�5�W� }������m�ׯů�� ���C���j�|�3� U�/���ӿ������ ]�Bρ��u�cυχ� ���Ͻ���5��Y��� M�;�q�_߁߃ߕ��� ���1߻�%��I�7� m�[�}�������	�� ����!��E�3�i��� ����Y���U������� A��h��1� ������[ @	sa��� ���3/W�K/ 9/o/]/�/�/�/��/ �/�/�/�/?G?5?k? Y?�?�/�?�/?�?�? �?�?OCO1OgO�?�O �?WO�O�O�O�O�O�O 	_?_�Of_�O/_�_�_ �_�_�_�_�_G_m_>o }_oqo_o�o�o�o�o �ooCo�o7�oG m[���o� ���3�!�C�i�W� ������}��Տ� ��/��?�e�����ˏ U������џ���+� m�R�d��=������ ��߯ͯ�E�*�i�� ]�K�m�o�������ۿ ��A�˿5�#�Y�G� i�k�}ϳ�����ϣ� ���1��U�C�e߻� �ϲ��ϋ�����	��� -��Q��x��A�� =���������)�k� P������q������� ����C�(g���[ Im����  ?�3!WE{ i������� �///S/A/w/��/ �g/�/�/�/�/�/+? ?O?�/v?�/??�?�? �?�?�?�?�?'Oi?NO �?O�OoO�O�O�O�O �O/OUO&_eO�OY_G_ }_k_�_�_�__�_+_ �_o�_/oUoCoyogo �o�_�oo�o�o�o 	+Q?u�o��o e������'� M��t��=�����ˏ ���ݏ�U�:�L�� %���m�����ǟ��� -��Q�۟E�3�U�W� i�����ï��)��� ��A�/�Q�S�e��� ݯ¿�������� =�+�Mϣ�ɿ��ٿs� �ϻ�������9�{� `ߟ�)ߓ�%ߣ��߷� �����S�8�w��k� Y��}�������+� �O���C�1�g�U��� y��������'��� 	?-cQ���� �w�s�; )_���O�� ���//7/y^/ �'/�//�/�/�/�/ �/?Q/6?u/�/i?W? �?{?�?�?�??=?O M?�?AO/OeOSO�OwO �O�?�OO�O_�O_ =_+_a_O_�_�O�_�O u_�_�_o�_o9o'o ]o�_�o�_Mo�o�o�o �o�o�o5wo\�o %�}����� ="�4����U��� y�����ӏ���9�Ï -��=�?�Q���u��� �ҟ�����)�� 9�;�M���ş���s� ݯ˯��%��5��� ������[�����ٿǿ ���!�c�Hχ��{� ϋϱϟ�������;�  �_���S�A�w�e߇� �ߛ������7���+� �O�=�s�a����� �������'��K� 9�o������_���[� ������#G��n ��7������ �aF�yg ������9/ ]�Q/?/u/c/�/�/ �/�%/�/5/�/)?? M?;?q?_?�?�/�?�/ �?�?�?�?%OOIO7O mO�?�O�?]O�O�O�O �O�O!__E_�Ol_�O 5_�_�_�_�_�_�_�_ o__Do�_owoeo�o �o�o�o�o%o
�o �o�o=sa�����o�!+q�$SE�RV_MAIL � +u!���O�UTPUT��$�@�RV 2��v  $� (�q�}��SAVE�7�	�TOP10 �2W� d  'ݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w����������ѿ�u��YP����FZN_CF�G �u�$�~����GRP� 2�D� ,�B   A[�+qD�;� B\�� � B4~�RB{21��HELL�C�u��j�k�2�|����%RSR�� �����
�C�.�g�R� ��v߈��߬�����	����-�?�Q��  �_�%Q���_����,p����Sޖ�g�2,pd��|���HK 1�� ��E�@�R�d� ���������������� *<e`r�~��OMM ������FTOV_E�NB�_���HOW_REG_UI��	�IMIOFWD�L� �^�)WAIT���$V1�r^�NTIM7���VA�_>)_UNIT��v��LCTRY�B��MB_H�DDN 2W� 2�:%0 �pQ/ �qL/^/�/�/�/�/�/��/�/�"!ON_ALIAS ?e�	f�he�A?S?e? w?�:/?�?�?�?�?�? OO&O8OJO�?nO�O �O�O�OaO�O�O�O_ "_�OF_X_j_|_'_�_ �_�_�_�_�_oo0o BoTo�_xo�o�o�o�o ko�o�o,�oP bt�1���� ���(�:�L�^�	� ��������ʏu�� � �$�Ϗ5�Z�l�~��� ;���Ɵ؟����� � 2�D�V�h�������� ¯ԯ���
��.�ٯ R�d�v�����E���п ���ϱ�*�<�N�`� r�ϖϨϺ���w��� ��&�8���\�n߀� �ߤ�O���������� ��4�F�X�j�|�'�� �����������0� B���f�x�������Y� ��������>P bt����� �(:L�p ����c�� / /$/�H/Z/l/~/)/ �/�/�/�/�/�/? ?�2?D?V?]3�$SM�ON_DEFPR�O ����1 �*SYSTEM*�0m6RECAL�L ?}9 ( �}]?�?�?�?OO)O �?NO`OrO�O �O�O;O�O�O�O__ &_�OJ_\_n_�_�_�_ 7_�_�_�_�_o"o�_ FoXojo|o�o�o3o�o �o�o�o�oBT fx��/��� ����>�P�b�t� ������=�Ώ���� �(���L�^�p����� ��9�ʟܟ� ��$� ��H�Z�l�~�����5� Ưد���� ���D� V�h�z�����1�¿Կ ���
�ϯ�@�R�d��vψϚ�-�5cop�y frs:or�derfil.d�at virt:�\temp\=>�147.87.1�49.40:80�08����)� }-��*.d�������~ߐߢ�5�
xyz�rate 61 �J�\�n����#�6� ���������߁����8�8����mpba�ck��q���)� �}/��mdbG�*������������7�3x��:\H���Z�[�pt�) }4��a����p������ ����W�r�':� �^�������K ]���/#/6�� l}/�/�/��O� �/??2D�/hy? �?�?��U/��?	O O./@/�?d/�?�O�O�,O:�$h:\su�pportIH�I=�>2611609�60:56058�9�O
__�,tp?disc 0_Ou@��O�O_�_�_�%t�pconn 0 �H_Z_l_�_o!o�'=�?6olptest.tp��HgG_uO�o �o�/�/K?koxo	 .?@?�od?�o���~��$SNPX_A�SG 2�����q� �P 0 '%�R[1]@1.Y1��y?��s%� !��E�(�:�{�^��� ����Տ��ʏ��� A�$�e�H�Z���~��� џ����؟�+��5� a�D���h�z�����ů �ԯ���
�K�.�U� ��d�������ۿ��� ���5��*�k�N�u� �τ��ϨϺ������ 1��U�8�Jߋ�nߕ� �ߤ����������%� Q�4�u�X�j���� ���������;��E� q�T���x��������� ��%[>e �t������ !E(:{^� �����/�/ A/$/e/H/Z/�/~/�/ �/�/�/�/�/+??5? a?D?�?h?z?�?�?�? �?�?O�?
OKO.OUO �OdO�O�O�O�O�O�O _�O5__*_k_N_u_ �_�_�_�_�_�_�_o 1ooUo8oJo�ono�o��o�d�tPARAM� �u�q ��	��jP�d�9p�ht��pO�FT_KB_CF�G  �c�u�sO�PIN_SIM  �{vn���p�pRVQSTP/_DSBW~r"t|�HtSR Zy� � & O?LPTEST����vTOP_O�N_ERR  �uCy8�PTN �Zuk�A�4�RING_PR�MB� �`VCNT_GP 2Zu:q�!px 	r���ɍ���׏��wVD>��RP 1�i p�y��K�]�o��� ������ɟ۟���� #�5�G�Y���}����� ��ůׯ�����F� C�U�g�y��������� ӿ��	��-�?�Q� c�uχϙϫ������� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�^�[�m��� �����������$�!� 3�E�W�i�{������� ��������/A Sew����� ��+=Ov s������� //</9/K/]/o/�/ �/�/�/�/�/?�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO)��PRG_COUN��:t�k�GuKBENB��FEMpC:t}O_UPD 1�{T  
4Or�O �O�O__!_3_\_W_ i_{_�_�_�_�_�_�_ �_o4o/oAoSo|owo �o�o�o�o�o�o +TOas�� ������,�'� 9�K�t�o��������� ɏۏ����#�L�G� Y�k���������ܟן ���$��1�C�l�g� y���������ӯ���� 	��D�?�Q�c����� ����ԿϿ�����)�;�d�_�q�=L_I�NFO 1�E��@ �2@����������� ��6���c80ͻ6���W��´ ���<LYSDOEBUGU@�@����d�If�SP_PA�SSUEB?x�L_OG  ���Ce��*ؑ�  V����  UD1�:\�ԘΥ�_MPAC�ݵE&�8�AV��X�A�SAV �!�������X����SVZ�TEM_TIME 1"��]�@ 0��2X�����������$T1?SVGUNS�@VE�'�E��ASK_OPTIONU@�E�A�A+�_DI���qOG�BC2_GRP 2#�I���~��@�  C����<Ko�CFG %�z��� ���`��	�.>dO �s������ �*N9r]� ������/� 8/#/\/n/v$Y,�/ Z/�/�/H/�/?�/'? ?K?]�k?=�@0s?�? �?�?�?�?�?O�?O O)O_OMO�OqO�O�O �O�O�O_�O%__I_ 7_m_[_}__�_�_�X � �_�_oo/o�_So Aoco�owo�o�o�o�o �o�o=+MO a������� ��9�'�]�K���o� ��������ɏ���#� �_;�M�k�}������ ��ß�ן��1��� U�C�y�g��������� ������	�?�-�c� Q�s����������Ͽ ����)�_�Mσ� 9��ϭ�������m�� �#�I�7�m�ߑ�_� �ߣ����������� !�W�E�{�i����� ����������A�/� e�S�u�w��������� ����+=O��s a������� 9']Kmo �������#/ /3/Y/G/}/k/�/�/ �/�/�/�/�/??C? ��[?m?�?�?�?-?�? �?�?	O�?-O?OQOO uOcO�O�O�O�O�O�O �O__;_)___M_�_ q_�_�_�_�_�_o�_ %oo5o7oIoomo�o Y?�o�o�o�o�o3 !CiW��� ������-�/� A�w�e���������� я���=�+�a�O� ��s�������ߟ͟� �o�-�K�]�o�ퟓ������ɯ���צ���$TBCSG_G�RP 2&ץ�  ��� 
 ?�   6�H�2�l�V���z���@ƿ�������(��d�E+�?~�	 HC����>���G����C�  A�.�e�q�wC��>ǳ33��"S�/]϶�Y��=Ȑ� C\  Bȹ���B���>���X�P���B�Y�z�"�L�H�0�$���� J�\�n�����@�Ҿ ���������=�Z�%�07����?3������	V3.0�0.�	cr35��	*����
���0������ 3���4�   {�CaT�v�}��J2��)������CFG� +ץ'� ,*������I����.<
� <bM�q��� ����(L7 p[����� �/�6/!/Z/E/W/ �/{/�/�/�/�/.�H� �/??�/L?7?\?�? m?�?�?�?�?�? OO $O�?HO3OlOWO|O�O ����Oӯ�O�O�O!_ _E_3_i_W_�_{_�_ �_�_�_�_o�_/oo ?oAoSo�owo�o�o�o �o�o�o+O= s�E���Y�� ���9�'�]�K�m� ������u�Ǐɏۏ� ��5�G�Y�k�%���}� ����ßşן���1� �U�C�y�g������� ӯ������	�+�-� ?�u�c���������� Ͽ���/�A�S��� ��qϓϕϧ������ ��%�7�I�[���m� �ߑ߳������߷�� 3�!�W�E�{�i��� �����������A� /�e�S�u��������� ������+a O�s��e��� ��'K9o] ������� #//G/5/k/}/�/�/ [/�/�/�/�/�/?? C?1?g?U?�?y?�?�? �?�?�?	O�?-OOQO ?OaO�OuO�O�O�O�O �O�O___M_�e_ w_�_3_�_�_�_�_�_ oo7o%o[omoo�o Oo�o�o�o�o�o! 3�o�oiW�{� ������/�� S�A�w�e�������я �������=�+�M� s�a���������ߟ� �_	���_ן]�K��� o�������ۯɯ��� #���Y�G�}�k��� ��ſ׿������� �U�C�y�gϝϋ��� ���������	�?�-� c�Q�s�u߇߽߫��� �����)��9�_�M� ����/����i���� ��%��I�7�m�[��� ���������������� EWi{5�� ������A /eS�w��� ��/�+//O/=/ _/a/s/�/�/�/�/�/ �/?'?��??Q?c?? �?�?�?�?�?�?�?O �?5OGOYOkO)O�O}Op�O�O�O�N  �@�S V_R��$TBJOP_G�RP 2,�E��  ?��V	-R4S.;\=��@|u0{S~PU >��U�T @�@LR	� �C� �Vf?  C���ULQ�LQ>�33�U�R�����U�Y?�@=��ZC��P�����R��P  Bȸ�W$o/gC��@g��dDb�^�㙚eeao�P&ff~�e=�7LC/kFaB o�o�P��P��efb-C�p�B�^g`�d�o�PL�P�t<�eVC\ � �Q@�'p�`��  A�oL`��_wC�BrD��S�^�]�_�S�`<PB��P�anaaF`C�;�`L�w��aQoxp�x�p:���XB$'tMP@�PCHS��n����=�P����trd<M�gE�2pb����X �	��1��)�W��� c������������ 󟭟7�Q�;�I�w����;d�Vɡ�U	�V3.00RSc7r35QT*�QT��A�� E��'E�i�F�V#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG��G#
�D���E'
E�MKE���E��ɑE�ۘE���E���F���F��F���F(��F�5��FB��F�O��F\��F�i��Fv��F���vF�u�<#�
<t����ٵ=�_��V �R�p�V9�~ ]ESTPARtp��HFP*SHR\�A�BLE 1/;[$%�SG�� �W�
G�G�G� WQG�	G�
G�GȖ�QG�G�G�ܱv�'RDI~�EQ�ϧ� ��������W�O_�q�@{ߍߟ߱���w�S]�CS !ڄ������ ������&�8�J�\� n������������� ] \�`��	��(�:� ����
��.�@�w��NUM  �EUEQ�P	P ۰�ܰw�_CFG �0��)r-PIMEBF_TTb��CSo�,VERڳ-B�,R 11;[' 8��R�@� �@&  ��� ����//)/;/ M/_/q/�/�/�/�/�/ ?�/?J?%?7?M?[? m?>�@�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_��_l_�Y@c�Y�MI_CHAN�8 c cDBGLV��:cX�	`�ETHERAD �?f�\`���?�_uo�oQ�	`RO�UTV!	
!��d�o�lSNMAS�KQhcba255.uߣ'9ߣY��OOLOFS_D�Ib��U;iORQCTRL 2		�Ϸ~T��� ��#�5�G�Y�k�}� ������ŏ׏�����.��R�V�PE_�DETAI/h|zP�GL_CONFI�G 8�	����/cell/$�CID$/grp1V�̟ޟ�������o?�Q�c�u����� (���ϯ������ ;�M�_�q�����$�6� ˿ݿ���%ϴ�I� [�m�ϑϣ�2����� �����!߰���W�i� {ߍߟ߱�%}F��� ����/�A�C�i�H�Eߞ�������� ��?��.�@�R�d�v� ������������� ��*<N`r� ������& 8J\n��!� ����/�4/F/ X/j/|/�//�/�/�/ �/�/??�/B?T?f? x?�?�?+?�?�?�?�? OO�?>OPObOtO�O��O�O���Us�er View ���}}1234567890�O�O�O�_#_5_=T�P��]_���I2�I:O�_�_�_@�_�_�_X_j_�B3�_ GoYoko}o�o�o o�op^46o�o1CU�ovp^5�o������	�h*�p^6 �c�u����������ޏp^7R��)�;�M� _�q�Џ��p^8�˟ ݟ���%���F�L�� lCamera�J���� ����ӯ���E~�� !�3��OM�_�q��������y  e��Yz��� 	��-�?�Q���uχ� ��俽���������>��e�5i��c�u߇� �߽߫�d������P� )�;�M�_�q��*�<� �i���������)� ��M�_�q�������� ��������<�û��= Oas��>��� �*'9K] f�Q������ �/�%/7/I/�m/ /�/�/�/�/n<�� ^/?%?7?I?[?m?/ �?�?�? ?�?�?�?O !O3O�/<׹��?O�O �O�O�O�O�?�O_!_ lOE_W_i_{_�_�_FOXG9+_�_�_oo(o :o�OKopo�o)_�o�o@�o�o�o ��	g�0�oM_q��� No����o�%�7� I�[�m�&l�n�� Ə؏���� ��D� V�h���������ԟ 柍�g�ڻ}�2�D�V� h�z���3���¯ԯ� ��
��.�@�R���3u F�鯞���¿Կ��� ���.�@ϋ�d�vψ� �ϬϾ�e�w���U�
� �.�@�R�d�ψߚ� ������������*� ��w���v���� ����w�����c�<� N�`�r�����=�w�� -�����*<�� `r�������x���  �� 1CUgy��������    -/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_�i_�  
��( � �%( 	 y_�_�_�_�_�_�_ o	o+o-o?ouoco�o�o�o�Z* � Q&�J\n ������o��� 9�(�:�L�^�p�� �������܏� �� $�6�}�Z�l�~�ŏ�� ��Ɵ؟���C�U�2� D�V���z�������¯ ԯ���
��c�@�R� d�v�����᯾�п� )���*�<�N�`ϧ� ���ϨϺ������� �&�8��\�n߀��� �߶���������E�"� 4�F��j�|���� ��������e�B� T�f�x����������� ��+�,>Pb ���������� (o�^p� ������ /G $/6/H/�l/~/�/�/ �/�//�/�/?U/2?�D?V?h?z?�?�/�`@� �2�?�?�?�3��7�P��!frh�:\tpgl\r�obots\m2�0ia\cr35?ia.xml�?;O MO_OqO�O�O�O�O�O�O�O ���O_(_ :_L_^_p_�_�_�_�_ �_�_�O�_o$o6oHo Zolo~o�o�o�o�o�o �_�o 2DVh z������o� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟�ݟ��&�8� J�\�n���������ȯ ߟٯ���"�4�F�X� j�|�������Ŀ־�8�.1 �?@8?8�?�ֻ� ֿ�3�5�G�iϓ�}� ���ϳ��������5߀�A�k�U�wߡ߿���$TPGL_OUTPUT ;�!��! �� ������,�>�P�b� t����������� ��(�:�L�^�p������������2345678901�� �������"�� BTfx��4�@����
}$ L^p��,>� �� //$/�2/Z/ l/~/�/�/:/�/�/�/ �/? ?�/�/V?h?z? �?�?�?H?�?�?�?
O O.O�?<OdOvO�O�O �ODOVO�O�O__*_ <_�OJ_r_�_�_�_�_ R_�_�_oo&o8o�_ �_no�o�o�o�o�o`o �o�o"4F�oT�|����\��} �����0�B�T�e��@������� ( 	 ��Џ��� ���<�*�L�N�`� ��������ޟ̟�� �8�&�\�J���n��� ������ȯ���"�������*�X�j�F��� ��|�¿Կ��C���� ��3�E�#�i�{�忇� ��S����������/� ��S�e�߉ߛ�y߿� ��;�������=�O� -�s���ߩ��]��� �����'����]�o� �����������E��� ��5G%W}�� ����g��� 1�Ug	w�{ ��=O	//�?/ Q///u/�/��/�/_/ �/�/�/�/)?;?�/_? q??�?�?�?�?�?G? �?O�?OIO[O9OO �O�?�O�OiO�O�O�O !_3_�O_i_{__�_�_�_�_�_�R�$T�POFF_LIM� >�op:�y�mqbN_SV`�  l�jP_�MON <6�)dopop2l�a�STRTCHK �=6�f� bVTCOMPAT-h��afVWVAR �>Mm�h1d ��o �oop`b�a_DEFPRO�G %|j%OLPTES�`H�l�_DISPLAY�`|n"rINST_�MSK  t| �^zINUSER��odtLCK�|}{QUICKMEN��dtSCRE�p�6��btpsc@dt�q��b*�_.��ST�jiRACE_CFG ?Mi��d`	�d
?��u�HNL 2@"|i����k r͏ ߏ���'�9�K�]��w�ITEM 2A��� �%$12�34567890<����  =<��П<��  !���p��=��c��^� ���������.���R� �v�"�H�ί��Я� �����*�ֿ���r� 2ϖ�����4�޿�ϰ� ��&���J�\�n���@� ��d�v��ς������ 4���X��*��@�� ���ߨ������� T���x������l� �������,�>�P��� ����FX��d���� ��:�p" ��o����� F6HZt~�� N/t/�/��// /2/ �/V/?(?:?�/F?�/ �/�/j?�??�?�?R? �?v?�?QO�?lO�?�O �OO�O*O|O_`O _ �O0_V_h_�Ot_�O_ _�_8_�_
oo�_@o �_�_�_Lodo�_�o�o 4o�oXojo3�oN�o r��o��s��S�B���z� 3 h��z ��C�:y
 P�v�]���~�UD1:\������qR_GRP� 1C��� 	 @Cp���@$��H�6�l�Z��|� ����f���˟���ڕ?�  
���<� *�`�N���r������� ޯ̯��&��J�8�Z���	�u�����s�SCB 2D� �����(�:��L�^�pς��|V_C�ONFIG E����@����ϖ�OUTPUT F�������6�H� Z�l�~ߐߢߴ����� �������#�6�H�Z� l�~���������� ����2�D�V�h�z� ��������������
 �.@Rdv�� �����) <N`r���� ���//%8/J/ \/n/�/�/�/�/�/�/ �/�/?!/4?F?X?j? |?�?�?�?�?�?�?�? OO/?BOTOfOxO�O �O�O�O�O�O�O__ +O>_P_b_t_�_�_�_ �_�_�_�_oo'_:o Lo^opo�o�o�o�o�o �o�o $����!� bt������ ���(�:�-o^�p� ��������ʏ܏� � �$�6�G�Z�l�~��� ����Ɵ؟���� � 2�D�U�h�z������� ¯ԯ���
��.�@� Q�d�v���������п �����*�<�M�`� rτϖϨϺ������� ��&�8�J�[�n߀� �ߤ߶���������� "�4�F�W�j�|��� ������������0� B�S�f�x��������� ������,>P a�t��������(:L/x���k}gV �K���//&/ 8/J/\/n/�/�/�/W �/�/�/�/?"?4?F? X?j?|?�?�?�?�/�? �?�?OO0OBOTOfO xO�O�O�O�?�O�O�O __,_>_P_b_t_�_ �_�_�O�_�_�_oo (o:oLo^opo�o�o�o �o�_�o�o $6 HZl~����o ���� �2�D�V� h�z��������ԏ� ��
��.�@�R�d�v� ��������Ϗ���� �*�<�N�`�r����� ����˟ޯ���&� 8�J�\�n����������Ż�$TX_SCREEN 1G�g�}�ipnl/��g?en.htmſ��*�<�N�`ϽP�anel setupd�}�dϥϷ����������ω�6� H�Z�l�~ߐ�ߴ�+� ������� �2�߻� h�z������9�g� ]�
��.�@�R�d��� ������������� }���<N`r�� ;1��& 8�\��������QȾUALR�M_MSG ?��� �Ȫ-/ ?/p/c/�/�/�/�/�/ �/�/??6?)?Z?%�SEV  -��6"ECFG �I��  }ȥ@�  A�1�   B�Ȥ
 [?ϣ��?OO%O 7OIO[OmOO�O�O�G~�1GRP 2J�;w 0Ȧ	 �?��O I_BBL_NOTE K�:�T��l�Ϣ�ѡ�0RDE�FPRO %+ (%N?u_Ѡc_�_ �_�_�_�_�_o�_o�>o)oboMo�o\INUSER  R]��O�oI_MENH�IST 1L�9 � ( _P���)/SOFTP�ART/GENL�INK?curr�ent=menu�page,1133,1�oDVhz~�(
50������q,��ued�it(rOLPTEST�M�_�q�|~|o ����ʏ܏� ���$� 6�H�Z�l�~������ Ɵ؟�������2�D� V�h�z������¯ԯ ���
��h9Rq��B� T�f�x���������ҿ ����ϩ�>�P�b� tφϘ�'�9������� ��(߷�L�^�p߂� �ߦ�5������� �� $����Z�l�~��� ��C�������� �2� �/�h�z��������� ������
.@�� dv�����_ �*<N�r �����[�/ /&/8/J/\/��/�/ �/�/�/�/i/�/?"? 4?F?X?C�U��?�?�? �?�?�?�/OO0OBO TOfO�?�O�O�O�O�O �O�O�O_,_>_P_b_ t__�_�_�_�_�_�_ �_o(o:oLo^opo�o o�o�o�o�o�o �o $6HZl~i?{? ������2� D�V�h�z����-� ԏ���
����@�R� d�v�����)���П� ��������N�`�r� ������7�̯ޯ�� �&���J�\�n�����������$UI_�PANEDATA 1N���ڱ�  	��}  frh/�cgtp/who�ledev.st�m���&�8�J�Y�)  riρ�@�� �ϫϽ�������Z�� )��M�4�q߃�jߧ� �����������%�7���[�7�� � �    ,��Ϙ����� ����E����:�L�^� p�������������� ��$H/l~ e������o�ܳ7�<N`r ����-���/ /&/8/�\/n/U/�/ y/�/�/�/�/�/?�/ 4?F?-?j?Q?�?�? %�?�?�?OO0O�? TO�xO�O�O�O�O�O �OKO_�O,__P_b_ I_�_m_�_�_�_�_�_ oo�_:o�?�?po�o �o�o�o�oo�o sO $6HZl~�o� ������ �2� �V�=�z���s����� ԏGoYo�.�@�R� d�v�ɏ����П� �����<�N�5�r� Y�������̯���ׯ �&��J�1�n���� ���ȿڿ����c� 4ϧ�X�j�|ώϠϲ� ��+��������0�B� )�f�Mߊߜ߃��ߧ� ��������P�b� t����������S� ��(�:�L�^���� i�����������  ��6ZlS�w�'�9�}���"4FX)�}�� l�����/j '//K/2/D/�/h/�/ �/�/�/�/�/�/#?5?�?Y?��C�=��$U�I_POSTYP�E  C�?� 	 e?�?��2QUICKME/N  �;�?�?��0RESTORE� 1OC�?  �L?��!6OCC1O��maO�O �O�O�O�OuO�O__ ,_>_�Ob_t_�_�_�_ UO�_�_�_M_o(o:o Lo^oo�o�o�o�o�o �oo $6H�_ Ugy�o���� �� �2�D�V�h�� ������ԏ��� �w�)�R�d�v����� =���П������*� <�N�`�r������� �ޯ���&�ɯJ� \�n�������G�ȿڿ������7SCRE��0?�=uw1sc+@u2K�U3K�4K�5K�6K��7K�8K��2USE�R-�2�D�T,�M�k�sUô�4��5��6ʴ�7��8���0ND�O_CFG P�;� ��0PDAT�E ����None�2��_I�NFO 1QC�@��10%�[���I� ��m߮��ߣ������� ���>�P�3�t��i�����<-�OFFSE/T T�=�ﲳ $@������1�^�U� g�������������� ��$-ZQcu����?�
����U�FRAME  ���*�RTOL_ABRT	(�!�ENB*GRP� 1UI�1Cz  A��~��~ ���������0UJ�9MS�K  M@�;N%8�%��/�2oVCCM��V��V�#RG�#Y�9����/����D�BH��p71C����3711?�C0�$MRf2_�*S�Ҵ��	���~XC�56 *�?�6����1$�5���A�@3C��. ��8�?��OOKOx1FOsO�5�51���_O�O�� B����A2�DWO�O 7O_�O8_#_\_G_�_ k_}_�__�_�_�_�_�"o�OFoXo�%TCC��#`mI1�i������� GFS��2�aZ; �| 23�45678901 �o�b�����o�� !5a�4BwB�`56� 311:�o=L�Br5v1�1~1�2�� }/��o�a��#� GYk}�p��� ����ُ�1�C�U� 6�H���5�~���ߏ����	���4�dSEL#EC)M!v1b3��VIRTSYNC��� ���%�SI?ONTMOU�������F��#bU��U�(u FR:\H��\�A\�� �߀ MC��LO�G��   UD�1��EX����'� B@ �����̡m��̡RO�BCL�1�H� ��  =	 �1- n6  G-������[�,S�<A�`=��͗���ˢ��TRAIAN⯞b�a1l�
0�d�$j�T2cZ; (aE2ϖ�i��;� )�_�M�g�qσϕϧπ�������	��F�S?TAT dm~2!@�zߌ�*j$i߾߮�_GE�#eZ;��`0�
� 02���HOMIN� f�U��U� P~�����БC�g�X����JMPERR {2gZ;
  �� *jl�V�7�������� ������
��2�@�q�hd�v�B�_ߠRE� �hWޠ$LEX��i�Z;�a1-e��VM�PHASE  �5��c&��!OFFX/�F�P2n�j�0�㜳E1@���0ϒE1!1?s33�����ak/�k�xk䜣!W�m[�� ���[����o3;� [i {����/ �O�?/M/_/q/� �/��//�/'/9/�/ =?7?I?s?�/�?�/�/ �?�??Om?O%O3O EO�?�?�O�?�O�O�? �O�O�O__gO\_�O E_�O�_�O�O/_�_�_ �_oQ_Fou_�_|o�o �_�oo�o�o�o�o;o Mo?qof-�oI� ����7�[ P���������ˏ ��!�3�(�:�i�[��ŏg�}������TD�_FILTEW�n��� �ֲ:��� @���+�=�O�a�s� ��������֯��� ��0�B�T�f�x����SHIFTMENoU 1o[�<��%��ֿ����ڿ�� ��I� �2��V�hώ� �Ϟϰ�������3�
��	LIVE/S�NAP'�vsf�liv��E��^��ION * Ub�h�menu~߃��`���ߣ���p����	����E�.�5T0�s�P�@� ���AɠB8z�z���}��x�~�P��c ���MEbЩ��<�0���M�O��q���z�W�AITDINEN�D������OK�1�OUT���S�D��TIM����o�G���#���C����b������REL�EASE������T�M�������_A�CT[�����_D?ATA r���%L����xRDI�Sb�E�$XV�R�s���$ZA�BC_GRP 1Ut�Q�,#�0�2���ZIP�u�'�&����[M�PCF_G 1v��Q�0�/� wx�ɤ� 	�>Z/  85�/0�/H/�/l$?��+�/ �/�/?�/�/???r?>�?  �D0�? �?�?�?�?�;����x�]hYLINuD֑y� ��� ,(  *VO�gM.�SO�OwO�O�M i?�O�O^PO1_�O U_<_N_�_�O�_�_�_ _�_�_x_-ooQo8o`�_�o�oY&#2z�� ���oC�e?�a?>N|�oq�����qA�$DSPHE_RE 2{6M��_ �;o���!�io| W�i��_��,��Ï�� �Ώ@��/�v���e� ؏��p���������l�ZZ�� �N