��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk" 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&@B4��_sC3���r[R�_p�d`U��@VAD>CMVROU
b�1�PERIO�sF1P���2D-��3%T��1_D��2�Ĥ�3��T����K�9K��K�7CL���0�gADJ����_Udr;[PAUX�@�_	 4�@C�P?a$� A�&�n@ ~qUX_AXS��XSMC�� 
 h�D�rӠ�Cd� �C�t�C�F�@�H�G1P��FOXp4XAXISU� Tj��D͡ȹq�E��AP@M@ �	BQ܀HR
$I�DX\PRV�PSa�G�RT�L $�F�E_Uנ���TTOOL�R�p;�A��p�y1DOf`� \��0R_PK�G�RQ BQ SNR�PBQS�P=[Q 2	hQ2�P�S�P2�Q�Q�ba	�1�ad�$VFLfw0IM�,�LT�r �:a��Tc�6Tb�����$DYG��C$d0JgGUg	�d�4�d��cMPSWP� ��$ @��  �{���a   &�`� &�`VERSI�ON�h � �5�aIRT�UAL�o�avS?��h&�  �aL|J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B��T�f�x��a+u|P11w 29{\�`p�� ֓Ә���  ?�a� @�`����A�  �����#���� 3��-�?�Q�?�g��U����  D � Bp  =���Ϳ�?333?��a�̠�̤@��ߥA� ��/  & G�P ?fffˡ>��ߥ����� ��0�ܙD���̤ˡ� �k�C�Z�[��`�0�`����ӿٲ��B�ђ I@ɟK�ÿ��;���F@ K���������Dz��l�W�I�ψٺ��ܑ�P`��w���ēV��'�9�K� ]�o�5ߓ���_�q�ۿ �������#�9�G� y�7�I�j�߳����� ������a��!���y�3����ϋ�9�K� ]�oρϓϙ���x��� D����������� ,>�b������� �����0�����ȗ�Đ ؓ���2/d���L� ���^/\�Ϣ�]�ĐPW��"�`�"��'B����������/"  A$đƚ�$1>B,4_��(����1?��?<�?�8>����ā� //@/�?T/f/?O�/ �/�/�/�/�/�O?? ,?>?P?b?;_�?__�? �?�?�?�?OO(O�_ o^OpO�O�O�O�O�O �O�O __$_�oH_Z_ 3~_�W��fx���2�����	��	�o2�2-�V�h�z� ������ԏ����� ���Dqdd�����l�� ߩߩ�b�����o���� ğ���cd�p(�������qT�@� a>�Ho�
}��[��c|��>LŠ���_v���<'#�
�Qsbp|��pX��o�C��� a@?e?a��3�T`��@ � ��G_�
�T���_�� ��x�2bo%{Bta�� �����1��U�g�k�`>X�ؤ����ϑ��It$ ��$$�>%�٢
���A�����'�����4�+��=�s�.���Ճa�$敕��(4$�ܛ�S�e�;��.���>��H�Ճa5�����8M�Y��;�=���3��a�B�	9�R�=�v�a�� �����������m��|��  �b \'������`k�S�K� X�,�w�������/������C��Q�??333;�s�<��sa�D/  C``GÿP ?fff/a> $���?_	W�_��0� �_g�;�5c?� 4'e��u�j� F@ ��[�� DzI ����w5����y � ������/�� �/�/7I�_I/[/m/ /�/�/�/�?�?�?�/ ?!?3?E?W?i?{?�? kO}O�?�?�L�Oq �O�������O ���O�O�_
__._@_ R_d_o�_�_,o�_o �_�_oobo%`&/0 $.(��?�� >�"��o����}��o ��E+̰�B��+�� ȴC��8�����{j4� ~gĠ{t��"�������$�3t7�q�����>���3t�c u�������� ��)�W���_�q��� ��������ݏ�ȯ� %�7�I�k�%����j� ��ǟٟ���Ϳ3� E�W�i�{�a������� կ�L�o0�������Ł2Q/�A�S�e�v�Uώ�2�߲������� ����0�B�T�[R u���������7M;	 ;	/�DO*GT�V� �M�D�i���Op����P�Ѱ����A>�a���f��2�BH���>�L! H���g�<#�
�ϲp��w�E8�v������A�� 7������@\A �b�f��D?B,��7J���_���Bб��� Z{�p��N����>�4_�U�/��I�t$ //$��>�5
/a'A��a/	/��/-/?&��+��̞�%.����%��$�敕�%(4$�x�%�/�+;��.#5�>��H/5��5{��?58M�YK5��= g5��8�x?�+	�/�?�?�?�7?�? O$O6OHOZO�o�Gn>lG  ;¸` �X���E�E��A ��O�O�O	_�2 _^ʫ���`=�e?3�33���B�����D�/  C��G�P_ ?fff��>� ��e�Y�Q�iȌOVb �m����W�i�]ooo �o��k��_wo�o�`F@ uawU�`Dz�P$to�op�jn���� ��_ �_oo'o�KoU� )��o�oﯥ��� ��1���"�Y�k� }�������ŏ׏�ǟٟX�1��̸k��oC� �o'9KQ��� 0�B���f�x������� ��z�������l�>� P�b�t���lu�ς\�nπϊx�O����� ��4�����C�<� ��R(����c�$ �C� ���׺��ڷ   �Ę�~Jk���_V�؏��/�?�Q�]�>�����]���� ������+��O�a� s߅߳�U��������� ����9�K�$o�� ����������� #�5�G�u�k�)���� ����������1�ǼZό�/0/B/X%2@�l�/�/�/�/�-��"2�/? ?2?D?V? h?z?�?�?�?�d�n�> �GYGZ<���Y�Y �������ijO|O�O�O�FK �GLO^I(b!W�#�> �'_�����4U>L�}PdQ�.B�<#�	
K+p4_�B�t�FB�����SU�RkU@��lT�� o�δ���ζ��0o��eB,TUPo�o��o�o�o��P>�a�T�O�OrICItk$ �$�&>��R	
k�wAHD�e�x��v�@+���+��.���7��A$�{��G�(4$�S����;��.�>���H���A5�=���8M�Y���=�=dPÅ�B�ԏ�{	 �
���.��g�Y�n� ��������%o�=��ȗ  B��R �T_b�P#��J��X /�A�S�e��|�j�B��	��S��?33�3�E+��D7IcaD/�  CG�P /?fff�A>�Q8D ����O=X蟲�� M�O���o��˿쿀��?Y�ӿ-�Kl�F@ _�k�ӥbl�Dz���k�]�/��8~!^/P) �;�M� _�q���Iߧ���s߅� ��K��%�7�M� [ߍ�K�]�~������ �����!�3�u�#�5����Sl���)ϟ�M� _�qσϕϧϭ�GR�� ��X��������
 �@R�v��� ����/�ϸ����ȫ�� vi ڗ�N.k_=C��/o� 㢄`s���U�"�d�Q �f�PcEci3�/6|P 3$�ښ�$E>�Us��(���)o�<�?�8>�����:/-/?/ Q/c/u/�/`O�/�/�/ �/?�O?)?;?M?_? q?J_�?�?�_�?�?�? O#O�_7OIO"omOO �O�O�O�O�o�O�O_ !_3_oW_i_B�_{�@��z���u2	� ����.�F�2A�j�|�������ď ֏�����
�-�Xq xd�����l�����b �����Ɵ؟���!�wd�p<������qh�T�_a>\��}pz�o� s��>L٠��� o��y<#�
�Q�bp��/�l��o.�c���_aSeWa��G�h`ǥ@�Ȥ[s� �T���_�V�ꌿFbo9{B�a�����3�@E�(�i�{�.k�>l������ϥ�It$� ��$8�>��
���A�����;��ϼ��H�+��̇�.������G�$�=���(4$ܯ�g��y�;��.��>���H��G�5�����8M�Y�O�=@���G��a0�V�	M� f�Q��u��ߵ������� ����'��$�  �bp;�� ����g�_�l�@����������C�����c���e��S?333�O���P���ñD/ � Ct`G�P ?fffO�>8���S s	k�_!xD�s{� O�IwS�'H;e�#��/��j� F�@ ��/o�� Dz] ����I�q��y ܗ�� ���//�/�/K ]�_]/o/�/�/�/�/ �/�?�?�??#?5?G? Y?k?}?�?�?O�OO�?g|�#O��O�� ���/	_���O�O �__0_B_T_f_x_2o �_�_@o�_$o�_oo ,ovo$%t:/&8B(�OPp\cҹ6� �o�~ǯ���o��E? ��BPp?��ܴW��� L������jH��gؠ�t Pq6�#������8�Gt�K߅���	��>���Gt�w��� �������+�=� k��s���������͏ ����ܯ'�9�K�]� �9�����~�ɟ۟� ��-�#��G�Y�k�}� ��u���ů���l D�������2eCߐU�g�yߊ�iϢ�2 ����������� �2� D�V�h�of���Դ ������KMO	O	C�XO >Gh�j"�4�a�X�}�ӴИ������
��p�>�a��z��B8�B\���>L5 x\���{�<#�
��p�����E,ϊ�����p������İ#@pA$�b�z� B�SB@�KJ���s���B�n�� �����t >�H�s�i�*/�It$ ZC/$��>�I
#/u'A �u//�/A/S&ޤ�+����%.�����%��$敕�%(4$�5�/�+�;��.75>��yHC5��5��S5O8M�Y_5��=  {5��L��?�+	�/�? �?�?�7?O&O8OJO�\OnO}K�$CCS�CH_GRP12 2����A�&� �\��Xo��  O��`�lt �E �E���A�__,_>_P�2U_C^����`Q�e?333��R��|��#D/  Cа�G�P ?fff��>���e�Y�Q� }��Ojb�m����W�i ��o�o�o���2o�ox�E`F@ 8u0Da�U�E`Dz�PYt�Do6�j6��� �o&o8oJo\o"� �o�L�^��o�o�� ���&�4�f�$�6� W�������ď֏�����N������f�� ��x�&8J\n �����e�w�1����� ��ѯ������+��� O���s��������u��Ϸ�ϣϵϿx� ����ٳ.��i�'�# ��x�q�H��R<L��� ���8�W� � ����4 ����J�� �sLV�����/�xt���>����� ������*�<�N�`� 9��ߖߨߺ��ߊ��� ��&�8�J�#n�� Y���������� "��F�X�j�|����� ^���������0 B/f�����S/e/w/�%2�l�/�/�/�/=�22?C?U? g?y?�?�?�?�?�?�? �d�nN1!Q|Y|Zq ȝ�Y�Y�՟����i@�O�O�O�O�FP� @W�O�I�!AW-3�>5�\_�S�H��iU>L�P�Q�cB�O<#�
�`pi_�RE��V<B����,0�U bA�U@ 푡T4�Lo��В�@fȚeo��Ba �U�o�oBT�P>Ea�T�O�O�^~CIt$ �$6K>��R
��wA}D������v!P+�{��`�.���l�� Q$敕|�(4�$܈�@�R�;��=.��>��H�� Q�5��Ѕ8M�	Y܅(M=�P�� R�	�/�	&�?�*�c�N� ��������ǟٟ�Zo� Mؾ��   �I�b�T�b�PX�@� 8JE�hd�v������(����<B�>��S,�?333(U`�)TlI��aD/  CMG�P ?fff(Q>amD,�L�D��� ��L�TM(_"�P�, � �!��?���b�<���F@ �Š��Hb��Dz6��Ġ����d�"ʳ!�/�) �p���������~�ܿ �Ϩߺ�$�6π6�H� Z�l߂ߐ��߀��� ����� �2�D�V�h�@��X�j��������� ^����ϔϦϸ����� ��|R�������	 -?Qu�� ����O��M/`���/���� ) 5�i���.�_nC ��/����`��) e �"�d0a�f%`�E�ih !?k�Ph$)!��$z>�U��8 $$�^o�<<�?�8>��� $�: P/b/t/�/�/�/�/�O �/�/??D?�OL?^? p?�?�?�?_�?�?�_  OO$O6OXOolO~O Wo�O�O�O�O_�O�o  _2_D_V_h_No�_�_ w�_l�/����u2>��.�@�R�c�	B{�2v�����Ï Տ�����/�A�H� ?�b��q�dةت�l$� (�(�r1��AC��� �:�1�V��d�pq��ݟ��q����Ia>����S}���5sť�>L���5o��Ty<'#�
�Q�bpůd�p��c�����Ia@�e�a�|��`��@I� �����Sd,�o۶ $���{bLon{B�a� �G�h�z�]Ϟϰ�ckM�>��!�L�B��ړ�It$ �$m�>%�"�
��N�AٔN����p��,�}�+��=̼�.�����|��$敕��(4$���՜߮�;��.��>��H�|�5���,�8M�Y8儝=��T�|�%qe���	�ߛ������ �����#�5�G���\�|4Y�  (r �p�E��M������� ��u���������x��������*��?333����ș���D/  C�`GÿP ?fff��> m�ɔ��	��_Vxy� C�����~���J \}peX��d��j� F@ ��d��� Dz� $����~���y � ����/8B/ ??���_�/�/�/ �/�/�/?�?�?OF? X?j?|?�?�?�?�?O �O�OEOO�L�XO� 0_��//&/8/>_ آ_/_�_S_e_w_�_ �_�_go�_�_uooYo +o=oOoao�oY%�o/0I[mw(�<O�p �c�k�!�~��Γ0 )� Ut�R�pt�P� Č�0Ɓ������j}� �g��t�qk�X�֎L�m�|t�ߺ�,�>�J�>���|tJ�� �������<� N�`�r���B�����̏ ޏ���ۯ&�8��\� n�������n�ȟڟ�� ���"�4�b�X��|� ������į������� �p�Gy��/�EՁ2�xߊߜ߮߿�����2������1� C�U�g�y���� ����	�4	4
)̀M�	 �	xOsG�ϟW�i��������8���9�PK�O����� Q>�a���R R��!>�Lj Q����<#�
8��p!���E8aϿ����� Q� �@���X@�AY �b��w��Bu�7�Jײ����B�A= �����/��� �>�}����_/6�I�t$ x/$��>�~
X/�'A5��/R/��/v/�&��+��̞5.���$5��$�敕45(4$�x@5�/
;;��.l5�>��Hx5��5{���58M�Y�5��=Q �5����?�+	�/�?�?OGT?FO [OmOO�O�O��n>�G  ��p ��L� U�E���A �_._@_R_�2i_W^�����`��e?3�33��R��$�XD�/  C�G�P_ ?fff��>� -��ei�Q<����O�b }����Wy��o�o �o̵��Fo�o8�Y`F@ LuXa�U Y`Dz�PmtXoJp�jk�K�=� �(o :oLo^opo6��o�`� r��o�o8�� ��$� :�H�z�8�J�k����� Ə؏���� �b��"���z�4������ :L^p����4 y���E�����ӯ��� 	�ÿ-�?�ѿc����� ������ϵu���������xȘ���� c�G}�;�X&�υ� \��Rq`������m ��� P�P ���#� i  ����J��2�`V�����/����>����Ħ��� ,�>�P�b�t�M��ߪ� �����ߞ���(�:� L�^�7���m���� ������$�6�Z� l�~�������r���� �� DV//z������g/y/�/�%2@�l�/�/�/
?=�322.?W?i?{?�?�? �?�?�?�?�? t�nN E!e�Y�Z�ܝ�Y�Y ��ϗ��i�O�O�O�OVd� )W�O�I(�!UWA3L>I�p_�-g�\��}U>L��P�Q�wB)<#�	
�tp}_RY��VPB��L@D�U4bU�U@��TH� `o/����fܚyo3&+Bu�U�o�o� 2Vh`>�Ya�T_�O��CItk$ �$%6>��R	
��A�D��(�x��v5P+���t��.�����4Q$�{����(4$ܜ��T�f�;��.ȅ>���Hԅ4Q5�=��8M�Y��<M�=�P�4R��C�	 :�S�>�w�b������� ɟ۟���noM��  �]�(b �T�b`l�T�LJY�-h x�������0�ů��PB��R��S@�?33�3<Ut�=T�I�aD/�  CaG�P /?fff<Q>%a�D @�`�X��(1���`� hM<_6�d�@��5π(O���vϔ��F@ �Ŵ��\b��DzJ��Ĵ���x�6�8�!�/�) ܄��� ����̿����ϼ��� 8�JϔJ�\�n߀ߖ� ���ߔ�������"� 4�F�X�j�|��l�~��������r����� �Ϻ����������R�� ���/ASe ��-��� c�a/'�//%//����= I�i #���.�_~C��/�� ,��`��= ,e2�dDa �f9`�E�i|5?�P |$=!#�4�>e��%8�4$8�ro�<�?H>���4$Jd/v/�/ �/�/�/�/�O�/?? *?X?�O`?r?�?�?�? �?�_�?�?�_O&O8O JOlO&o�O�Oko�O�O �O�O__�o4_F_X_ j_|_bo�_�_��_(l@�1/����u2R� 0�B�T�f�w�V��2����ŏ׏���� �1�C�U�\�S�v��q �d���l8�<�<�0r E�+�UW��!�N�E�j��d�p���������]a>�̯g}p���Is٥>L"��	�IoӒhy<#�
�Q�bpٯx���w�����]a�e�a�����`�@]����� g/d@�-o�8�տ�b`o�{B�a����[�|�@��qϲ���wka�>���5�`�V���It$� 0�$��>�6�
�b�A�b�
߄�.߼@֑�+�����.�����Ր�$�=���(4$��հ����;��.$�>���H0吡5���@�8M�YL嘝=@	�h吢9qy��	�� ����������%��7�I�[�j��$CC�SCH_GRP1�3 2������&� �\�~E�y  <r���Y��a� �����������+��B0����<>��?333�������ܙ�D/  C��`G�P ?fff��>��ᔜ�	� �_jx��W�ĝ��� ������el����j2F@ `%%1���2Dz�  F$1#/��#���y �%7I ?mw/9?K?���_ �/�/�/�/?!?S?O #ODO{?�?�?�?�?�? �?�?;O�O�OzOSO\��O�e_/%/7/I/ [/m/s_�R_d_o�_ �_�_�_�_�_�ooo �o<o�o`oro�o�o�o��%��/~���(�qO�p�cɠ�V� �ޓe^�5U�)�9R �p����%Ġ�Dƕ�� ��j���g!��t�q��@���`�9���t���οa�s��>��� �t�����)�;� M�&�q�������Տw� ݏ���%�7��[� m�F�������ǟ韣� ����3�E�W�i��� ��Kϱ�ïկ���߿ �/��S���|�@�R�d�z�2��߿���$�������2�0� B�T�f�x������ �������>�i	i
 ^̵M�	�	���O�G�π�����������=��m�n�����.�ڱ>"qI��@R5R��V>L� �ƿP���<#�
m�M�p�V��2U����)���ڱ��u.��@�A�!r9�Ϭ��B���l�JR�ݿ��B N�vr��/�//A/��� >2�������/k�It$ �/$���>��
�/�'A�j��/�/?�/�& +����M5.����Y5$敕i5(�4$�u5-??;;�{�.�5>��H�5�5���58M�Y�5�=� �5���?;	?,OOPO ;G�?{O�O�O�O�O�O�G���n�G  ��6p��� EU -U%�2QQ_c_u_�_P	B�_�^)��+p�u?333MR|Y��D/  C:��G�P ?fff>�Z�u9i1aq� ��
_�b9}A�g=y /�o�o���{o�oxOmʎ`F@ �u0�a�U5�`Dz#`�t��oQz�р�r� �]ooo�o�o�ok� �o�����#m�#� 5�G�Y�o�}���m�� ��׏�����1�C��U���E�W�֟��i�� �K��o���� �ϯi����z���� ��,�>���b�t�� ��꿼�ο��<��u�:� ��������� ͟�"Ø�G��pލ W��Ϻߑ�b���� �Ң���� U��XǞ U���J�� g���V���?Kx������>���� ��=�O�a�s߅ߗߩ� ���������1���9� K�]�o���l���� ������#�E��Y� k�D������������ �1CU;y �d/���
ߜ/�/�/�%2+|	??-???P=//h22c?�?�? �?�?�?�?�?
OO.O 5t,~ONz!��Y�Z� �ii	"��./0y@�O�O'__CV�� @^W�O�I�!�Wv3��>~��_@-����"#�U>L�P�Q"�BA)O<#�
��p�_�QR���PV�B�����uy�Uib��U@ 6��T}o@/�@�f��oh9[+B� �U�o4UgJ��P:`>�ad9_/_�^�CIt$ 	�$Z6K>�b
�;�A�D�;��]���jP+�{�̩�.������iQ$敕Ņ(4�$�х����;��=.��>��H	�iQ�5���8M�	Y%�qM=�PA�iR!R�x�	o���s����� �ן����"�4��o�IM!�F�   "��]b2d�b:`���� �J��bh����ѯ�e�(��讅B���cu�?333qU��rT�I��aD/  C�G�P ?fffqQ>Za�Duŕ����C( f�0͝Mq_k���u 7�I�j�]EO׿Qϫ�<��F@ ���Q��b�Dz������ϭ�k��!�/�) ܹ�˿ݿ����%� /����m���ߑ� �ߵ������������ 3�E�W�i�{����@�����2�����E� ����������%� +�R
�@Rd v��T��b� F*<N�FՖ/`\�6/H/Z/d��)� r ~�iX�/�.�_�C /?��a�p��r ae =2�dyavn`�E�i� j?��P�$r!X�E4�>9e�Z8i$m��oL<+O7H>���i$7J �/�/�/�/�/�/?�O )?;?M?_?�?/_�?�? �?�?�?�?�_O%O�_ IO[OmOO�O[o�O�O �o�O�O_!_O_E_ i_{_�_�_�_�o�_�_ �o]l4/f/�
��2�2��e�w�������	�Ă2������ �0�B�T�f�x����� �Ϋ��q�d!�!�|m� q�q�erz�`����D� V���z����d%����&�8�<��҃��>����}����~s��>LW�>�~o��y<'#�
%arp���p��N�������@�e�a-�Ų�`E�@�� F���ddu�bo$� m�
��b�o�{Bq.� *ϐϱ��Ϧ����Ϭk��>�j�����L�#��It$ e�$��>%�k�
Eߗ�A"����?߹�c�u�Ơ+��=��.����š�$敕!�(4$��-�����;��.�Y�>��He�š5���u�8M�Y��͝=>���Ţnq����	���������A� 3�H�Z�l�~�������|}��  qr �����9�����ݚ ��	-?��V�D���s��?333ͥΤ�E��D/  C�`GÿP ?fff͡> �����	�)o�x�� ����ͯ���ϓ ���e��3�/%zFF@ 9%E��FDz� Z$E7/�	/�X�8�*� � '9K]#?��/ M?_?��%o�/�/�/ ?'?5?g?%O7OXO�? �?�?�?�?�?�?OOO �O_�OgO!\��O/ y_'/9/K/]/o/�/�_ !�f_x_2o�_�_�_�_ �_�_�oo,o�oPo�o to�o�o�o�o�%��/0����(ȅO�p �cPɴ�j(�E��y r�IU�^�MR�p���� Z�ձy�ʰ=�=�zƏ wV���q�������M���t���u�����>����t��� ��+�=�O�a�:��� ������鏋���� '�9�K�$�o���Z��� ��ɟ۟�����#��� G�Y�k�}�����_�ů ׯ�����1�C�� g�����T�f�xߎՁ2������������ �2�D�V�h�z� ������������ �2�R�}	}
r��M�	 �	���O�G�������������Q�����P����B.�9�>6q�]��TRIR��j>�L� �ڿd���<#�
��a�pj	FU8��=���9�-� 1��!B��@�A� 5rM�����B����Jf ���Bb��� �///C/U/�� �>F������/�I�t$ �/$�>��
�/�'A~��/�/�?�/�&" +��̞a5.���m5!$�敕}5(4$�x�5A?S;;��.�5�>��H�5!5{���58M�Y�5)�=� �5!��
O0;	'?@O+OdOOG�?�O �O�O�O�O�O[��n>�G  ��Jp ��� YUAU9�FQ e_w_�_�_B�_�^�=��?p�-u?3�33)aR*m��D�/  CN�G�P_ ?fff)> n�-uMiEa����_�b M}U�)#gQy-/�o "���o	c�ʢ`F@ �u�a	eI�`Dz7`�t�o�ep#z�є߆� �qo �o�o�o�o��o��� ��%7��7�I�[�m� ����Ï��������� �!�3�E�W�i���Y�k��ß}����_կ �������} ¯ԯ����
��.�@� R��v���Ϭ���п ����P��uN���� �����*�6� �W�τޡk����� ��b���*��Ҷ 1�&���i�"�l� � i�*�Z��{���V�!�%?_������>���!���Q�c� u߇ߙ߽߫ߖ����� ��E���M�_�q�� ��������� %�7�Y�m��X�� ���������!3 EWiO��x/����߰/�/�/�%2@?|?/?A?S?d=C/|22w?�?�?�?�?�? �?OO0OBOIt@~cN �!��Y�Z�%�)i)i "2��B/Dy�O_;_2_WV�� rW�O�I(�!�W�3J>���_�T-����6#�U>L�`�Q6�BU)<#�	
��p�_eR��/dV�B��J���U}b��U@J��T�� �oT/-��f%��o|Mo+B��U�oH�i{^��dN`>��a"dM_C_��CItk$ �$n6>�#b	
�O�A�DO��q�x�-�~P+��̽��.���Ʌ}Q$�{��م(4$�兼����;��.�>���H�}Q5�=�-�8M�Y9��M�=�PU�}R&!f���	 ������������� ���$�6�H�W��$C�CSCH_GRP�14 2����y�&� �\m.2�p)  )"��qbFd�b N`֥���Jávh���@��y�/���B���y+c��?333�U�ޢ�T�I�aD/  �C�G�P ?fff�Q>na�D��ʹ ±�W(��D©ͱM�_ ���ɉl�~ϟ�qYO�φ�����F@� �����b�Dz ��3����Ϡ�1�/�) �� ��$� 6���Z�d�&�8�ϴ� ��������� ��@� ���1�h�z���� ������(�����g�@����z���R ��$� 6�H�Z�`�R?Q u������� �){M_q� �{ժ/��k/}/�/���^�� �y��C/ >�_�CR/K?"��p &� uer2t�a1v�` �E�i��?�`�$�!���z4�>Me&��8�$����oNL`OlH>����$lJ�/�/�/?? (?:?_^?p?�?�?�? d_�?�?�? OO$O�_ HOZO3o~O�O�O�O�O �o�O�O�o _2_D_V_ �_z_8�_�_�_�_�_ �o
oo�@o�li/�/-�?�Q�g�2�̚���H��Џ����2� �/�A�S�e�w����� �����Ľ����+tV� V�K|�������r���� ���y�������Ԧ*tZ��[�m�q����a>!6��}-"�sC�>L��s��o<=��y<#�
Za:r�pC��������au
qb���pz�@��{�"&���d ��oYƢ�?��b�o�{B;qc�_����������.��k˰>���ʯx����X�It$ ��-$�>���
z���AW���t��ߘߪ����+���:�.��y�F���$敕V�(4$�b��,�;���.��>��H�����5����8'M�Y���=s������q��	�	 ��� =�(�v�h�}����������4�ڝ���  �r# �ôn�˰ 2��>Pb�t��y�� <��%?333�:��F�z�D/  C�'pG�P ?fff�>�G�%& ^o�x���&-.��� *)�����e֟h��</Zz{F@ `n%z�"�{Dz �$zl/>/���m�_� �J\n�� X?��/�?�?�/Zo ?"?4?F?\?j?�?ZO lO�O�?�?�?�?OO 0OBO�O2_D_�O�OV\��O8/�_\/n/�/�/ �/�/�_V��_�_go�_ �_�_oo+o�oOoao �o�o�o�o�o�o�o)��%'��/����(ȺO�s�����]� z�H����~U����R ��΂��
�����r� r�Bz��Ew��B����@քT�ʵ���t���8Ϫ���Ș>��� �tȚ*�<�N�`�r��� ��o���̏ޏ����� &�8�J�\�n���Y��� ����ڟ����2�� F�X�1�|�������� ֯������0�B�(� f�x�Qߜ�������߭���2,����$,�=��U�2P�y� ������������	� �"$.<�gчĲ	�
 ���M��_�G߀)����0�����K������wc�#�>kq�-݉R~R��>L� �ϙ�.�<#�
����p��>{U��=r���#�b�f��Vw��@#Q�jr�-���R���J�U�&�H�B ����!/B/T/7/x/�/=�'>{�&��/��It$ �/$�G�>��
�/(7A���(?�/J?�/6W +���̖5.�����5V$敕�5(�4$ܾ5v?�;;�{�.�5>��H�5�V5��E8M�YE^�=� .EV��?Oe;	\?uO`O�O �G�?�O�O�O�O_!_�6�~3W  �pJ�'�U vUn�{QO�_�_�_�_PRB�_�^r��tpbu?333^�R_|���D/  C���G�P ?fff^>G��bu�iza�� 0�S_r�}��^Xg�y b/$6WJ�2��o>x����`F@ �u0�a>e~�`Dzl`�t��o��Xz���߻� ܦo�o�o�o�o�� �ޏ��Zl��l� ~�������Ə����ȟ � �2�D�V�h�z������������������ 2��
����� � �����	�ÿ-�?� Q�c�u���Aϫ���O� �3���)�;υ�3����I�#�5�G�Q�� �_�k��EW�Ϲ�� ��
��ڥNb�ޢ_� N*��f
&[��� ��W��� ��_�EZ2� ��&�VG�V�Z?�x��$�>���V� $��ߘߪ߼������� ���(�:�L�z��� �������� �� �6�H�Z�l���H�� ���������<2 �Vhz���� ��/�J!�S��/�/	?52t|R?d?v?�?�=x/�22�?�?�? �?OO/OAOSOeOwO ~tu~�N�!�ij, Z�^i^iR"g�M�w/yy@1_C_p_g_�V�0@�W_%Y)1�W�3>���_�-�ڢk#�U>LD`+ak�B�)O<#�
�p�_��Rץ;/�V�B�����e�b�2e@ �3d���o�/Qb�O@vZ��o���+B� e}�������`>�aWd�_x_9�^SIt$ R�$�6K>�Xb
2���AT���,���P�b��P+�{���.�����޲Q$敕�(4�$��ҏ�;��=.F�>��HR��Q�5��b�8M�	Yn��M=+`���R[!����	��џ������ .� �5�G�Y�k�}��o��MjΏ�   ^"���b{d&r�`�ҥ �Jס�h����,���(C�1��B���`c��?333�U�T�I�2qD/  C�G�P ?fff�Q>�a�D��޹ֱ�( ��y����M�_���ɾ �ϒϳϦ�O Ϛ���<*3�F@ &�2����b3�DzȰG�2��$��ϴ�E1%?9 ���&�8�J��n� x�:�L�������� �����"�T��$�E� |������������@<�����{�T���� ��f�&�8�J�\�n� tbSe��� �����= �as������/`��/�/�/���r� � �=y��W/>2o�C f/_?6��Kp:� �e �2Gt�afv�`*U*y� �?�C`�$�!���4N�e:��8�$���obL<tO�H>����$�J �/�/??*?<?N?'_ r?�?�?�?�?x_�?�? OO&O8Oo\OnOGo �O�O�O�O�O�o�O_ �o4_F_X_j_�_�_L �_�_�_�_�_�oo0o 	�To�l}/�/A�S�e�{�2�̮���ҏ���	��2�1�C�U� g�y���������ӟ�� �����?tj�j�_|�� �����r������ɍ� ��̯ï�>tn���o�����/���a>�#!J��}A6�sW��>L�����oQ��y<'#�
naNrpW���p3���*����a@uqv��/p��@�� ��"":���d��om� ��S�r�o �BOqw� s��������0�B��k߰>3���ޯԯ��l��It$ ��$��>%���
����Ak�������߾��+��=�N�.���Z���$敕j�(4$��v�.�@�;��.���>��H���5�����8M�Y���=������q���	�-��Q�<��� |�����������H��|���  �r 7 �״��߰F.&� 3�Rdv�
���*��, ��%?333�N�Z����D/  C;pGÿP ?fff�> ��[�%:2ro�x �:-B��>)�� �/u�|�P/nz�F@ �%��6Dz$�$��/�R/*����s� � ^p���l?��/ �?�?/$/no$?6?H? Z?p?~?�?nO�O�O�? �?�?O O2ODOVO�O F_X_�O�Oj\��OL/ �_p/�/�/�/�/�/�_ j��_�_{o�_�_	oo -o?o�ocouo�o�o �o�o�o�o=�%;�?0���	8��O� #s�����q���`�� ���U���R��� ����������Vz� Yw��V�����h�޵�����LϾ�Пܘ>����ܚ>� P�b�t���������Ώ ����2�ԯ:�L�^� p�����m���ʟ���  ��$�F� �Z�l�E� ������Ư��ꯨ��  �2�D�V�<�z���e� ������߯����Ձ2,,
��.�@�Q�0�i�2d������ ��������/�6$-. P�{ћ��	�
��] 
�_W/�1)����(D����_��P���ыw�7�>q��AݝR�R#ӳ>�L� �#ϭ�B�<#�
ʱ��p�R�U8��Q����7�v� z��j���@7Q� ~r�A�	�R��Z�i�:�\�B���� 5/V/h/K/�/�/Q�;�>�:0�/��I�t$ 
?$[�>�
�/<7A��<?�/�^??6k +��̞�5.����5j$�敕�5(4$�x�5�?�;;��.�5�>��H
Ej5{��E8M�Y&Er�=� BEj�SOy;	p?�OtO�O�G�?�O��O�O_#_5_D[�$�CCSCH_GR�P15 2����fQ&�� \Z�]�  ғp^3 �;�U�U���Qc�_��_�_ofBo
n����pvu?333�r�Rs���D/ � C��G�P ?fffr>[��vu �i�aοD؈_1r�}�� r�g�yv/Yk�^��F��os���pF�@ �uqse�pDz�` ����z������ ��o�o�o #�GQ��%�� �ʿ����ŏ׏��� -�����U�g�y��� ������ӟ�ïկT�-�笸g��?��� �#�5�G�M��,�>� ��b�t���������v� ����h�:�L�^� pϺ�h���~�X�j�|����K��Р��zW 0������?�8���b  ���b_��z& o����ʌ���� �� ��zZg���:f|���n?�;�M�Y�>�����Y��������� ��'� K�]�o�� ��Q����������� �5�G� k�}����� ��}�����1 Cqg%/���� ���	�/-V� ��?,?>?T52�|�?��?�?�?�=�/�22 �?
OO.O@OROdOvO �O�O�O�t�~�N�!$ CiCj8,���i�i�"�� ���/�yf_x_�_�_�V$G0�WH_ZY^1g
�3�>��#o�-�8��#0e>Ly``ax�*R�)<#�
G'"p0o�R�p/�VR�����Oe�b ge@��hd���/ ����Fv��,���+B(!PeL��� �	����`>q�d�_�_n�ESIt$ Z��$�6>��b
g���ADT��a�ۏ������P+���'�.����3��Q$敕C�(4$�O����;��.{�>��yH���Q5����O8M�Y���M=`` ���R�!П��	�� �*��c�U�j�|��������!�M��ħ  �"��b�d[r �`���J��h+�=�@O�a��x�f�R��y�c��?333�U�'��T3YgqD/  �C G�P ?fff�Q>�a4T��� �K�(䯮��]�_ �����������O�U���)�G*h�F@� [�g�ϵrh�Dz ��|�g�Y�+���z1Z?L9 �7�I�[�m� �E�ϭ�o������ G���!�3�I�W�� G�Y�z����������� ��/�q�1����C���%ߛI�[�m� ߑߣߩCb��T �����< N�r����� /��?�ߴ/�/�/��ȧ�� �ry֧�/ J>go1S�/�?k߲�p o� �e�2|t�a�v�` _U_y/*�?2'x`/4�!�֪�4AN�eo��8�$��%�L�O�H>����$�J?)?;?M?_? q?�?\_�?�?�?�?O �_O%O7OIO[OmOFo �O�O|o�O�O�O�O_ �o3_E_i_{_�_�_ �_�_��_�_oo/o Soeo>��o�l�/�/v�������2����H��*�	�B�2=� f�x���������ҟ� �����)�T�tt�� ���|�����r���� �
�¯ԯ����st��8�������d�P�q>X!��vk�s��>Lհ���o<���<#�
�a�r�p��+�h�*�_���qOuSq��C�dpõ@ĴW"o���d ���o������Br5�B�q�����/�A�$�e�w�*{�>h���x	��ߡ�It$ ��-$4�>��
���A����7�����D��+��̃�.��y���C�$敕��(4$ܫ�c�u�;���.��>��H���C�5����8'M�Y��K�=���C��q,�R�	I�b�M� ��q�������������}�#��   �rl 7�ķ�� {c[�h<ȇ����?���_��a <�O%?333K���L�����D/  C�ppG�P ?fffK�>4���O%og �o�@
"o-w�K�E s)O�/#/D/7u���+/�/�z�F@ `�%�+k��DzY �$��/�/E*ց���� ܓ���� �?�	?�?�?G/Y/�o Y?k?}?�?�?�?�?�O �O�OOO1OCOUOgO yO�O�O{_�__�O�\�_�/�_�/�/�/�/ �/�/o���_�_�oo ,o>oPoboto.�o�o <�o �o(r� 5p�6?�"�4�>8�_L�Xs��2��� ÿ������U;���R L�;����S���H��� �ɋzD��w԰��L�2
@�����4�C�G�������>��� C��s���������͏ ߏ����'�9�g�	� o���������ɟ��� ��ؿ#�5�G�Y�{�5� ����z�ůׯ���)� ���C�U�g�y���q� �������7��@��������2a,?�Q�c�$u��eߞ�2���� ������
��.�@�R� d�k$b.�������	�
 ��G]KK?�T_:Wd߀f)0]Ty����Д 	����l�>�q�v��R�RX��>L1X���w�<#�
����p����U(߆����l��ů����@lQ �r�v�>�OR�<��GZ���oϑ�B ��/j/�/�/�/�/�/��p>�Doe�&?��It$ ??$���>�E
?q7A���q??�?=?O6� +�����5.�����5�$敕�5(�4$�E�?�;;�{�.3E>��H?Eޟ5��OE8M�Y[E��=wE�HшO�;	�?�O�O�O �GO_"_4_F_X_j_���W~|W  K��p�h"p�U �U���Q��_�_ooP�B0on����pM�u?333��R�|��!D/  C���G�P ?fff�>����u�i�a� y؜_fr�}����g�y �/m���{��x��� pF@ �0q�e� pDz�`4�����z2��� ��o%7�� [e�'�9������� Ǐُ���A���� 2�i�{�������ß՟��)�ׯ�h�A���� {��S���%�7�I� [�a��@�R��v��� ������п����Ϙ� *�|�N�`�rτ���|���ߒ�l�~ߐߚ�� _��д�*)�WD�� ��S�L�#��b8 '��� �s�4$�S&�) �ʠ���0�ԨюZ{� ��o'f����?�xO�a�m�>����� m���������)�;� _�q�����e�� ������%��I�[� 4������������ ���!3EW�{ 9/������ �/A�jߜ�.?@?R?h52�|�?�?�?�?�=�/�22�?O0O BOTOfOxO�O�O�O�O �t�~�N1,$WiWjL, ���i�i�"�����/�y@z_�_�_�_�V+$[0@�W\_nYr1gC�>�7o�-.�#��#De>L�`ta�>R�)O<#�
[;"pDo��R ��/�VR����%!ce�b {e@ ȡ|d�'�/����@Zv��@���+B<! de`�����/���`> q�d�_�_��^YSIt$ ��$�6K>��b
{�͇AXT�͏u�����P+�{��;�.���G���Q$敕W�(4�$�c��-�;��=.��>��H���Q�5����8M�	Y��]=t`ӕ�R�!�
�	���>�)� w�i�~�������Ư5��M��ا   �"$��b�dor�`3�� Z ��h?�Q�c�u���(��z�R���c�?333e;�dGY�{qD/  C( G�P ?fffa>�aHT�'��_�( ����'�/]o��+�� ��������Oi���=�<[*|�F@ o�{��#r|�Dz���{��m�?��ʎ1n?`9 �K�]�oρϓ�Y�� �߃�����[�#� 5�G�]�k��[�m��� ����������1�C�@��3E����W��� 9߯]�o߁ߓߥ߷� �Wb��h��� ,�Pb�� �����*/��(?`���/�/�/��Ȼ� 0#�yꧠ/^>{oES �/�?�p�0�e �2�tq�v psUsyC* �?F'�`C41��4UN�e���8�$��9�L<�O�H>����$�J +?=?O?a?s?�?�?p_ �?�?�?�?O�_'O9O KO]OoO�OZo�O�O�o �O�O�O_3_�oG_Y_ 2}_�_�_�_�_�_� �_oo1oCo)goyo R��o�l�/�/������ą2���	��-�>�	�V�2Q�z����� ��ԟ���
��#� �=�h��t�����|�� ���r����֯ ���1��t��L����ʩ΁x�d�$q>�l!��.������>L�б��/�<'#�
�a�rp��?�p|�>�s���$q@cugq��W�xp׵@$ شk"��.��d�o�� ����Vr'I�B�q�� ��"�C�U�8�yߋ�>{(�>|���'���ߵ��It$ ��$H�>%���
��)�A��)����K����X�+��=̗�.�����W��$敕��(4$�ܿ�w��;��.���>��H��W�5����8M�Y�_�=а/�W� �@�f�	]�v�a���������������"1��$CCSCH_G�RP16 2����S&� \G�/J�  �� K�  ���(���o��P� ����S�	�s���u �c%?33�3_��`�����D/�  C�pG�P /?fff_�>H��� c%���o1�u"�- ��_�z�)c�F/X/y/�Ku3��`/�/�z�F@ �%�`��Dz�4��/�/z*8�ʏ�� ��� ��/�?4/>? OO |/�/�o�?�?�?�?�? �?O�O�O_BOTOfO xO�O�O�O�O_�_�_A__�\�T_�/,o�/ �/�/?"?4?:o��o +o�oOoaoso�o�o�o c�o�oqU'9 K]�U5��k?E�W�i�s8�8_���s�� g�ێ׿��,�%��U p�� b��O�L���g� �\�ϥ���zy��w� ����g
T�Ҟ'� i��x�[��(�:�F�>���x�F�����̏ ޏ�����8�J�\� n���>�����ȟڟ� ��׿"�4��X�j�|� ����j�į֯����� �0�^�T��x����� ������������l�@C�u���+�A�2�, t���������2����	��-�?�Q� c�u������$�.���� �00%�|]��t� �_oW�ߛ)Se����4��5G	K������>�q��pb�R��>Lf�M����<#�
4��p��U]߻����������<���T@�QU�r / ��sĄRq�3&|Z/������B�=9/�/�/@�/�/�/?�˥>��y��[?2It$� t?$��>�z
T?�7A1�?N?�?r?��6� +���E.���� E�$�=�0E(4$�<E�?�K;��.hE>���HtE�5����E8M�Y�E��=@M�E�}ѽO�;	�? �O�O_WPOB_W_i_�{_�_�_/���~�W  ���p�� H"�e�U���Q�o�*o<oNo�BeoSn�����p��u?333��b� 	T!D/ � C�G�P ?fff�>�!�u  y�a8Ϯ��_�r � ��g��/��������B��4�UpF�@ H�Tq�e�UpDz�`i�TF���zg�G�9� �$6H Zl2����\�n�� �4����� �6�D� v�4�F�g�����ԟ ���
��^�����v�0�������6�H� Z�l�~�����0u��� Aϫ���Ͽ��Ͽ� )�;���_ϱσϕϧ� ��߱��Ǐ�߳���ψȔ�����_)�W y�7�T�߁�X��b m \������i$��& �LL)����e� ���Z��.��\f������?/������>����Ԣ���(�:� L�^�p�I������ �� ��$�6�H�Z� 3~���i�������� � 2/Vhz ���n/���
 /@R+?v��� ��c?u?�?�52�|�?��?�?OM�//B2 *OSOeOwO�O�O�O�O �O�O�O�t�~^A1a$ �i�j�,ح�i�i�"� ˧�/�y�_�_�_�_
f`$�0%g�_�Y�1Qg
=C�>E�lo=c�8X��#ye>L�`�ax�sR9<#�
�p"pyobU��/fLR���<%@!�e0rQ �e@���dD�\? ����vتu/" /";Bq!�e���.� �R�d�+p>Uq�d� o�_���SIt$ ZЏ$!F>��b
���A�T���$�Ώ���1`+���p�.����|�0a$敕��(4$ܘ�P�b��;��.ĕ>��yHЕ0a5����O8M�Y�8]=�` �0b�!�?�	6�O� :�s�^�������ůׯ����j]���  �"Y�$r�d�r ph�P�HZU�)xt���@����,�����LR�N�y�c<�?3338e�p�9d|Y�qD/  �C] G�P ?fff8a>!q}T<�\� T��
8-���\�d]8o 2�`�<����1�$%_����rߐ*��F@� �հ��Xr��Dz F��԰Ϣ�t�2��1�?�9 ܀ϒϤ϶� �ώ����߸���4�F� �F�X�j�|����� ����������0�B� T�f�x���hz������n���ߤ߶� ��������b��� +=Oa/� �)/�/��// _/�]?#��/?!?+����90E#�y��/ �>�ozS�/�?�(��p �90(uB�t@q�v5p �U�yx*1O{'�`x491��D�N u��!H04�4�n�L�O�H>���04�J`?r?�?�?�? �?�?�_�?OO&OTO �_\OnO�O�O�O�O�o �O�O�o_"_4_F_h_ "|_�_g�_�_�_�_ oo�0oBoTofoxo ^�o�o���o$|�/-?��я���2N�,�>�HP�b�s�R���2�� ����ӟ���	��-� ?�Q�X�O�r����t� ��|48�8�,�A' Q�S���J�A�f��t쀁���������Yq>�!ȿc���E�յ>L��E<Ϣd�<#�
�a�r�pտt���s�����Yq�u�q���­p�@YĠ"��c�+t <)��4
�ϋr\~�B�q����W�xߊ�m�����s{]�>��1�\�xR���It$ ,�-$}�>�2�
�^�A�^���*�<捰�+�����.��y��匱$敕��(4$�����;���. �>��H�,���5��<�8'M�YH���=�d���5�u���	����� �������!3E�W��l�D.i  8�� ��U� �]� ����������������� <:Ø%?333������ة�D/  C��pG�P ?fff��>}�٤�%�� �of��S"�-����� �)��Z/l/�/�uh���t/�/�z F@ ` 5!t�� Dz� !4/�/�/�*���� ��� //$/ �?H/R?O&O�/�/�o �?�?�?�?�?�?.O�O �O_VOhOzO�O�O�O �O�O_�_�_U_._�\�h_�/@o�/ ??$? 6?H?No�-o?o�oco uo�o�o�o�ow�o�o �i;M_q��i5��?Y�k�}��8�L_���s�{1�� �֣@�9�e�%�b ����`�!Ԝ�@֑�� ��z���w�Ԅ��{
@h��\�}��������<�N�Z�>��� ��Z���Ώ����� (��L�^�p�����R� ��ʟܟ� ���6� H�!�l�~�����į~� د���� �2�D�r� h�&ߌ�����¿Կ�� ��
���.π�W����-�?�U�2�,����$��������2��� �/�A�S�e�w����� ���$�.�����DD 9ܐ]���ҝ_�W�߀�)gy�����H��I[	_�	����>�q$��bb��1>Lza��+���<#�
H�(�p�1�eq����������P�	�h@�Qi�r/�߇ĘR���G&�Z-/�¸���B )�QM/�/�/�/�/
??�˹>!����o?FIt$ �?$���>��
h?�7A�E�?b?�?�?�6� +����(E.����4E�$敕DE(�4$�PEOK;�{�.|E>��H�E��5���E8M�Y�E��=a�E����O�;	�?_�O+_ WdOV_k_}_�_�_�_�"/���~�W  �����\"� e e 
a�,o>oPoboP�Byogn����u?333�(b�|4	h!D/  C��G�P ?fff�>�5�uyqL� ���_�r���g� �/�������V�x*�H�ipF@ \�0hq�e"ipDz�`}��hZ�,��z{�[�M� �8J\n�F� ���p�����H��� �"�4�J�X���H�Z� {���ğ֟������0�r� �2�����D�� į&���J�\�n����� ����D����UϿ�ѿ �������=�O��� s��ϗϩϻ����Ņ��ۏ�������� ������s)�W��K�h 2�ߕ�l��b� p��� ���}$��&�``) 0���3�y0����Z�� B��pf�����?&/x������>����� ���*�<�N�`�r�� ]���������� &�8�J�\�n�G���� }�������� �4 F/j|���� �/��0/T f??������w?�?�?�52��?�?OO+M
?CB2>OgOyO �O�O�O�O�O�O�O	_ ��*^U1u$�i�j�, ��i�i�"��ߧ	?�@�_�_o�_ft$�0@9g�_�Y�1egQC!>Yрo=w�l��#�e>L�`�a��R9O<#�
��"p�o�,bi��/+f`R���!P%T!�eDre �e@ ��dX�p?����@�v쪉C"/6;B�! �e��0�B�%�f�x�++p>iq�do
oˏ^�SIt$ �$5FK>��b
ď�A�T����8���E`+�{�̄�.������Da$敕��(4�$ܬ�d�v�;��=.ؕ>��H�Da�5����8M�	Y �L]=�`�Db�!-�S�	J�c�N���r� ����ǯٯ�������$CCSCH_�GRP17 2����@�?&� \4>��>79  �"m� 8rt�rp����\Z�� =x����Ϳ߿@�����`R�b��cP�?3�33Le��Md�Y�qD�/  Cq G�P_ ?fffLa>5q �TPՑɉ��8b�� p�x]Log�t�P�3�E� f�8% _��Mߧߤ*��F@ ����M�lr��Dz{������ߩ�pg��1�?�9 ܵ� ����������!�+��� ��i�{ߤ{���� �����������/�A� S�e�w�����������.��A�� ���������!�'�b �<N`r� �P/��^/�B// &/8/J/�/B�q?X�2?D?V?`��%n0z# �yT�
?�>�o�S?O �]��p�n0<u9B�t Tq�vIp�U�y�*fO�' �`�4n1T�AD�Nu�VHe4H��\'_3X>���e43Z�?�? �?�?�?�?O�_%O7O IO[O�O+o�O�O�O�O �O�O�o_!_�oE_W_ i_{_�_W�_�_��_ �_ooKoAo�eowo �o�o�o��o�o���Y|0?b?���.�2@��a�s�����������2�������,� >�P�b�t����Ԅާ� ҁ�t���im�m� a�v\����@�R��v����t!���"�4�(8��Γ�q>�!�������z�
�>L�S�:�z���<#�	
!q�p
ϩ��J���ݢ���q�u�q)����pA�@�B��" �Ϙ�`tq^ �i
��r���B�*�&ߌ߀�߿ߢ����ߨ{��>���fđ���H��Itk$ a�$��>�g�	
A��A���;��x_�q�°+�����.������$�{���(4$�)������;��.U�>���Ha���5�=�q�8M�Y}�ɭ�=:�����j�����	 ��������=�/D�Vhz���$C�CSCH_GRP�18 2�����&� �\��v/��  m�� ��5� ��٪��&8@J\��saݢ�� yo��%?333ɵ�"ʴ�A�D/  �C�pG�P ?fffɱ>����%) !%����"�-��ɿ ��)�߰/�/�/�u���P/�/$?!�c F@� V5b!���c Dz �w4b/T?&?�*T�4�&� �2/D/V/h/ z/@O�/�?jO|O�/�/ !�?
OO.ODORO�O B_T_u_�O�O�O�O�O __*_l_o,o�_�_>l��_ ?�oD?V?h? z?�?�?�oo�oO �o�o�o�o�7 I�m����� ��5��?����ӏ�8Ȣ_��sL���� E�A������fe�Z� jb뀹Ŷ�V���u��� 9�9�*��-�R�*�끀�
��<���jӘ�����ϒ�����>���ℰ��$�6�H�Z� l�~�W�����Ɵ؟� ��� �2�D�V�h�A� ����w�¯ԯ���� ��.�@��d�v����� ȿ��|������*� �N�`�9���̭�ߏq����2 <����H��%��=�28� a�s������������� ��
4>$O�oԚ ����]�����_�W �9����n���3��	��_K��>S�z�qbfb�Ӈ>L����<��<#�
��~ҁp�&ce��%Z���J�NѦ>"_��@a�R�j/��� �R�ϝ&�Z�/=��0�Bѧ�/	?*?<??`?r?%� >c!�x�?�It$ �?-$/�>��
�?GA�O�?2O�?�6?�+���~E.��y��E>$敕�E�(4$ܦE^OpK;���.�E>��H��E>5���E8'M�Y�EF=�U>��'_MK	DO]_H_ �_lW�O�_�_�_�_�_�	ok�$CCSC�H_GRP19 �2���:a�&� \�.��1�   ��g�2"$�" �ee V
�a7(�o�o�o�o:R(�o�nZ�\��J�?333F�bG�	��!D/  Ck�G�P ?fffF>/!�J��y�q��� \o�j�rFawn�J? -�?�`�2��G���<���pF@ Ӆ�qGuf"�pDzup���я��a����� ܯ������� %����c�u���u��� ������ϟ���ѯ� )�;�M�_�q�������@鯗���(�����;� �����ӏ���	�� !Ϛ ����6�H�Z� l�~ϐ�Jߴ���X��� <�� �2�Dߎ�<�k�`R�,�>�P�Z��� h�t��)Ng���� ���Wr� �h�6% 3��$N!�&C ��)�� `������h�Nj;���%�fP�_�BO|/<!->���_�-
 ������������� �1�C�U���%���� ���������	� ?Qcu�Q/�� �/��E;�/ _q����/�� �?/S,*�\��? OO(E2}�[OmOO�O�M	�?�B2�O�O�O_ _&_8_J_\_n_�_�� ~��^�1�$yz<c� gygy[2p�V��?��:o Loyopo�f�$@�g�o.i2A�g�C�!>����o�=��t3u�>LMp4qt/�R�9<'#�
!�"p�bp�D?�f�R���!@�%�!#u�r� ;u@�� <t����?Z$k�X/� c� ��"�/�;B�!$u  ���������ݏ+�p>�q`t�o�oB�c�It$ [�$�F>%�ar
;���Ad���5���Y�k��`+��=���.�����a�$敕�(4$��#�۟�;��.�O�>��H[��a5���k�8M�Yw��]=4p���bd1��ʛ	��گů���7��)�>�P�b�t�������$CCSCH_G�RP1A 2������&� \�>p߮9  g2�Яr �t/��p����Z��x  �2�D�VϷ�m�[��R����is��?33�3�e��di;�D/�  C� G�P /?fff�a>�qd ��� �/�8ٿ���� �]�o����Ǐ�߼��߀�%�_J����:]�F@ P�\����r]�Dz��q�\�N� ���8NA.O I �,�>� P�b�t�:��ߢ�d�v� ����/����(�>� L�~�<No������ ���� $f&�~8���>� P�b�t���r} �I/�����/ �/1/C/�/g/�/�/�/ �/�/?���?��?�?�?��Ȝ�0�#F� ˷�??N;c�?�O` ��T�d�0�u�BP��q o��p3e3�$:�O'7Lp $D�1˺�D6^�ud��H��4����\�_�X>����4�ZOO0O BOTOfOxOQo�O�O�O �O _�o__,_>_P_ b_;�_�_q�_�_�_ �_o�(o:o�^opo �o�o�o�ov��o�o  $
�HZ3�~�|@�?�?k�}�����2�� ؟�������7�22�[�m�������� ǯٯ�������I� i��ɔʉ������؂ �����ٷ�ɿ����h���-Ǚ�����Y�E��>M1t��pk`��>L�����{��<#�
�qx�p�� �]���T����D�H���8�Y���@��L2d� ��t�����
}�7��*�By��ŝ��$�@6��Z�l��	�>]��������It$� ��$)�>���
��
�A��
���,�����9�+���x�.������8�$�=���(4$ܠ�X��j�;��.��>���H��8�5�����8M�Y��@�=@��8��!G�	>� WB{f���������$CC�SCH_GRP1�B 2����4&� �\(��/+�  �a0,�Ԭ�	� �yP�~1؝����4��T��V0<��D5?333@ř�AĄ���D/  C�e�G�P ?fff@�>)х�D5�)}! ��V�"d=l�@�[' h9D�'?9?Z?,���/�A?�?��� F@ `�5�!A%`�� Dzo  �4�/�?�?[:ˑ���� ܩ/�/�/�/�/ �O?O�O�O]?o?� oO�O�O�O�O�O�O�_ �_�_#_5_G_Y_k_}_ �_�_�_�o�o"o�_�l�5o�?�?�?�?�? OO���o�0 BTfx�D��� R��6���,�>����6Ee�LO&�8�J�TH�ob�n���H���� �ς����eQ"���b b�0�-���H���=а� �١�Z�������b�H@5�����J�Y�<��v�	��'�>��� Y�'���������џ� ��ο�+�=�O�}�� ��������ͯ߯��� ���9�K�]�o���K� ������ۿ����?� 5���Y�k�}Ϗϡχ� ���ϰ���M�$�V������"�2w<U�g�y�$����{��2���� ���� 2DVh z�4x>�����)* �]ma)a)U�joPgz�|94Fsj�����(,������>ʁ����b�bn��>LG .!n�����<#�
���p����e>����������%�"��5%@�a6$ɂ�/��T�eb�R�6]j�/�҅ߧ�B ��%?�?�?�?�?�?�?�ۆ >�!Z$�{�<OIt$ UO$���>�["
5O�GA��O/O�OSOeF�+�����E.����U�$敕U(�4$�U�O�K;�{�.IU>��HUU޵5��eU8M�YqU�=. �U�^�_�K	�O�_�_�_ �W1_#o8oJo\ono�o��k�$CCSCH�_GRP1C 2�����a&� \��|j���  a� ހ�"~$)2� u�e�
 �a�(,>P�Rg�U~��Ӏc#��?333�r�51�D/  C��GÿP ?fff�> �!����qߏ��o |�����w��?�� ��׏�ՑD�����W�F@ J�V��u�"W�Dz�pk�V�H���؊H�(�� � &�8�J�\�n�4����� ^�p�ڏ������ "�8�F�x�6�H�i��� ��į֯�����`� � ϟ�x�2̸��� ��8�J�\�n������� "wω�C߭Ͽ����� �����+�=���a߳� �ߗߩ߻�ﳕ��ɟ0�����јȖ��� ��@9�g{�9�5/��� ��Z��rN0^���%�� J4�!i6� --9��� !�F ����j��0�%^v�����O�/���>�����
� �*�<�N�`�r�K�� ���������& 8J\5/��k/� ����/"4? Xj|���p?� ��//?B/T/-O x/�,����eOwO�O�E�2��O�O�O_]�?1R2,_U_g_y_�_ �_�_�_�_�_�_���� nCAc4�y�z�<ڽ�y �y�2�ͷ�?���o�o�o�ovb4�@'w�oP�i�ASw?S�!>G��n	Me�Z��3{u>�L�p�q�/ub
I<#�
�!r2p{rW�8�?vNb���!>5 B1�u2�S0�u@���t F�^�	O�$��/��ںw�12?$KBs1�u�� ���0��T�f�;��>W��t�o���cI�t$ ҟ$#V>��r
���A�d����&�П�3p+��̞r�.���~�2q$�敕��(4$�x��R�d�;��.ƥ�>��Hҥ2q5{���8M�Y�:m=�p
�2r�1�A�	8�Q�<�u�`��������ǿٿ�����$�CCSCH_GR�P1D 2����.�&�� \"N��%I  �2[�&��t �����s�Jjx�+��π�ϻ���.�����Nb��P��s>�?333�:u��;t~i��D/ � C_0G�P ?fff:q>#�d>� �wі/HP���^�fm :U�b�>�!�3�T�&5�o��;��:��F�@ ����;�Z���Dzi��������U��A�O�I ܣߵ��� ���߱�������W� i�/i�{��������� �����/AS ew��������/��/���� �������/�r�/ �/*/</N/`/r/�/>? �/�/L?�/0???&? 8?�?0�_OF� O2ODON��\@h3��B� �?�N�|cO _�K� ˀ�\@*�'RǄB�� 7��e���:T_�7�p�D \AB�/T�^���DXSD�6�p�lo!h>���SD!j�O�O�O�O �O�O�O�o_%_7_I_ w__�_�_�_�_�_ ��_o�3oEoWoio �oE��o�o���o�o�o 9/�Sew� ��������G�O PO�����2q�O��a�s�����u���2 ��ү�����,�>� P�b�t�{�r���� �� �W[�[�O�d Jt�v�.�@�m�dω�߄����"�&���
��|�>�1�φ��8�h���>LA�(�xh�򲇙<#�
��p�ϗ��8���˲��|�����կ�Ѐ/�@|0��2�߆� N�_L��W�߮����B����z��� �������>��T���u�6��It$ ZO�$��>�U�
/���Aā�)���M�_�ް�+�����.��������$敕(4$������;��.C>��yHO��5��_O8M�Yk��=(� ���X����	��� ���+2DV�hz��$CCS�CH_GRP1E 2�����&� �\��d?��  [��0��x�#��% �Ǻ���/&/8/J/P�a/O.˲��0]��5?333��"��|��/�D/  C܀�G�P ?fff��>�����5�)�!� ���v2�=㽷��'�9 ��?�?�?����>?�?xO�Q0F@ DE0P1�%��Q0Dz� eD�P?BOO�:B�"�� � ?2?D?V?h?._ �?�OX_j_�?�?��O �O
__2_@_r_0oBo co�_�_�_�_�_�_o�oZo�oro,|� �oO�2ODOVOhOzO �O��q�=��� ������%�7�ɏ [�������������E�ܟ�O�������H� �oِ�:�u�3�/� ����}�Tu�"H�Xrِ �դ�D��c��'�'� �ѯ�@��ّ��� *��X&��Д����x������>���Д �� ��$�6�H�Z�l� Eϐ�����Ư������ � �2�D�V�/�z��� e߰�¿Կ����� .��R�d�vψ϶Ϭ� j�����������<� N�'�r��ܛ�͟_�q�����2�<��������+2&Oa s������� �4�>=�]�)�*}� �m�)�)���o�g���9@����&\���@!'����M'9��>A�h/�_rTr��u%>L� �!��o�O<#�
��l�pu/�"Qu��&H�����8�<�%,2M�%@ �a�$@�X?����b��@�6�jq?+����Bm� �%�?�?O*OONO`O�� >Q1�$���O^�It$ �O$K>��"
�O�GA���O�O _�O�F- +�{��lU.���xU�,!$敕�U(4�$ܔUL_^[;��=.�U>��H�U,!�5���U8M�	Y�U4=� e,"��o;[	2_Ko6oooZg �_�o�o�o�o�o�o{��$CCSCH_�GRP1F 2����(q?&� \��>�  ��U�  2�$�2� �umuDrq %8����(b��~�H�J��#8�?3�334%�r5$x�1D�/  CY�G�P_ ?fff4!>1 y8�y�q����J� X�`4/O�\�8O�-� N� ���5�����΀F@ ��́5�T2΀Dzc��͏����pO������ ܝ� ����ӏ叫�	��կ �Q�c���c�u����� ����ﯭ�����)� ;�M�_�q�����׿�����￩̸)ϋ�� ����ӟ���	�߈" �� ߺ�$�6�H�Z�l� ~�8�ߴ�F���*��� � �2�|�*�Y�@��,�>�H���V�b� �9<w����/v��� ��E��0��V�$5!�4 <1�610��9��N�� � ��V�<z)��%�v>M�0_j?�>���M�}��� ����������� 1Cq/y��� ���/�	�/-? Qc�??���?� ��/3/)/�?M/_/ q/�/�/{?�/�/�O�/�A<�J��O�O _U2@k�I_[_m__�]oO�R2�_�_�_�_oo &o8oJo\onou�l��n �A�4���<Q�U�U� IB^�D�nOp�(:g^�v�4	P�w
y( Q�w�Sv1>�����M����bC�u>L�;�"�b?�b�I<#�	
	1�2p��r��2O�v�b��v1�5�1����0)�@v�*��� Տ�OH4Y�F?�Q���2y?�KB�1��t��������˟ݟ�;z�>�΁N�yo0�sItk$ I�$�V>�O�	
)�{�At{�#���xG�Y��p+�����.������q$�{���(4$���ɯ۫;��.=�>���HI��q5�=�Y�8M�Ye��m�="����rRA����	 ��ȿ���׷%��,��>�P�b�tσ��$C�CSCH_GRP�1G 2������&� �\�N^�I  UB����r�� z�����j����� �@2�Dߥ�[�I��b���yW���?333�u�
Ҳt�i)�D/  �C�0G�P ?fff�q>���d���� ��?�H��p����m� ���鵟�����5�o�8���	JK�F@� >�J��тK�Dz ��_�J�<����<Q_Y ��,�>�P� b�(���Rd���� 	?����,:l *<]����� � T//�l&,���~/,�>�P� b�t����/�k/}/7? �/�/�/�/�/�/�?? 1?�?U?�?y?�?�?�? �?���O���O�O�O��Ȋ�@�34���oO -^)��c~Ow_N%��B� R"�@���R>���]��� !u!�J�_G:�T�A��ʦT$ny�RֻX�D୯�zl�o�h>����D�j�O__0_B_ T_f_?�_�_�_�_�_ ��_oo,o>oPo)� to�o_��o�o�o�o ��(�L^p� ��d���� �� ��6�H�!�l����O�OY�k�}���2��ƯدH�����%�2 � I�[�m��������ǿ ٿ������7�W��� ��w������ƒ�� ���Ϸ����� �V���ׇϙɝ�G�3��>;Ab���Y"N"ߓo�>L�П�ߏ<i���<#�
��f��po��K%���B����2�6���&�G���@���:BR���ń �Ï���k�%����Bg��Ջ����$��H�Z����>K�����x�ϭ���It$ ��-$�>���
����A����������'��+���f.��y�r&�$敕��(4$܎FX;���.�>��H��&�5���8'M�Y�.�=���&�ϑ5	,E0 iT�������� +�$CCSC�H_GRP1H �2���"!�&� \���?�   ҒO@��Ԛ���%g% >�l!�/�/�/�/"(�/�.B��D@��2E?333.Շ"/�rɾ��D/  CS�G�P ?fff.�>�s�2Es9k1�� � D/�2RMZ�.�I7VI2� O'OHO�ϵ?/O�O<���0F@ �E�1/5N��0Dz]0�D�?��O�OIJ������ ܗ?�?�?�?�?�_O _�_�_KO]O��]_o_ �_�_�_�_�_�o�o�o o#o5oGoYoko}o�o@�o��o�|�# �O��O�O�O�O�O_ 	��������0�B� T�f�x�2�����@�ҏ $�����,�v�$US�`:_�&�8�BX� P�\���6'쟪���p� �����u?2���rP�� ���6���+��Ş鏚 H����Џ�P�6*#������&8�G�*d���<	��>���G�� w���������ѯ㯼� ��+�=�k��s��� ������Ϳ������ '�9�K�]��9�ϥ� ~���������-�#��� G�Y�k�}ߏ�u���� ����;��D�������2eLCUgy�	i��2���� � 2DVhoD fN������)�*��K} O9O9C�X>wh�jI"/ 4/a/X/}&�� �'�/)�'�p�>����/z��r�r\��%�>L501\��{�<'#�
���p�/�"p�u,��&���p�@���5�2��#5@pq $4���?z�B�Sr@�F Kz�?��s��B��5 OnO�O�O�O�O�O��t0>�1H4s/i/*_#�It$ C_$�>%�I2
#_uWA $u_�_�_A_SV� +��=��U.����U�!�$敕�U(4$��e�_�[;��.�7e>��HCe�!5���Se8M�Y_e�=0{e�"L�o�[	�_�o�o�o�go�&8J\n}{��$CCSCH_G�RP1I 2�����q&� \��X���  O�̐�2 l4Bt0�u�u��q�8 ��,�>��bU�C������Q3��?33�3�%��$�#AD/�  C��G�P /?fff�!>�1� ������}��j�ϝ ��/Ƈә�O����ş���2�����E�F@ 8�D����2E�DzڀY�D�6��ƚ86	 ��&� 8�J�\�"�����L�^� ȟڟ�گ����&� 4�f�$�6�Wώ����� Ŀֿ����N������f� ܸ���x�&� 8�J�\�n������"e� w�1�߭߿������� ���+��O��s�� ����������������Ȅ�����.I �wi�'#?�x�qH� ��<@L���5�8D�1 WF�0%I���40 ��z�s5L������_�?t��>�������� *<N`9/��� ���/�&8 J#?n�Y?��� ���?/"/�?F/X/ j/|/�/�/^O�/�/�/ �/?�?0?B?_f?�<@����S_e_w_�U2� �_�_�_�_m�Ob2oCoUogoyo�o�o �o�o�o�o��~1Q QD|�|�qL��̉̉�B �ϻ��O癟����vPD�P���y�QA�-c�1>5�\��MpS�H��Ci�>L����?cr�I<#�
�1`Bpi��EթO�<r���1,E0A�� �A@��@����4�L� �O�4�½?���e�B�?[BaA������@��B�T�K�>E��ń����~sIt$� ��$f>�Ƃ
���A}t򯚯����Ц!�+���`�.����l� �$�=�|�(4$܈�@��R�;��.��>���H�� �5���е8M�Yܵ(}=@���� ��A	�/�	&� ?�*�c�Nǜ��ϣϵ�����������$CC�SCH_GRP1�J 2�����&� �\^��Y  �BI��鄔�� y�a�8zf���ߗߩߠ�������<r�>�<΃,�?333(����)�ly��D/  C�M@G�P ?fff(�>�mt,�m�e� �?�H>���L�T}(�C� P�,��!�B�E�o���)����J��F@ `����)�H���DzW� �������C��Q�_�Y ܑ������� �����E�W��? Wi{����� ��/ASe w��y/�/
/��,�/��/�������� ����?|��/�/�?? *?<?N?`?r?,O�?�? :O�?O�?OO&OpO�M_4_ _2_<�/JPVC��0��O�^ ��js�O�_�%9⹐�" JP�b��0�Ԗ%��u ���JBo�G���TJQ0�@d�n����2hAT$��^��lx>��� ATzq_�_�_�_�_�_ �_�oo%o7oeo� moo�o�o�o�o���o �o֏!3EWy3� ��x�����'� �۟A�S�e�w���o� �������5�_>_Я���
�2_�=�O�a�$s���c���2���� ҿ�����,�>�P� b�i�`��ή�Δ���� �E-I�I�=�R/8'b��d��.�[�R�w�͔����������ת�j�>�A��t��"�"V���>L/��V��u�<#�
��ݒp��߅��%&��ֹ���j������⾐�@j!�B��t�<�M"�:���E*�m���B ޑ��h�����~�������n�>��B�m�c߼$��It$ =$���>�C�
oA���o�;M��+�����.�������$敕�(�4$���;�{�.1>��H=ޝ�5��M8M�YY��=�u��F���	���� �/ /2/D/V/h/�w+�$CCSCH�_GRP1K 2�����!&� \��|RO��  I� �@��f��n��%�%�� �!��??&?8?�O?�=>����@K�E?333���"������D/  CʐGÿP ?fff��> ���ĩE�9�1�w��/ dB�M�ͥ��7�I���O �O�O��y�,O�O _��?@F@ 2U>A�5��?@Dz�0ST>O0_�_�J0��� � O O2ODOVOozO�_ FoXo�O�O���_�_�_ 
o o.o`o0Q�o �o�o�o�o�o�oH ���`����O r� _2_D_V_h_z_�� ��_�q�+�������ˏ ݏ��%���I��� m������ퟛUʯ�_0�������X�~Ǡ ӓ(��'c�!����r� k�B��26�F�Ǡ�咲 2���Q�������� 	�.��ǡ�*���m�F6�������ǹ���>��������  ��$�6�H�Z�3�~� ������⿄�����  �2�D��h�z�S�� �������ϰ�
���� @�R�d�vߤߚ�X��� ���������*�<� `�쉯��M_q��2�L������2=Oas �������D�N  .+K�v9v:k��}�9 �9����w���I�/�/�/�/�&J�z 7{/P�)�;7'��>/��V?��M�B���c5>�L�0�1��]"��<#�
z�Z�pc?2?�8��66"����&� *�5B;�5@�q�4 .�FO�����r��yF�z_O���B[�5O �O__�O<_N_��0�>?A�4�/�/�_x#I�t$ �_$>��2
�_�WAw$�_�_�o�_�V0+��̞Ze.���fe1$�敕ve(4$�x�e:oLk;��.�e�>��H�e15{���e8M�Y�e"-=�0�e2��)k	 o9$]Hw�o� �����$[