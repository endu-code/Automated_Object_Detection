��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER� q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS�	 DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� �ERE-   � �0�B{!F S{T� M�DTR>S$STD6XlQCWFA� 7X�QCW�"�YV�"eS/ �A7  � $�@TINvd@�0SUL� ��R_@ 3 $}@ SW@��RO�RR%	 ��P�T� �@JUx� �SqFS4D6'
 �2P�0_@c�FOL[d!$FCIL� jjE�P��C�S�aDIG4RC�_SCA��cI�NTTHRS_�BIdA�dSMAL��bCOL�bG��`� �� ��_�IVTIM�$t!0B"$S?0~xCCBDDN���-qI2wT2wDEByUdA\!SCHN�"TOfa0�! � Q0 mr<0V� �;!�r�AUTTUNN� TRQa�uE40�N �qFS3AXG  � 1eb}t�r5I�v	"G_gr7 l �!�3@�WEIGH�q�2 UuS_5QF(�T2��WA� 	pEsNTERVA�; - Q��� S!�t�AS0S�{$J-_STA�p� JQg���1(�*��2��3��W���� hqx��"COG_�X�Y�Z�ҁCM�p?�p�܂RSLT�4��D�P�D��	"_�p_�q�7  �~�b#0V�ROUNDCMVP�ERIODA�1P�UU3F2D�'TM01� �Ƒ_D���GAMMc1�TWRXI�K�K�MK��CLbP�&O00�ADJ�GAu�U�PDB�A:p%0/ ,$M"P30f��� d�:pG �p"��HCD�G]V�#GVY��Z�GJDO5�,q��S��7$R��E_8@{t٣�pAPHBCy��$VF6��P��2L��蘨@IL [����;���;�d@���RG���NEW_���r�Q}���ڡN�5OBOA@fY�sW2/�G<�	����ȴ�\�2�E�KP�NUC?NPRGOV��Ŝ�@`d_TW�c,�G�E^!NV2#C�c0�@�WTS�TRL�_SKI2!$SiJ�Q��NQpGW���	"��7 \ m;0FR]b� � CMDC���T�b���TO?��� �5گ���_�Ah 0 '�>�ALARM�_��*�TOT6�FRZn l�,!Y 3��X!�� mӥ�X �Œ`X �ʕ�U#��2��2
�X#Z�N��FIX�8��F�"d��IT�`IB�PN_d��CH�%���_DFL _�BF2N�ڶ�3����� ��3�"�����ʷ�(� ����3��3
��X��DIA����/#� ���%��� ��[1��g1�[���Z���#��!���%����$0�@
p��7F��D,�� HA�pU�5����v�FSIW6K �2PN@�`R>!��PHMP�`HCK%���>0G�'*#eb A����pNT��p^H	��HUFRzs�3��A��UgvCa��$v0Q ��i��@p@p � � SI0��  �5�I�RTU_��� %S�V 2���  � �6>0]@�]	Q�EF@� �oP�  ��  � �/@/'/9/K/U%@pd@p
m hK�/w/�/�/ �(��$��/� �/�/ ?.8e"�/?J?\?r? 8?�?|?�?�?�?�?�? �?>O4ObOO�OTO�O �OjO|O�O�O�O_�O (__\_f_�_B_�_�_ �_�_ o�_$o�_Ho>o o^b�/�ot��%�/�o��o�k	MC:� 5678  A�fsdt1 78901234qx#5w  	q 6xz.Ops�3'��j l�o�o����������,�5�DMM c�)5�A ���x�������=���O�R 2	Q� "��m��_� tu�B?)D�N�S4D 
FQ�!tY�d�!Ls`|�q`rƈ̀?�l��B𴐠�$ ON�FIG �}(�[ � ������i!�� 2��,
Hand guide���?�3��� � �X��с��ь��g#�=���A��ύ�������p �ݯ�(��L�7�p�x[����m*�� ����ʿܿ� ��$� 6�H�Z�lɌ��ό��� ���������
�C�E�]I 2Q�(�0� -�zՀ�F�M���_`πB��<��d�C�  ��uq�=#�
_aNnk=(��K����̥�@��e��=D�y���_a;�����8I��_aIt�$ �$F�>�s��k"���Q�Fۀ3]儢ѯǯ����!�/�``+��=���.�����_a�$敕��(4$������>�E���B<~w%�_a8�E�y5�;�j�A��Ҝ�Q�>��]�_a?��m���஑����~u1�?�3�3����0�:�o ����0�����LSB��~uq�ӻ���m�S]���/8��� ��� t�	eF|���P]��߯���x�n��;�.��z��3�'	���,��B���4*� 2/V��%D�DGH  *%v�+� �^-��
�/��/u/F~u�J/l/�)AI��/�/�?/ A��n5��p��4vO?�;)�7�?�?�o�?�8J�hq�?�?zyjG�_F?SIW Q��9 ��O�O�Ou�