��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGDsEV��RCM+ ;$Z <��QSIZ�X|�� TATUSW�MAILSERV~ $PLAN� �<$LIN<�$CLU���<${TO�P$CC�&sFR�&�JEC�!}�%ENB � �ALARl!B�TQP�3�V8 S��_$VAR9M �ON
6��
6APPL
6PA� 5B 	7'POR��#_�!�"�ALERT�&�2U�RL }�3A�TTAC��0ER�R_THRO�3UaS�9z!�800CH- �Y�4MAXNS_�1�AMOD4�AI� $B� �(APWD  �� LA �0�ND�ATRYQFDEL�A_C@y'>AERS�I�A�'ROtIC�LK�HMR0�'� X�ML+ :3SGFReM�3T� XOU�3�PING_�_COAPA1�Fe3�A�'C�25�B_AU�� k �6R,2COU�!H!U�MMY1RW2?��RDM*� $�DISc �SMeB�	"�BCJ@b"CI2AIP�6EXPS�!�P�AR��TCL��
 <(C�0�S�PTM�E� PWR���X�X�Qo !l5��!�"%�7�I�CC�%� kfR��0leP� _DLV���YNo3 �<oNbX_�P~#Z_�INDE
C�`OFYF� ~UR�iD���c�   ts �!�`MON�r%sD�&rHOU�#�EWA,vSq;vSqJvL�OCA� Y$Nޅ0H_HE����@I"/ 3 $GARPz&�1F�#W_\ �I!F�`;�FA�Dk01#�HO�_� INFO�sEL	% P K � !k0WO` �$ACCE� L�VZk�2H#IC�E�L�  �$<�s# ���k���%
��
`�K`SQi�w��5|�I�0ALh�z�'0 ��
���F��]����܅�$� 2ċ$b�w��@����� č��!r��Z���4���Ċ!�147.87.?224.20h�S���96����܁܁�3�_{p_  �ċ� bfh.ch̟�1�C�U�g� y���������ӯ^�� _FLTR  ���π �����B���n�nxč2n���rSH�PD 1�ĉ  P!
�robstatison֯՚!k�.�Q�ſ������� �޿?��c�&χ�J� �Ͻπ��Ϥ����)� ��M��"߃�Fߧ�j� �ߎ��߲���%���I� �m�0��T��x�� ������3���W�� {���P���t������� ������Sw: �^�������= a$Zׯ$� _L�A1��x!1.�ğP��1�Q255.�%�S���2 ��E �//*/<&3F/�� l/~/�/�/<&4�/�50�/�/??<&56?��0\?n?�?�?<&6�?�%@�?��?�?
O1�?P���MY� MY���c��� OQ� �VN<�O �O_�O+_=_O_"_s_�_NPd_�_�_�_�_ �_o!o3o�_Woio{oVNLoM��o�l�o�Ao
.@U}�iRConnec�t: irc\t//alertsE ����Pu�����1�C�UуP_R8�d��H�~��� ����Ə؏���� �2�D�V�S$���8�(p����o͟ߟ���QA8��d�A�@�B4��j�h9�Q+�n�@DM_�A+�~�SMB 	X��8%ğVO��߯���_CLNT 2
X� 4C�ɯ0��l �c�B�T���x���Ͽ ������)�;��_��q�Pϕ��MTP_CTRL ��%���ϙdc���ߋ�@�?�*�c߳l��N����@{�Vߵ�Ƥ�������ѓC���USTOM d{���}�@ }��DTCPIPu��{��h�E�TELҮ{��A���H!�Ta�t�çr�oblolr�  ����!KCL����F��!C�RT��������?!CONS&�����n+���