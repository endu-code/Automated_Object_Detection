��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��#� �8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�? �RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DIS�� S�MB�	"�BC�J@"CI2AI<P6EXPS�!�gPARQ#�SCL�/
 <(C�0��SPTM�E� PW�R��X�V��Ro� l5��!�"%,�7�ICC�%� �kfR�0leP� _D�LV��YNo"3 <oNbX_�P~#?Z_INDE
C�`gOFF� ~UR�i�D��c�  � t �!�`MO�N�%sD�&rHOU�#EWA,vSq;vSq�JvLOCA� Y{$N�0H_HE�K��@I"/ 3 $ARPz&�1�F�W_\ �I!F�`;FA�Dk01#��HO_� INFOv�sEL	% P dK  !k0WO`� $ACCEF� LVZk�2H#�ICE�L���$<�s# ���k���%
��
`�K`SQi��  �55|�I�0ALh�z�X'0 ��
���F����P���܅�$.� 2ċ�� w������� č���!r�Z���4����Ċ!147.8�7.224.204h�S���96�����܁܁3�_{p_ � ċ� bfh.ch̟�1�C� U�g�y���������ӯ�^�� _FLTR � ��π ��
������n�nxč�2n��rSH�PD �1ĉ  P�!
robsta�tion֯՚!k�.�Q�ſ���� ����޿?��c�&� ��JϫϽπ��Ϥ�� ��)���M��"߃�F� ��j��ߎ��߲���%� ��I��m�0��T�� x��������3��� W��{���P���t��� ����������S w:�^���� ��= a$Z�ׯ$ _L�A1>��x!1.�ğ�P�1�Q25c5.%�S���2��E �//*/<&3F/�� l/~/�/�/<&4�/�50�/�/??<&56?��0 \?n?�?�?<&6�?� %@�?�?�?
O1�?P���MY� MY���c��?� Q� �VN<�O�O_�O+_=_O_"_s_�_NPd_�_�_ �_�_�_o!o3o�_Woio{oVNLoM��o �l�oAo
.@U�}iRConn�ect: irc�\t//alertsE����Pu�����1�C�UrуP_R8�d��H� ~�������Ə؏���@� �2�D�V�S$���8�(p����o͟ߟH��QA8��d�A�B4��j�h9�Q�+��@DM_�A�+��SMB 	X�8%ğVO��߯����_CLNT 2]
X� 4C�ɯ 0��l�c�B�T���x� ��Ͽ������)�;���_�q�Pϕ��MT�P_CTRL ��%���ϙdc��� ߋ��?�*�c߳l��N���@{�Vߵ�zƤ����������C��USTOM �{���}�@ �}�DTCPIP�u�{��h�E�TKEL�{��A��ЏH!Ta�t�çroblolr��  ���!K�CL���F��!CRT����������!CONSH&����n+���