��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ��5/IRTU�AL-9LOO�R G��DD?8�?�������k,  1 <DwH82 ������%'����))%��Z�Z]/�o/�/S/�/�/�-_ ��/�/�/;�$MN�U>AP"�� 8���=��?{���<�i��t-�ｇD	?x
� ?tt>2q�n>|l���F��9������0���+�?�&������S�R��������Ѯ���w<S����ʢ�Č���C�-b{5��3��?��;�[��?��7J��j:>�e:>��@�0������AzD����#�
{5��x�?�o;'���7ue��'�&��0��0�<�i�8�/�ȭO�Ę��^���{5?}�z�B��>d����O0f>>����@�>��?�yBB��h�?�%"�=%&C */fO��_O�O�O�O�O��O�E��?���A�H
T��߉������1��<�H)��ʠ �_�� C���%7�NUM  ��>�� "5TOO=L/?4 
E3�O��_�O�_�_  ¢�����ZDCF���_�_e?�+����YC�;��_o=e�1#�B�1�CG���)o;o�V��?�zC���aoso �o�_�o�o�o�o�/l�����33C�@:RW1PfTIVyWV#