��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETGcs��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S�ETHOST� � �DNSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM� !�* �D $PRIM�AR_IG !$?ALTERN1��<WAIT_TI�A �� FT�� @� LOG_�8	�CMO>$DNLD_FI:��SUBDIRCAP�5� �8 .� 4� H�A�DDRTYP�H NGTH��Y�z +LS�&$ROBOT2�PEER2� MA�SK4MRU~O�MGDEV�����RCM+� ;$Z ��QS�IZ�X�� TA�TUSWMAIL�SERV $P�LAN� <$L�IN<$CLU����<$TO�P7$CC�&FR�&��JEC�!�%EN�B � ALARl!B�TP�3��V8 S��$VA5R9M ON
6���
6APPL
6PAp� 5B 	7POR��#_�!�"ALER�T�&�2URL �}�3ATTAC���0ERR_THRO�3US�9z!�8�00CH- Y�4MA�XNS_�1�NAMOD�AI� �$B� (APoWD  � LA ��0�NDATRYQFDELA_C@y'>AERSI�A�'�ROtICLK�HM8R0�'� XML+ :3_SGFRM�3T� �XOU�3PING_�_COPA1�Fe3��A�'C�25�B_A�U�� k 6R,2CO�U�!H!UMMY1zRW2?�RDM*}T $DIS�]� SMB�	"&�BCJ@"CI2�AIP6EXP9S�!�PARQ$�R{CL�
 <(yC�0�SPTM�E� PWR��X�ViQ{SMo l5Ȥ�!�"%�7�ICC"�%� kfR�0le=P� _DLV��Y)No3 <oNb�X_�P~#Z_INsDE
C�`OFF� ~UR�iD��c� �  t ��!�`MON�%sD\�&rHOU�#EWA�,vSq;vSqJvLOC�A� Y$N�0H�_HE���@I�"/ 3 $AR�Pz&�1F�W_�\ �I!F�`;FAp�Dk01#�HO_� oINFO�sEL	%G P K  !�k0WO` $oACCE� LVtZk�2H#ICE��L���$�s# �S��k���
��
`�rK`SQi��P��5|�I�0AL`h�z�'0 ��
����F����P�܅��$� 2ċ T"�w������� č��!r�Z���4����Ċ!147�.87.224.�20h�S���96�����܁܁3�_{p_�  ċ� ?bfh.ch̟� 1�C�U�g�y����������ӯ^�� _FLT�R  ��π *��������n�ndxč2n��rSH�P�D 1ĉ � P!
robs?tation֯՚!k�.�Q�ſ ��������޿?�� c�&χ�JϫϽπ��� �����)���M��"� ��Fߧ�j��ߎ��߲� ��%���I��m�0�� T��x�������� 3���W��{���P��� t������������� Sw:�^�� ����= ah$Zׯ$ _L�A�1��x!1.��ğP�1�Q�255.%�S	���2��E �//*/<&3F/��  l/~/�/�/<&4�/�@50�/�/??<&56?���0\?n?�?�?<&6 �?�%@�?�?�?
O1��?P��MY� MY��c���� Q� �VN<�O�O_�O+_@=_O_"_s_�_NPd_ �_�_�_�_�_o!o3o �_Woio{oVNLoM ��o�l�oAo
.�@U}iRCo�nnect: i�rc\t//alertsE���� Pu����1�C��UуP_R8�d��H�~�������Ə؏ ���� �2�D�V�S$���8�(p����o ͟ߟ��QA8�	�d�A�B4��j�h�9�Q+��@DM_�A+��SMB 	X�8%ğVO���߯���_CLNTw 2
X� 4C�ɯ0��l�c�B�T� ��x���Ͽ������ )�;��_�q�Pϕ���MTP_CTRL ��%���ϙd c���ߋ��?�*�c�d�l��N���@{��Vߵ�Ƥ��������ѓC��USTOOM {���}�@ }�DTCP+IPu�{��h�E.�TEL�{��A=���H!Ta�t��çroblo�lr�  ���!KCL���F�>�!CRT����������!CO#NS&����n+���