��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d PPINFO{EQ/  ��L A �!�%�!� H� �&�)EQUIP 3� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1dQDDd!OE4LA� �R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Dc@�D5�F6�F7*�F8�F9�G0�G�G@JA�E�GbA�E�G1�G!1�G �F�G2�B!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HO30IO�0� }%�SMACRO�ROREPR�X� D+��0��R{�T UT�OBACKU��0 �)DE7VIC�CTI*0�A� �0�#�`B�S�$INTERVA�LO#ISP_UN9I�O`_DO>f7�uiFR_F�0AI�N�1���1c�C�_WAkda�jOF�F_O0N�DEL��hL� ?aA�a1bc?9a�`C?��P��1E��#sATB��d��MO� �cE' D [M�c���^qREV�BI5Lrw XI� Qr�R  � O�D�P�q$NO^PM�Wp�t�r/"�w� �u�q�r��0D`S p =E RD_E�pCq�$FSSBn&$�CHKBD_SE�^eAG G�"$SLOT_��2=�� V�d�%��3 �a_EDIm  � � �"���PS�`(4%$EP<�1�1$OP�0�2��a�p_OK�UST1P_C� ��dx��U �PLACI4!��Q�4�( raCOsMM� ,0$D冀���0�`��EOWBh@BIGALLOW�G (K�"(2�0VARa��@�2B �p�BL�0OUy� !,Kvay��PS�`�0�M_O]����CCFS_UT~p0 "�1�3�#�ؗ�`X"�}R0  4�F IMCM�`O#S@�`��upi �_�p��BA!���M�/ h�pIMPEE_F�N��N�`��@O��r�D_��~�n�Dy�F� dC�C_�r0  T0� '��'�DI�n0�"��p�P�C$I������F�t7 X� GRP0�z�M=qNFLI�<7��0UIRE��$�g"� SWITCH^5�AX_N�PSs"�CF_LIM�� � �0EED��!��qP�t�`P�J_dVЦMODE�h�.Z`�PӺ�ELBOF� �������p� ���3���� F@B/��0�>�G�� �� WARN	M�`/��qP��n�wNST� COR-�0bFLTRh�T�RAT�PT1�� $ACC1a��N ��>r$ORI�o"6V�RT�P_S��pWCHG�0I��rQT2��1�I��T��I1��� x �i#�Q��HDR�BJ; CQ�2L�3�L�4L�5L�6L�7�L� N�9s!$�O`S <F +�=��O��#92��LLEC�y�"MULTI��b�"N��1�!���0T��� �STY �"�R`�=l�)2`�p���*�`T  |�  �&$��۱m��P�Ḻ�UTO���E��EXT����ÁB���"2� (䈴![0������<�b+��� "D"���ŽQ���<煰kcl�9�# ���1��ÂM�ԽP���" '�3�$ L� E���P<��`=A�$JOBn�T����l�TRIG3�% dK�������<���`\��+�Y���_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`��Z���0� �C�P_�P��@ ( @�F RO.��&�t�I9T�c�NOM�
�����S����P`T)"w@���Z�P�d���RA�0��2b"�����
$T����MD%3�T��`U31��ʩp(5!HGb�T1�*E�7�c�KAb�pWAb�cA4#YNT��>�PDBGD�� *(��PUt@X���W���AX��a��ewTAI^cBUF��"0!+ � l7n�PIW�*5 P�7M�8M�9
0�6}F�7SIMQS@�>KEE�3PAT�n�^�a" 2`#�"!_�L64FIX!,C ���!d��D�2B�us=CCI�:FPCH�P:BAD�aHCE hAOGhA]HW�_�0>�0_h@�f�Ak���F��q\'M`#�"H�GE3�- l�p3G��@FSOES]FgHBSU��IBS9WC��. `{ ��MARG쀜���FACLp�SLEWxQe�ӿl�BMC�/�>\pSM_JBM��� �QYC	g�e��R��0 ā�CHNv-�MP�$G� �Jg�_� #��1_3FP$�!TCuf!À�#�����d�#a��V`&��r�a;�fJR�о�rSEGFR�PIyO� STRT��N��cPV5�B�!41�r��
r>İ�b��BBO�2` +�[���,qE`&�,q�`y�Ԣ}t��yaSCIZ%���t�vT�s�� �z�y,qRSINF}Oбc���k��`��`�`L�ĸ T`7�gCRCf�ԣCC/��9��`a�uah�ub'�MIN��uaDs�#�G�D�YC��C�����e`�q0��� �EV�q�F�_�eF��N@3�s�ah��Xa+p,�5!�#1�!VS�CA?� A��s1�"!3 ��`F/k� �_�U��g��]��C�� �a�s�.bR�4� ����N����5a��R�HANC��$cLG��P�f1$+@�NDP�t�AR5@N�^��a�q���c��ME`�18���}0��RAӆ��AZ 𨵰�%O��FCTK��s`"r�S�PFADIJ�OJ�ʠ�ʠ���<���Ր��GI�p�BMP�d�p�Dba���AES�@	�K�W_���BAS�� �G�5�  M�I�T�GCSX[@@�!62�[	$X���T9��{sC��N�`�a~P_�HEIGHs1;�W�ID�0�aVT ACϰ�1A�Pl�<����EXPg���|���CU�0MMENU���7�TIT,AE�%)�a2��a�δ�8 P� a�EDr�E.`��PDT���REM.��AUTH_KEY  ��$���� �b�O	�.a�}1ERRLH� �9c \� �q-�OR�D�B�_ID�@l �PU�N_O��Y�$SCYS0��4g�-�I��E�EV�#q'�P�XWO�� �: G$SK7!f2%�Td�wTRL��; �'�AC�`��ĠIND&9DJ.D��_��f1���f���PL�AF�RWAj���SD�A���A+r|��UMgMY9d�F�10d��&���J�<��}1PR�� 
3�POS���J�= �M$V$�q�PL~�!>���SܠK�?�����CJ�@����ENE�@T��A���S_��RECOR��B�H 5 O�@=$LA�>$~�r2�`R��`�q�b`�_Du�&�0RO�@�aT[�Q� �b������! }У��PAUS���dETgURN��MR�U�  CRp�EWyM�b�AGNAL:�s2$LA�!�?$PX�@$P��y A �Ax�C0 #ܠDO�`X�k��W�v�q�GO_AWAY��MO�ae����]�CSS_CCwSCB C �'N��CERI��гJ`u�QAP�}�\�@�GAG� R�0��`��{`��{`O�F�q�5��#M�A��X��!�L�L�D� �$ ���sU�D)E%!`��>�OVR10W�,��OR|�'�$ES�C_$`�eDSBIOQ��l ��B�VIB&� �c,��p���f�=pSSW�l��f!VL��PL��>�ARMLO
��`a����d7%SC ��bALspH�MP Ch �Ch �#h �#h 5�UU���C�'�C@�'�#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$�4�C�P3Wұ46�$VOLT37$$`�*�^1��$`�O1*�$o��0RQ�Y��2b4�0DH_THE����0SЯ4�7ALPH�4�`��D�7�@ �0�qb7�rR�5�88� ×����"��Fn�M�ӁVHBPFUAFL�Q"D�s�`�THR��i2dB�����G(��PVP���������
��1�J2�B�E�C�E�CPSu�Y@��Fb3 ���H�(V�H:U�G�@
X0��FkQw�[�Na��'B���C INHBcFILT���$ ��W�2�T1�[ ���$���H YАAF�sDO��Y�Rp�  fg�Q�+�c5h�Q0�iSh�QPL���W<qi�QTMOU�#c �i�Q\��X�gmb��vi��h�bAi�fI�aH!IG��ca	xO��ܰ4��W�"vAN-u!���	#AV�H!P�a8$P�ד#p�R_�:�A�a�T"�N80�X�MCN���f1[1�qVE�p��Z2;&f�I�QO�u�rxZ�wGldDN{G|d���aF>!�9��aM�:�U�FWA�:�M l���X�Lu��$!����!l�ZO����0%O�blF�s�13�DI�W�@��Q���_�|�!CURVA԰&0rCR41ͰZ�C<� r�H�v���<�`��<�(�f�CH�QR3�S����t���Xp�VS_��`�ד�F��ژ����?NST�CY_ E L����1�t�1��U��U24�2B�NI O7�x�����DEVI|� F��$5�R�BTxSPIB�P����BYX����T���HNDG��G H tn���L��Q�C���5��Lo0 H���f��FBP�{tFE{�5�t��T��I�DyO���uPMCS�v�>�f>�t�"HOT�SW�`s�?ELE��J T���e�2���25�� O� ��HA7�E��344�0%Ғ�ܘ�A�K �� MD�L� 2J~PE ��	A��s��tːÈ�s�JÆG!��rD"��0������\�TO��W��	��5�OP�SL{AV�L  \0INPڐ���`%ن�_CFd�M� $��ENU��O�G��b�ϑ]զP�0�`ҕ�]�IDMA0�Sa��\�WR�#���"]�VE�$a�SK�I�STs��sk$��2u���J�������	��Q���_SVh�E�XCLUMqJ2M!ONL��D�Y��|�P�E ղI_V�A�PPLYZP��HI�D-@Y�r�_M�2��VRFY�0��r�<1�cIOC_f��"� 1������O��u��LS���R$DU/MMY3�!���S=� L_TP/Bv��"���AӞ�ّ Ns ���RT_u.�� N�G&r[��O D��P_BA��`�3x�!$F ��_5���H��N����� �� P $<�KwARGI��� �q�2O[�_SGNZ�Q �~P/�/P�IGNs�l�$��^ sQANNUN�@�T<�U/�ߴ�LAzp]	Z�d�~��DEFwPI��@ R @�F�?IT�	$TOTA%��d���!mP�EM�NIY�CS+���E�A[��
DAYS\�AD�x�@��	� �E�FF_AXI?�T�I��0zCOJA ��ADJ_RTRQ��Up��<P�1D �r5̀Ll�T�p? ]P�"p��m8tpd��V 0w��G��������SK��SU� ��CTR�L_CA�� W>�TRANS�6PIDLE_PW����!��A�V��V_��l�V �DI�AGS���X� �/$2�_SE�#TAC���t!�!0z*L@��RR��vPA��4�p ; SW�!�! �  ��ol�U��o3OH��PP� ��sIR�r��BRK'#��"A_Ak���x 2 x�9ϐZs2��%l��W�pt*�x%RQD�W�%MSx�t5AX��'�"��LIFEC�AL���10��N �1{"�5Z�3{"dp5�xZU`}�MOTN°9Y$@FLA�cZgOVC@p�5HE	>��SUPPOQ�ݑ�Aq� Lj (C�1_�X6�IEYRJZRJW�RJ�0TH�!UC��6�X�Z_AR�p��Y2��HCOQ��Sf6AqN��w$N�ICTE��Y `��CACHE�C9�M�P�LAN��UFFIQ@�Ф0<�1	���6
�O�MSW��EZ 8�KEY�IM�p��TM~�S�wQq�wQ#���N�O�CVIE� �[ A�BGL��/�}ӛ?����D?��D\�p�ذST��! �R� �T� �T� �T	��PEMAIf�ҁ|P��_FAUL�I]�Rц�1�U�о�R�DTRE�?^< $Rc�u�S�% IT��BU!FW}�W��N_� 'SUB~d��C|��8Sb�q�bSAV�e�b�u �B��� �gX�^P �d�u+p�$�_~`�e�p%yOTT����s�P��M��OtT�LwAX � ��X~`9#�c�_G�3
P�YN_1�_�D��1 �U2M���T��F��H@ g�`� 0p��Gb-s7C_R�AIK���r�t�RoQ�u7h�q'DSPq��rP��A�IM�c6�\����s2��U�@�A�sM*`I�P���s�!D��6�T!H�@n�)�OT�!6��HSDI3�ABSC���@ Vy���� �_D�CONVI�G���@3�~`	F�!�pd��psq�SCZ"���sMER�k��qFB��k��pEiT���aeRFU:@�DUr`����x�CAD,���@p;cHR�	A!��bp�ՔՔV+PSԕC���	C��pTQғSp�_cH *�LX� :cd�Rqa�| ����W� �U��U��U�	�U�TOQU�7R�8R�9R���0T�^�1k�1x�1���1��1��1��1*��1ƪ2Ԫ2^�k�U2x�2��2��2��U2��2��2ƪ3Ԫ%3^�3k�x�3���To���3��3��3ƪ54Ԣ%�XTk!0�d <� 7h�p�6�p�O��p����NaFDR^Z$eT^`V��Gr����䂴2REMr� Fj��BOVM�z�A�TROVٳDT�`-�MX<�I�N��0,�W!IND�KЗ
w�׀�p$DG~q36��P�5�!9D�6�RIV������BGEAR�IO�%K�¾DN�p��J��82�PB@�CZ_MCCM�@�1��@U���1�f ,②a?� ���PI�!�?I�E��Q�"����`m���g� _0Pfqg RI9e���b�ETUP2_ 3h � �cTD�p�〪�! a���]�bB;AC�ri T�P�b��`�) OG��%p���p��IFI�!`�pm�>��	�PT�"���MR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4�@��Uk��� �T�FS#p�Tl �P���e�qP�p$GEX_���1M�2��2� 3�5��9G ���m ��Ѝ��SW�eOe6DEBcUG���%GR���pU�#BKU_�O�1'� �@PO��I5�5MSf��OOfswSM���E�b�A�0��_E �n �0 ���TERM�oN�ORI+�p�GSM_���b�q��A�r�UP�Rs�� -�1��n�$�' o$SEG�,*> ELTO���$USE�pNFIAU"4�e1���#$p$UFR���0ؐ0O!�0����OT�'��TAƀU�#NST��PAT��P�"P'THJ����E�P r�PV"ART�``%B`8�abU!REL:�aSHFT��V!�!�(_SH+@M$����� ��@N8r����OsVRq��rSHI%0���UN� �aAYLO����qIl����!8�@��@ERV]��1 �?:�¦'�2��%��5�%�RCq��EA�SYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba���
5Po��0�p6OR2�MY� `GR��t2b5n� � ��j��a�Uu Ԭ")�.��TOCO!S�1POP ��`�pC��������Oѥ`REPR3��aO�P�b�"ePR�%WU.X1���e$PWR��I�MIU�2R_	S�$VcIS��#(AUD���Cv" v���$H���P_ADDR��H�G�"�Q�Q��QБR~pDp1�w H� SZ�a��e�0ex�e��SE��r���HS��MNvx ���%R́��OL���p<P��<-��ACROlP_!QND_C��ג�1<�T �ROUPT��BI_�VpQ�A1Q� v��c_��i���i��h�x��i���i��v�AC&k�IOU��D�gfsxu^d�y $|��P_D��VB`bP�RM_�b$�HT�TP_אHaz =(��OBJEr��P���$��LE�#|�s`{ � ��.u�AB_x�T~��S�@�DBGLVKRL�YHIT�COU�BGY LuO a�TEM��`e�>�+P'�,PSS|��P�JQUERY_wFLA�b�HW���\!a|`u@�PU�b�PIO��"�]��ӂ/dԁ=dԁ�� ��IOLN��}��z��CXa$SLZ��$INPUT_&g�$IP#�P��'�&��SLvpa~��!��\�W�C-�B��IO^�pF_ASv��$L ��w �F1G�U�B0m!����0HY��ڑ����U;OPs� `�������[�ʔ[�і"�[PP �SIP�<�іI�2���?P_MEMB��i`7� X��IP�P�b�{�_N�`����`R�����bSP����p$FOCUSB�G�a�PUJ�Ƃ �  � o7JOG܄'�DIS[�J7��cx�J8�7� I�m!�)�7_LAB�!�@�A��APHMIb�Q�]�D� �J7J\���� _K�EYt� �K^ՀLMONa����$XR��ɀ��WATCH_��3��&�EL��}Sy~���&s� �Ю!V�g� �CTR3򲓥��;LG�D� �R���I�
LG_SIZ����J�q IƖ�I�FDT�IH�_�jV�G� �I�F�%SO���q �ƀ����v��ƴ��K�S ����w�k�N����E��\���D'�*�U�s5��@L>�n4�DAUZ�EA�p0Հ�Dp�f�GH�B�qBOO���3 C���PIT����� ��REC��SCRN����D_p�aMARGf�`��:� ��T�L���S�s���W�Ԣ�Iԭ�JGM�O�MNCH�c��F�N��R�Kx�PRG�v�UF��p0��FW�D��HL��STP���V��+���Є�RES��H�@�몖Cr4@��?B��� +�O�U�q���*�a28����Gh�0PO��������M8�Ģ��EX��TKUIv�I��(� 4�@�t�x�J0J� ~�P��J0��N�a�#�ANA��O"�0VA�IA��dCLEAR~�6DCS_HI"��/c�O�O�S�I��S��IGAN_�vpq�uᛀT�dn� DEV-�LLAL �°BUW`��x0T<$U�E�M��Ł����P��A
�R��x0�σ�a��@OS1�2�3���_�`� ��ࠜh�AN%-���-�IKDX�DP�2MRO�X�Գ!�ST��Rq��Y{b! �$E&C+��p.&A&p�P���`� L���ȟ%Pݘ��T\Q�UE�`�U���_ � �@(��`�����# �MB_PN@ �R`r��R�w�TRIqN��P��BASS\�a	6IRQ6�@{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?0�?RIAt�MID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCESH?R`�BMhPa����BD4��B�q`�`�F_A�J�C[��O�H� K��� \ȶ��bTf$� ��LI��q�SREQUIR�E�#MO�\�a�XD�EBU���AL� M䵔 �p���P�c�AA�AN��
Q�qa�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N�i�PST9� � �4��LOC�RI쀀�EX�fANGx��AQODAQ䵍��@$��9�ZMF�����f��"��%8u#ЖVSUP�%��FX�@IGGo�� �rq�"��1��#B��$���p%#by���rx���vbPDAT�AK�pE;���� �aIIN*� �t�`MD�qI��) �v� �t�A�wH�`���tDIAE��sAN�SW��th���uD��)ED�`ԣ(@$`�� PCU_�V06�ʠ�d�PLOr�$`��R���B���B�pp������ARR2�E��  ��V�A�/A d$CALII�@��G~�2���!V��<$R�S�W0^D"��ABC~�hD_J2SE�Q\�@�q_J3M�
G�G1SP�,��@PG�Bn�3m�u�3p�@���JkC���2'AO)IyMk@{BCSKP^:�ܔ9�wܔJy�{BQ�ܜ�����`_A1Z.B��?�EL��YAOCMP�c|A)���RT�j���1�ﰈ��@1�������Z��SMG��pԕf� ER!��,0[INҠACk�p����A�n _���@����D�/R��3DIU��CDH�@
�:#a�q$V�Fc6�$x�$���`�@���b��̂�E��H �$BEL�P����!ACCEL����kA°IRCS_R�p�@�T!��$PS�@B2Lʀ���W3�ط9�< ٶPATH��.�Dγ.�3���p�A_ ��_�e�-B�`C����_MG�$DDx��ٰ��$FW�@��p����γ����DE���PPABN�R?OTSPEEup��O0��DEF>Q���ʀ$USE_���JPQPC��JYh����-A 6qYN�@�A�L�̐�L�MO�U�NG��|�OL�y�INCU��a���ĻB��ӑ�AENCS���q�B�����D�IN�I�����pzC��VE�����23�_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��PR9C����MOS� gT�MOpp�@-GPERoCH  M�OVӤ �����!3�yD!@e�]�6�<�� ʓA����LIʓdWɗ��:p83�.�I�TRKӥ�AY����?Q^���m��b��`p�CQ�� MOM�B?R�0u��D����y�0Â��DU�ҐZ�S_BCKLSH_C����o�n� ��TӀ���
c��CLALJ��A��/PKCHKO0�SNu�RTY� �q���M�1�q_
#c�_U�MCP�	C���SC�L���LMTj�_AL�0X����E� � �� ���m�0h���6��PC����!H� �P�ŞCN@�"sXT����CN_��1N^C�kCSF����V6����ϡj���nnCAT�SHs �����ָ1���֙����������PA���_	P���_P0� e���0O1u�$xJG� P�{#�OG���TORQU(�p�a�~���`�Ry������"_W�� ^�����4t�
5z�
5UI;I ;Iz�F�``�!��_8�1��VC��0�D�B�21�>	P�?�B�5JRK�<�2�6~i�DBL_SM�Q:&BMD`_DLt�&BGRV4
Dt�
Dz���1H_���31�8JCcOSEKr�EHLN�0 hK�5oDt�jI��jI<1�J�LZ1�5Zc@y��1cMYqA�HQBTHWM�YTHET09�N�K23z�/Rn�r@C�B4VCBn�CqPASfaYR<4gQt�gQ4V�SBt��R?UGTS���Cq��a��P#��<�Z�C$DUu ���R䂥э2�Vӑ��Q��r�f$NE�+pI�s@�|� �$R�#QA�'UPeYg7EBHBALP!HEE.b�.bS�E�c �E�c�E.b�F�c�j�F�R�VrhVghd��lV��jV�kV�kV�kV*�kV�kV�iHrh�f��r�m!�x�kH�kH��kH�kH�kH�iOJclOrhO��nO�jUO�kO�kO�kO�kO�kO�FF.bTQ����E��egSPBAL�ANCE��RLE6�PH_'USP衅F���F��FPFUL�C�3��3��E��1=�l�UTO_p �%�T1T2t���2N W�����ǡ��5�`(�擳�T�OU���>� INSEG��R��REV��R���DI�FH��1���F�1�;�OB��;C���2� �b�4LCHgWAR��i�ABW!~��$MECH]Q��@k�q��AXk�P���IgU�i�� 
p���!����ROB���CR��ͥ� ��C��_s"T �� x $WEgIGHh�9�$ccd�� Ih�.�IF �N��LAGK�8SK���K�BIL?�OD���U��STŰ�P��; �����������
�Ы�L��  �2�`�"�DEBU�.�L&�n��PMMY9��NA#δ9�g$D&���$���� Q   ��DO_�A��� �<	���~��L�B$X�P�N��+�_7�L��t�OH  ��� %��T���ѼTx�����TICK/�C�T1��%������!N��c�Ã�R L��S���S�����PRO�MPh�E� $IR� X�~ ���!�MAI�0��j���_9����t�l��R�0COD��FU`�+�ID_" =������G_SUFF�<0 3�O����DO��ِ��R��� �ن�S����!{�����u�	�H)�_FI���9��ORDX� ����36��X�����GR9�S��ZDTD���v��ߧ4 *�L_�NA4���K��DEF_I[�K���g�� _���i��Ɠ�š���IS`i �萚���"��e����4�0Bi�Dg����D� �O��LOCKE A!uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ� {����}��v�Ա� ��g������^��� K�Փ����!w�N��P'���^���,`�W�\�[R�� �sTEFĨ �OULOMB_u��0�VISPI�TY�A�!OY�A�_FRId��(�SI���R�����R�3���W�W���0��0_,�EAS%��!�& "����4p�G;� h� ��7ƵCOEFF_Om���m��/�G!%�S.�߲CaA5����u�GR`� � � $hR� �X]�TME��$R�s�Z�/,)�ER��T;�:䗰�  �]�LL��S�_3SV�($~��q��@���� "�SETU��MEA���Z�x0�u������� � � �� ȰID�"���!*��&"P���*�F�'��A��)3��#����"�5;`*��RE�C���!�t�SKy_��� P	�?1_USER��,���4���D�0��VEL@,2�0���2�5S�I��|��MTN�CFG>}1�  ���=Oy�NORE��3�l�2�0SI���� ��\�UX-�ܑP�DE�A $K�EY_����$gJOG<EנSVIA`�WC�� 1DSWy�x��
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��|�����z�� �@_ERR���! ��S L�-���@���s0BB$BUF�-@X1{ ��MORn�� H	�CU�A 3�z�1Q�
��3���O$��FV��27ࡐbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ųp0=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	����y�z=q�#�}1� @�@;���O&E�RI#A��
N��@X�s�f�tQ��PL}1�,RTv�m�ATU}SRBTRC_T(qR��B �����$ �pƱ��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���U1P(4����PX��؆��q��3�w� �P�G�5� $SUB������t�JMPWAITO�,�s��LOyCFt�!D=�CVF	ь�y����R`�0��CC_C�TR�Q�	�IGN�R_PLt�DBTeBm�P��z�BW)�d���0U@���IG�az��Iy�TNLN��"Z�R]aK� N��`B�0�PE�s���r��f�wSPD}1� L	��A�`gఠ�S��UN��{���]�R!�`BD�LY�2���y �_PH_PK�E��2?RETRIEt��2��b�p0���FI��B� ����8� �2��0DBGL�V�LOGSIZ,$C�KTؑUy#u��D7�_�_T1@�E�M�@C\1aA����R���D�FCHECKLK� ��P�0����@�&�(bLEc�" PEA9�T���P�C߰iPN�����ARh� 0���Ӯ�PO�B?ORMATTnaF��f1h���2�S��U�Xy`	��LB��4��  rEITC�H��8PL)�AL?_ � $��XPRB�q� C,2D�!���+2�J3D���{ T�pPDCKyp���oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYLOYA��m�_1t�2t���J3AR��؀�x�֏�laTIA4��u5��6,2MOMCP@�����������0Bϐ�AD��������PUBk`R��;���;����tQ��z4�` I$PI\Ds�oӓ1�yՕ�w�2�w�Z��I
��I��I���p����n���y�e`�9S|)bT�SPEED� G��(�Е��/���Е �`/�e�>��M��ЕSAMP�6V��/���ЕMO�@ 2@�A��QP���C��n� ����������LRf`kb`�ІE9h�EIN0 9��7S.В9
yxPy�GAMM%�S���D$GETH)bP�cD]��2
��IB�q�I�G$H�I(0;A��LRE�XPA8)LW VM8z)��tg���C5�CHKKp4]�0�I_��h` eT��n�q��eT�,���� �$^�� 1�iPI� RCH_D�313\��30LE�1�1\�o(�Y�7 �t�MSWFuL �M��SCRc��7�@�&��%n�f�SV���PB``�'��!�B�sS_SAV�&0ct5B3NO]�C \�C2^�0�mߗ�u� �a��u���u:e;��1���8��D�P����� ����)��b9���e�GE�3��V�d�M�l�� � �YQL��QNQSR lbfqXG�P�RR#dC Qp� �S:AW70�BA�B[�CgR:AMxP�KCL�H���W�r�(�1n�g�M�!o�� q�F�P@}t$WP �u�P r��P5�R<� RC�R��%�6�`��P� ��qsr X��OD��qZ�Ug�ڐ>D� -��OM#w�J? \?n?�?�?��9�b"��8�PL]�_��� |��X0��bf�Ӏqf��q`�ڏgzf��E�ڐ� d�Fb�"�����FdPB��P�M�QU�� �{ 8L�QCOU!n5�QTHI�HOQBnpHYSY�ES��FqUE�`�"�O���  �P�@\�SUN���Cf�O���� P��Vu��!<����OGRAƁcBe2�O�tVuITe ��q:pINFO������{�qcB��OI��r� (�@SLE�QS��q��p�vgqS����� 4L�E�NABDRZ�PTIONt�����Q���)��GCF��G�$�J�q^r�� R����U�g�@bOS_sED����� �F�R�PK��E'sNU߇وAUT$1܅COPY�����n�00MN����PRUT8R �Nvx�OU��$G[r|f��bRGADJ����*�X_:@բ$P�����P��W��P��`} ��)�}�EX�kYCDR|�NS.�9�F@r�LGO�#��NYQ_FREQ�R�W� �#�h�TsL�Ae#����ӄ �CcRE� s�IF�ᶕsNA��%a�_}Ge#STATUI`<e#MAIL������q t�������EwLEM�� �/0><�FEASI?�B ��n�ڢ�vA�]� � I�p��Y!q]�Lt#A�ABM���E�pr<�VΡY�BASR҈Z��S�UZ��0�$q���RMS_TR;�qb ���SY��	�ǡ��$���>C��Q`	� 2� _�TM������̲��@ �A��)ǅ�i$D�OU�s]$Nj���P�R+@3���rGRIyD�qM�BARS �#TY@�Aa O�p�)�� Hp_}�!�����d�O�P/�� � 9�p�`POR�s��\}���SRV��)����DI&0T����P� #�	�#�4!�5!��6!�7!�8� ��PF�2��Ep$VALUt��%���ֱf�F.��� !;�.1�q�����(F_�AN�#�ғ�Rɀ|(���TOTAL��,S��PW�Il��REGEN�1�c�X��ks(��a���`T1R��R��_S� ��1ଃV�����⹂Z�E��p�q��Vr���7V_H��DA�S�����S_Y,1�R4�S�� AR�P2� >^�IG_SE	s��d��å_Zp��C_��~��ENHANC�a�� T ;�8������INT�.���@FPsİ_OVRsP�`p�`��Lv�҂o��7�}��Z�@�SSLG�AA�~�2 5�	��D��S�BĤKDE�U�LvE���TE�P���� !Y��
�J��$2�IL_MC�x r#_��`TQ�`��q���'j�BV�C�P_� �0�M�	V1�
VU1�2�2�3�3�4�4�
�!����� � m�A�2IN~VIBP���1��2�2�3�3
�4�4�A@-±йS2���p� MgC_Fp+0�0�L	11d���M50Id�%"E� S`�R/��@KEEP_H/NADD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0��#i��#REM�"@�$��½%�!�(U}��e�$HPWD  �`#SBMSK*|)G�qU2:�P~	�COLLAB� ��!K5�B�� ��g��pITI1{9p#>D7� ,�@FLAP���$SYN �<M��`C6���UP_�DLYAA�ErDE�LA�0ᐢY�`A�D�Q� �QSK;IP=E� ���Xp�OfPNTv�A�0P_Xp�rG�p�RU@,G ��:I+�:IB1:IG�9J T�9Ja�9Jn�9J{�9J�9<��RA=s� X���4�%1�QB>� NFLIC�s�@�J�U�H�LwNO_aH�0�"?��RITg�]�@_PA�pG�QO� ��^�U���W��LV�d�NGRLT�0_q��O�  " 8��OS��T_JvA V�	�APPR_WE�IGH�sJ4CH�?pvTOR��vT��LCOO��]�+�tVJ�Є��ғA�Q�U�S�XO1B'�'�{�J2P���7�X�T�<a43 DP=`Ԡ\"<a�q\!��RDC��L� ��рR��R�`� �R�V��jr�b�RGEp��*��cN�FLG�a8�Z���SPC�s��UM_<`^2TH�2NH��P.a 1�� m`EF11��� lQ �!#� <�p3AT� g�S� &�Vr�p�tMq�Lr<���HOMEwr�
t2'r�-?Qc(u��w3'r��������w4'r�'�9�K�]�o����w5'r뤏��ȏڏ���
�6'r�!�3�E�W�(i�{��7'r힟���ԟ����8'r��-�?�Q�c�u��S$0�q�p�� sF�`�`)a�"`P����a�`/���-�IO[�M�I֠��qPOW=E�� ��0�Zatep�� y�5��$DSB OGNAL���0Cp�m�S2323�� Ɍ~`��� / ICEQP��PEp��5PsIT����OPBx0ޣ�FLOW�@TR`vP��!U���CU�M��UXT�A��w�ERFAC�� U���ȳCH��� tQ  _��>�Q3$����OM���A�`T�P#UPD�7 A�ct�T��UE�X@�ȟ�U EFA8: X"�1RSPT��ѧ��T ��PPA��0o񩩕`EXP�IAOS���)ԭ�_�0��%��C�WR�A���ѩD�ag֕`ԦFR�IENDsaC2UFx7P����TOOL���MYH C2LENGTH_VTE���I��Ӆ$SE�����UFINV_t���RGI�N{QITI5B��Xvl��-�G2-�G17� w�SG�X��_��UQQD=#���AS��d�~C�`��q�� ��$$C/�S�`������S0)`����V�ERSI� ��])`�5��I���������AAVM_�Y�2 �� 0  �#5��C�O�@�r� r�	 �����S0���������� ������
?QYf�BS���1��� <- ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O��O�O�OiCC�@XgLMT��C�7  ��DIN�O�A\�Dq�EXE�HPV_��ATQz
���LARMRECOV �RgLMDG *��5�OLM_IF' *��`d�O�_ �_�_�_j�_'o9oKo<]onm, 
��o db��o�o�o�o^���$� z, A  � 2D{�PPIN�FO u[ @�Vw������� �`�������*� �&�`�J���n�����DQ����
��.� @�R�d�v����������a
PPLICATf��?�P��`�Handl�ingTool �
� 
V8.3�0P/40Cpɔ_LI
883���ɕ$ME
F�0G�4�-

�398�ɘ�%�z��
7DC3x�ɜ
�Noneɘ�Vr���ɞ@�6d� Vq_A�CTIVU��C\죴�MODPye��I��HGAPONp���OUP�;1*�� i�m�����Қ_����1�*�  �@���� ����Q���Կ濸@�
����� g���5�Hʵ�l�K�HTTHKY_��/�M�SϹ��� ������%�7ߑ�[� m�ߝߣߵ������� ���!�3��W�i�{� ������������� �/���S�e�w����� ����������+ �Oas���� ���'�K ]o������ ��/#/}/G/Y/k/ �/�/�/�/�/�/�/�/ ??y?C?U?g?�?�? �?�?�?�?�?�?	OO uO?OQOcO�O�O�O�O �O�O�O�O__q_;_ M___}_�_�_�_�_�_�_kŭ�TOp��
��DO_CLEAN�9��pcNM  !{衮o�o�o�o�o���DSPDRY�Rwo��HI��m@ �or����������&�8�J���MAXݐWdak�H�h��XWd�d���PL�UGGW�Xgd��P�RC)pB�`�k�aS�Oǂ2DtSEGF0�K� �+� �o�or����������%�LAPOb�x��  �2�D�V�h�z�����య¯ԯ�+�TOT�AL����+�USE+NUO�\� e�A��k­�RGDISPWMMC.���C6�&z�@@Dr\�OMpo��:�X�_STRI�NG 1	(�
��M!�S��
��_ITEM1Ƕ  n����� �+�=�O�a�sυϗ� �ϻ���������'��9�I/O S�IGNAL���Tryout M�odeȵInp�y�Simulat{eḏOut��OVERRLp� = 100˲In cycl��̱Prog A�bor��̱u�S�tatusʳ	H�eartbeat�ƷMH Fauyl	��Aler� L�:�L�^�p����8������ Scû Saտ��-�?�Q�c�u� ���������������);M_q��WOR.�û���� ��+=Oa s�������8//'.PO���� M �6/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?H"DEVP.�0d/�?O *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�J_\_n_PALT 	��Q�o_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o�_GRIm�û9q�_ as������ ���'�9�K�]�o� ������'�R	�݁ Q����)�;�M�_� q���������˟ݟ����%�7�I�ˏPREG�^����[����� ͯ߯���'�9�K� ]�o���������ɿۿ��O��$ARG_�� D ?	����0�� � 	$O�	+[D�]D��O�e��#�SBN_CON?FIG 
0˃����}�CII_SAVE  O������#�TCEL�LSETUP �0�%  OME�_IOO�O�%M�OV_H������R�EP��J��UTOoBACK�����FRA:\�o� Q�o���'�`��o��ҟ��= �� f�o������*�!�3�`�Ԉ��f�������� ��o�{��&�8�J�\� n�������������� ����"4FXj| �������끁  ��SYS�UIF.SV V� T.TP D �MP 6.VD GIF 7N`r�o�NLQ���f�WINI�Po����c�MESSAG�����8��ODEC_D����z��O�0��c�PAUSM!!��0� (783�U/g+(Od/�/ x/�/�/�/�/�/�/? ??P?>?t?1�0$: ?TSK  @-��<T�f�UPDT���d�0
&XWZD�_ENB����6S�TA�0��5"�XI�S��UNT 2�0Ž� � 	 ���z���eng��-뷛�S��o�U@��H�����tL�Oo�}Cw�gJ�^����.�O��O�O�O/_2FMET�߀2CMPTAA���@�$A�-�@���@����@���]5���5�(d5���P5�r�5F*5�338]�SCRDCFG }1�6��	��Ź�_�_oo (o:oLo��o�Q���_ �o�o�o�o�o�o]o �o>Pbt���o9�i�GR<@M/��sUP_NA��/�	i��v_ED��1�Y� 
 ��%-BCKE�DT-�'�GE�TDATAU�o�9A��?�j�H�o�f��\��A��  ���2�&�!�E���:IB���~�ŏ׏m����3��&۔�� D��ߟJ�����9�ǟ�4���ϯ�(���@�]�o�����5N� �����(�w��)�;�ѿ_��6ϊ�gϮ� (�CϮ���ϝ�+��7��V�3�z�(��z� ����i����8��&���~�]���F�ߟ�5����9~������]����Y�k�����CR�!ߖ���W� q���#�5���Y��p$�?NO_DEL��r�GE_UNUSE���tIGALLO�W 1��(�**TEM*�S	$SERV�_GR�V� : REG�$�\� �NUM�
��P�MUB ULA�YNP\PM�PAL�CYC10#6 $\ULSU�8:!�Lr�BOX�ORI�CUR_���PMCNV6�10L�T4DLI�0��	����BN/`/r/�/��/�/�/�/���pLA�L_OUT ��;���qWD_AB�OR=f�q;0IT_R_RTN�7�o	�;0NONS�0�6� 
HCCFS_U?TIL #<�5�CC_@6A 2#; h ?�?�?O�#O6]CE_OPT;IOc8qF@�RIA_Ic f5�Y@�2�0F�Q�=2q&}�A_LI�M�2.� ���P�]B��KXʊP
�P�2O�Q�R�B�r�qF�PQ 5T1)TR�H�_:J�F_PARAMGoP 1�<g^�&S�_�_�_�_�VC��  C�d�`��o!o`�`�`�
`�Cd��Tii:ah:e>eBa�GgC�`~� D� D	�`m�w?��2HE �ONFI� E?�aG�_P�1#; ���o1C�Ugy�aKPAU�S�1�yC ,�������� �	�C�-�g�Q�w���@������я���rO�A��O�H�LLECT_�B�IPV6��EN. QF�3�ND�E>� �G�7�1234567890��sB�TR�����%
 H�/%) �������W���0� B���f�x���㯮��� ү+�����s�>�P� b����������ο� �K��(�:ϓ�^�|�:�B!F� �I|�IO #��<U%�e6�'�9�K���T-R�P2$��(9X�t�Y޼`%�̓ڥH���_MOR�3&��=��@XB� �a��A�$��H�6� l�~���~S��'�=�r�_A?�a�a`��@K(��R�dP��)F�ha�-�_�'�9�%
�k��G� ��%yZ�%��`�@]c.�PDB��+����cpmidbag��	�`:������p��N  #��@��.���]ܭ@s<�V^��@sg�$�fl�q>��ud1:���:J��DEF *�ۈ��)�c�b?uf.txt�����_L64FIX ,������l/ [Y/�/}/�/�/�/�/ 
?�/.?@??d?v?U? �?�?�?�?�?�?,/>#__E -���<�2ODOVOhOzO�O6&I�M��.o�YU>�c��d�
�IMC��2/����dU�C�Ӌ20�M�QT:Uw�C�z  B�i�A����A���Au��gB3�*C?G�B<�=w�i��B.��B����B��5B�$�D�%B���e�zVC�q�C�v��D���D-l�E\D��n�j��B9"��22�o�D|����� ����C�C�����
�xObi�DY4cdv`D��`/�`�v`s]E�D D��` E4�F*�� Ec��FC���u[F���E���fE��fF���3FY�F��P3�Z��@�33� ;��>L��T�Aw�n,a@��@e�5Y���a���`At��w�=�`<#�*�
��?�ozJRSMOFST (��,bIT1��D @3���
д�'�a��;��bw?��ߚ<�M�NTEKST�1O�CR@��4��>VC5`A��w�Ia+a�aORI`C6TPB�U�C�`4�s��r��:d�*��qI?�5��qT�_�PROG ���
�%$/ˏ�t��N�USER  �U�������KEY_T�BL  �����#a��	
�� �!"#$%&'()*+,-./���:;<=>?@A�BC�GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~�������������������������������������������������������������������������������͓���������������������������������耇�������������������������LCK�
�����STAT/��s_�AUTO_DO ��	�c�INDTO_ENBP���Rpq�n�`�T2����ST�Or`���XC�� �26�) 8
S�ONY XC-5�6�"b����@���F( А�HR50w���>��P�7b�t�Aff����ֿ� Ŀ�� ��C�U�0�yϋ�fϯ� �Ϝ��������-ߜ��TRL��LETE�ͦ ��T_SCREEN �ڟkcs���U��MMENU 1=7�� <ܹ� ��w��������� K�"�4��X�j��� ����������5��� k�B�T�z��������� ������.g> P�t����� �Q(:�^ p����/�� ;//$/J/�/Z/l/�/ �/�/�/�/�/�/7??  ?m?D?V?�?z?�?�? �?�?�?!O�?
OWO.O @OfO�OvO�O�O(y��?REG 8�y�����`�M�ߎ�_M�ANUAL�k�DwBCO��RIGY��9�DBG_ERRML��9�ۉq�ر_�_�_ ^QNU�MLI�pϡ�pd�
�
^QPXWOR/K 1:���_5o�GoYoko}oӍDBT;B_N� ;������ADB__AWAYfS�q/GCP 
�=�p�f�_AL�pR��bbRY��[�
�WX_�P 1<{y�n�,�%oc��P��h_M��I�SO��k@L��sON�TIMX��
�ɼ�vy
��2sMO�TNEND�1tR�ECORD 1B΋� ���sG�O�]�K��{�b���� ����V�Ǐ�]���� 6�H�Z��������� #�؟������2��� V�şz��������ԯ C���g��.�@�R��� v�寚�	���п��� c�χ�#ϫ�`�rτ� ��Ϻ�)ϳ�M��� &�8ߧ�\�G�Uߒ�� ������I������4��� �p7�n���ߤ� ���������"��� F�1���|�������� [�����i���BT�f���bTOLEoRENC�dB�'r��`L��^PCSS�_CCSCB 3IC>y�`IP�t} �~�<�_`r �K�����/�{��5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O��O�O�O_�~�LL� D��&qET�c��a C[C��PZP^r_ A�J� p� �sp��Q<GPt[	 A�p�Q�_�[? �_�[oU��p�P�pSB�V�c�(a�PWoio({h+�o�X�o�o�Y��[	r�hL�W��N:p����}6ګ�c��a�D@VB��|��G���+?��K� �otGhXGr�So�����eB   =���Ͷa>�tYB�D� �pC�p�q�aA"�H�S�Q-��q���u�d�v�����AfP `; 0���D^P�֨p@�a
�QX THQ����a aW>� �a9P��b�e:��L�^�h�Hc�́PQ �RFQ�PU�z�֟�o \^��-�?��c�u�X���zCz�ů�b2�Щ�RD�����l)*����S ̡0��]�0�.��@���EQ�p��F�X�ѿ�Uҁп�VSȺNSTCY 1E�
�]�ڿ��K�]� oρϓϥϷ������� ���#�5�G�Y�k�}���ߒ��DEVIC�E 1F5�  MZ�۶a��	� ��?�6�c���	{䰟����_HNDGD �G5�VP���R�LS 2H�ݠ��/�A��S�e�w����� ZPA?RAM I�Fg�He�RBT 2-K��8р<��WPVpC�C��,`¢PQ�Z�z��%{�C��2�jMTLU,`"nPB, s� �M� }�gT�g��
#B��!�bcy� [2Dchz�����/��/gT#�I%D��C�` �b!�R��A��A�,��Bd��A5��P��_C4kP�!�2�C��$Ɓ�]�f�fA�À��B�� �| ���/�/�T (��54a5�} %/7/d?/M?_?q? �?�?�?�?�?O�?O O%O7OIO�OmOO�O �O�O�O�O�O�OJ_!_ 3_�_�_3�_�_�_�_ �_o�_(ooLo^oЁ =?k_IoS_�o�o�o�o �o�o�o#5G �k}����� ��H��1�~�U�g� y�ƏAo�Տ���2� D�/�h�S���go���� ԟ����ϟ���R� )�;���_�q������� ���ݯ�<��%�7� I�[�m��������� }�&��J�5�n�Yϒ� �Ϗ��ϣ�ѿ���� ��F��/�Aߎ�e�w� �ߛ߭���������B� �+�x�O�a���� ��������,���%�b� M���q����������� ����L#5� Yk}��� � �61CUg �������� 	//h/���/w/�/�/ �/�/�/
?�/.?@? I/[/1/_?q?�?�?�? �?�?�?�?OO%OrO IO[O�OO�O�O�O�O �O&_�O_\_3_E_W_ �_?�_�_�_�_�_"o oFo1ojoE?s_�_�o m_�o�o�o�o�o0 f=Oa��� �������b� 9�K���o���Ώ��[o ��(��L�7�I����m������$DCS�S_SLAVE �L���ё���_4D�  љ��CFoG Mѕ��������FR�A:\ĐL-�%0�4d.CSV�� � }�� ���A Vi�CHq�z����p��|�����  ������Ρޯ̩ˡҐ-矩*����_CR�C_OUT N�������_FS�I ?њ ����k�}����� ��ſ׿ �����H� C�U�gϐϋϝϯ��� ������ ��-�?�h� c�u߇߽߰߫����� ����@�;�M�_�� ������������� �%�7�`�[�m���� ������������8 3EW�{��� ���/X Sew����� ��/0/+/=/O/x/ s/�/�/�/�/�/�/? ??'?P?K?]?o?�? �?�?�?�?�?�?�?(O #O5OGOpOkO}O�O�O �O�O�O _�O__H_ C_U_g_�_�_�_�_�_ �_�_�_ oo-o?oho couo�o�o�o�o�o�o �o@;M_� �������� �%�7�`�[�m���� ����Ǐ������8� 3�E�W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿� ��'�P�K�]�oϘ� �ϥϷ���������(� #�5�G�p�k�}ߏ߸� ������ �����H� C�U�g������� ������ ��-�?�h� c�u������������� ��@;M_� ������� %7`[m� ������/8/ 3/E/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO�sO�O�O�O�O�C�$�DCS_C_FS�O ?�����A P �O�O_?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo ~o�o�o�o�o�o�o�o 72DVz� ������
�� .�W�R�d�v������� ������/�*�<� N�w�r���������̟ ޟ���&�O�J�\� n���������߯گ� ��'�"�4�F�o�j�|� ������Ŀֿ�������G�B�T��OC_RPI�N_jϳ��� �ς��O����1�Z�U��NSL��@&�h߱� ��������"��/�A� j�e�w������� ������B�=�O�a� ���������������� '9b]o� ������� :5GY�}�� ����///1/ Z/U/g/y/�/�/�/�/ �/�/�/	?2?-???Q? z?u?��ߤ߆?�?�? �?OO@O;OMO_O�O �O�O�O�O�O�O�O_ _%_7_`_[_m__�_ �_�_�_�_�_�_o8o 3oEoWo�o{o�o�o�o �o�o�o/X Sew����� ���0�+�=�O�x� s���������͏ߏ� ��'�P�K�]�o������ �PRE_CH�K P۪�A ~��,8�2x��� 	 8�9�K���+�q���a� ������ݯ�ͯ�%� �I�[�9����o��� ǿ��׿���)�3�E� �i�{�YϟϱϏ��� ��������-�S�1� c߉�g�y߿��߯��� �!�+�=���a�s�Q� ����������� ���K�]�;�����q� ������������#5 �Ak{�� ����CU 3y�i���� ��/-/G/c/u/ S/�/�/�/�/�/�/? ?�/;?M?+?q?�?a? �?�?�?�?�?�?�?%O ?/Q/[OmOO�O�O�O �O�O�O�O_�O3_E_ #_U_{_Y_�_�_�_�_ �_�_�_o/ooSoeo GO�o�o=o�o�o�o�o �o=-s� c������� '��K�]�woi���5� ��ɏ��������5� G�%�k�}�[������� ן�ǟ����C�U� o�A�����{���ӯ�� ��	��-�?��c�u� S�������Ͽ῿�� ���'�M�+�=σϕ� w�����m������%� 7��[�m�K�}ߣ߁� ���߷����!���E� W�5�{��ϱ���e� ������	�/��?�e� C�U������������� ��=O-s� ���]���� '9]oM�� �����/�5/ G/%/k/}/[/�/�/� �/�/�/�/?1??U? g?E?�?�?{?�?�?�? �?	O�?O?OOOOuO SOeO�O�O�/�O�O�O _)__M___=_�_�_ s_�_�_�_�_o�_�_ 7oIo'omoo]o�o�o �O�o�o�o!�o1 W5g�k}�� ����/�A��e� w�U�������я��o ����	�O�a�?��� ��u���͟����� '�9��]�o�M����� ����ۯ��ǯ�#�ů G�Y�7�}���m���ſ �����ٿ�1��A� g�E�wϝ�{ύ����� ��	�߽�?�Q�/�u� ��e߽߫ߛ������� �)���_�q�O�� ������������ 7�I���Y��]����� ����������!3 WiG��}�� ��%�A�1 w�g����� �/+/	/O/a/?/�/ �/u/�/�/�/�/? �/9?K?�/o?�?_?�? �?�?�?�?�?O#OO GOYO7OiO�OmO�O�O �O�O�O_�O1_C_%? g_y__�_�_�_�_�_ �_�_o�_+oQo/oAo �o�owo�o�o�o�o �o);U__q� �������%� �I�[�9����o��� Ǐ�����ۏ!�3�M ?�i��Y�������՟ �ş����A�S�1� w���g�����������ӯ�+�=��$DC�S_SGN Q�K�c��7m� �29-MAR�-19 10:2�5   O�1�4-JANt�08�:38}�����? N.DѤ���𖲸���h�x,r�Wf*σ�^M���  O�VERS�ION [��V3.5.13��EFLOGIC� 1RK��  	����P�?�P�N�!�PRO�G_ENB  ⸴6Ù�o�ULSOE  TŇ�!�_ACCLIM�Ư��Ö��W?RSTJNT��c�;�K�EMOx̘���� ���INIT �S.�G�Z���OPT_SL ?	,���
 	R5�75��Y�74^�6Z_�7_�50��1���2_�@ȭ��<�TO�  Hݷ���V.�DEX��dc�����PATH A[�A\�g�y���HCP_CLN�TID ?��6�� @ȸ����I�AG_GRP 2�XK� ,`���� �9��$�]�H�����1�23456789q0����S�� |��������!�� ��H���;�dC�S���6���� �.�Rv� f��H��// �</N/�"/p/�/t/ �/�/V/h/�/?&?? J?\?�/l?B?�?�?�? �?�?v?O�?4OFO$O jO|OOE��Oy��O �O_�O2_��_T_y_�d_�_,
�B^ 4 �_�_~_`Oo�O&oLo ^oI��Tjo�o.o�o�o �o�o �O'�_K6 H�l����� ��#��G�2�k�V� ��B]���Ǐُ��������(��L�B\Dr�x�@��PC�����4  79?֐�$��>��� :�����ߟʟܟ����CT_CONFI/G Y��Ӛ��egU���STBF_TTS�ǁ
��b����Û�u��O�MAU��|��M_SW_CF6�Z���  �OCVI�EW��[ɭ������-�?�Q�c�u� G�	�����¿Կ��� ���.�@�R�d�v�� �ϬϾ�������ߕ� *�<�N�`�r߄�ߨ� ����������&�8� J�\�n���!���� ���������4�F�X��j�|����RC£\�e��!*�B^�������C2g{�SB�L_FAULT �]��ި�GPM�SKk��*�TDI�AG ^:�ա�I��UD1:� 6789012�345�G�BSP �-?Qcu�� �����//)/�;/M/� �
@�q��/$�TREC	P��

��/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO�0OBOi/{/xO�/UM�P_OPTIONk���ATR¢l��	��EPMEj��OY�_TEMP  ?È�3B�J�Ps�AP�DUNI���m�Q��YN_BR�K _ɩ�EMGDI_STA"U��aQSUNC_S1`ɫ �FO�_�_�^
�^dpOoo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{�E�����y �Q��� �2�D�V� h�z�������ԏ� ��
��.�@�R�d��z �������˟��� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i��������� ÿݟ�����/�A� S�e�wωϛϭϿ��� ������+�=�O�a� {�iߗߩ߻�տ���� ��'�9�K�]�o�� ������������� #�5�G�Y�s߅ߏ��� ��i�������1 CUgy���� ���	-?Q k�}�������� �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?u?�? �?�?��?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_m?w_�_�_�_�?�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9Ke_W� ���_�_���� #�5�G�Y�k�}����� ��ŏ׏�����1� C�]oy�������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;���g�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�_�i�{ߍߟ߹� ����������/�A� S�e�w������� ������+�=�W�E� s������ߧ������� '9K]o� ������� #5O�a�k}�E ������//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-?GY c?u?�?�?��?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_Q?[_m__�_ �?�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/I_ Sew��_��� ����+�=�O�a� s���������͏ߏ� ��'�A3�]�o��� ����ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����9� K�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ���ߑ�C�M�_�q� �ߝ��߹�������� �%�7�I�[�m��� ������������!� ;�E�W�i�{��ߟ��� ��������/A Sew����� ��3�!Oa s�������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? +=G?Y?k?!?��? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	_#?5??_Q_ c_u_�?�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o -_7I[m�_� �������!� 3�E�W�i�{������� ÏՏ����%/�A� S�e�q�������џ �����+�=�O�a� s���������ͯ߯� ���9�K�]�w��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����������'�1� C�U�g߁��ߝ߯��� ������	��-�?�Q� c�u��������� ��m��)�;�M�_�y� �������������� %7I[m� �������! 3EWq�{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/�/+?=?O?i _?�?�?�?�?�?�?�? OO'O9OKO]OoO�O��O�O�O�O�O�O? ��$ENETMO�DE 1aj5�  0�054_F[PR�ROR_PROG %#Z%6�_�Y�dUTABLE  #[t?�_�_�_g�dRSEV_NUM� 2R  ��-Q)`dQ_AUT�O_ENB  �PU+SaT_NO>a �b#[EQ(b W *��`��`��`	��`4`+�`�o�o�oZdHIS%c1+PSk_ALM 1c#[� �4�l0+�o;M_q��r�o_b``  #[�aFR�zPTCP_VER !#Z�!�_�$EXTL�OG_REQ�f9�Qi,�SIZ5�'��STKR�oe�~)�TOL  1{Dz�b�A '�_BWD�p��Hf���D�_DI�� dj5SdDT1KRņSTEPя�P���OP_DOt�QF�ACTORY_T�UN�gd<�DR_?GRP 1e#YNa�d 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ�ԟ ���1��U�@�y�d��v�����ӯ����LW
? J�'��,��tۯ�j�U���y��B�  B୰�>��$  A@��s�@UUUӾ����Ͼ��E�� E�`F@ F�5U/��,��L���M���Jk�Lz�p�JP��Fg{�f�?�  s���9�Y9}��9��8j
��6��6�;���A����O ��� �� I �������[FEATUROE fj5��JQ�Handl�ingTool �� "
P�English �Dictiona�ry�def.�4D St�a�rd�  
! �hAnalo�g I/OI�  �!
IX�gle� ShiftI�d��X�uto So�ftware U�pdate  r�t sѓ�mati�c Backup~�3\st���ground E�dit��fd�
Camer�a`�Fd�e��Cn?rRndIm����3�Common� calib U}I�� Ethe��n��"�Monit{or�LOAD8��tr�Relia�by�O�ENS�Da�ta Acquiys>��m.fdp�?iagnos��]��i�Document VieweJ���870p�ua�l Check �Safety*� �cy� �hanceod Us��Fr�����C �xt. oDIO :�fi��s m8���end��ErrI�L��S�������s  t P%a�r[�� ����J944FCTN Menu��ve�M� J9l�T�P InT�fac�{�  744��G���p Mask �Exc��g�� R�85�T��Pro�xy Sv��  �15 J�igh�-Spe��Ski>
� R738Г�~�mmunic���ons�S R7���urr�T�d�02�2��aю�conn�ect 2� J�5��Incr��s�tru,Қ�2 R�KAREL �Cmd. L��u�a��R860hR�un-Ti��En�vL�oa��KU�e�l +��s��S/�Wѹ�7�Lice�nse���rod�u� ogBook�(System)��AD pM�ACROs,��/�Offs��2�NDFs�MH�� �����MMRC�?��O�RDE� echS�top��t? � 84fMi$�|� 13dx��]е��܏���Modz�witchI�VP��?�:��. sv��2Optm�8�2���fil��I ��2g� 4 !+ulti-T�����;��PCM funY�Po|���4$��b&Regi� r\ �Pri��FK+�7���g Num �SelW  F|�#�� Adju����60.��%|� �fe���&tatuď!$6���%��  �9 J6RDM Robot)��scove2� 5;61��RemU�=n@� 8 (S�F3Servo�����)SNPX� b�I�\dcs<�0}�Libr1��OH� �5� fl�0��58��So� =tr�ssag4%G /91�p ���&0���p/I�� � (ig TMIL�IB(MӋ�Firm����gd7���s�'Acc����0�XAsTX�Heln���*LR"1��Sp�ac�Arquz�iOmulaH��� Q�n��Tou�Pa�D�I��T��c��&���ev. f.sv�USB po���"�iP�a�� � r"1Unexcept��`0i$/���n�H59� VC&�r��[6���P{�<�RcJPRIN�V�;� d T@�TSP� CSUI�� r��[XC��#Web� Pl6�%d -c�1R�@4d������I�R66?0FV�L��!FVGridK1play C�lh@X����5RiR�R.@�~��R-35iA|���Ascii��8�"��� 51f�c�Upl� � (T�����S��@rit�yAvoidM l�`��CE��rkδCol%�@�Gu"F� 5P��j}P�����
 B�L�t� 120C C� o�І!J�D�P��y��� o=qz�b @DCS b ./��c��O��q��D`�; ���qckpgaboE4�DH@��OTШ�main �N��1.�H��an�.��A> aB!FR�LM���!i ���M�I Dev�  (�1� h8j��spiJP��� �@��Ae1�/�r���!hP� M-2� i��߂^0ii�p6�PC���  iA/'�Pa�sswo�qT�RGOS 4����qedav�SN��Cli����G6x Ar�� �47�!���5s�DsER��Tsup>Ryt�I�7 (M�aΪT2DV�
�3D Tri-���&���_8;�
�A�@D�ef?����Ba�: deRe p 4�t0��e�+�V�s�t64MB DR;AM�h86΢�FRO֫0�Arc�� visI�ԙ�n<��7| ), �b��Heal�wJ�\h���Cell`��p� �sh[��� Kq:w�c� - �v�b��p	VCv�tyy�ys�"Ѐ6�u�t��v�m���xs ���TD_0��J�m㖙` 2��a[�>R �tsi�MAILYk�/F2�h��ࠛ 90 H��F02�]�q�P5'���T10C��5����FC��Uz�F9�GigEH��S�t�0/A� if��!2��boF�dr�i=c �OL�F�S����" H5�k�OPT ��4�9f8���croP6��@��l�ApA��Syn.(RSSG) 1L�\1y�rH�L� (2x5�5�d�p�CVx9����estb�$SР��> \pϐ�SSF�e$�tex�D o���A�	� �BP���a�(R00��Qirt��:���2@)�D��1�e�VKb@_l Bui, n��WAPLf��0��1Va�kT�XCGM��D���L����[CRG�&a�YBU��YK�fL��pf��k�\sm�ZTAf�@�О�Bf2�и��V#�s�d��� r���CB��@�
f���WE��!!��
���T�p��DDT�&4 Y�V�`��EH����
�#61Z��
�R=2�
&�E (Np��F�V�P K�B���#��Gf1`?G���H�р?eI�e ����LD�4L��N��7\s@����`���M��deSla<,��2�M�� "L[P��`?@��_�%�����S��M-F�TSO�W�wJ57��VGF��|�VP2֥ 5\ b�`0&�cV:���T;�T� �<�ce,�?VPD��$
eT;F��DI)�<�I�a\so<��a-�6Jc6s6�4L�M�bV9R�h���Tri� � ���5�` �f�@�������P
� ����`>��Img PH�[�l��I/A  DVP�S��U�Ow���!%S�Skastdp�n)ǲt�� SWI�MEST�BFe�00��-Q� �_�PB�_�Rued�_�T��!�_�S ��_bH573o2c2��-oNbCJ5N�Iojb)�Cdo�cxE��o�_�lp��o �TdP�o�c�B�or�2 .rٱ(Jsp�Efr�SEo�f1�}�r3s RGoeELS��sL����s������B	��S\ $�F�ryLz�ftl�o~�g�o ���������?������P  �n�&�"�l  ��T�@<�^��Y��e��u8Z���alib��Γ��ɟ3����f��\v ��e\c��6�Z�f�T�v�R �VW���8S��UJ9�1����i�ů[c91�+o�w8���847�:��A4�j��Q���t6�m���vrc.�����HR���ot8�0ݿ��  ���8ޯ�460�>eS0L�97���U���Ϧ�60.� g�н�@+��'�ܠ�Ϻ�8co&��DM߱U"����d�ߕpi�߲T! �&�na;�� ���u%��ⅰI��lo`R�d��1a59gϘ�ŭ���95�ϔ�R����1��?��o�#� �1A�/���vt{�U�Weǟ���ￇ73�[���7�ρ�C WL��62K�=fR���8��������d����2�ڔ����@��@" "http�����t7 ��� v R7��78�����4�� ��TT�PT�#	��eP#CV4/v߀�j�Q�Fa7��$N�0�/2��rIO�)/;/M/6.sv3�64i�oS�l? torah?*�|`�?��AM/�?
??p.?0�k/��1 JO0��� ,O�tro���0[P��OB4c.K?�g�'�)�24g?�� (1B�Od�\iOA5csb�?U_�?vi�/i��/�/Wn��`�o%�Fo�4l�$of���oXF I)xo�cm3p\7��mp���d�uC��lh����o(AA�_Bt� �o]6P���m�I?�w�@���na$O��4*O0wi�8%P�?"�bsg?�]7��YEM���8woVJ̇/ե11?o��DMLs�BC��7J��\���(�52�XFa AP�ڟ<�v�`/ş�aqs����/OIf��1�9��VRK���ph�քH�5+�=�IN/¤SckiW�/�IF�0�_�%��fs�I�O�l����"<𜿚$�`����\jԿz5bON�vrouς�3(�ΤH (DϮ��?sG ��|��F�Ou������ �D)O��*�3P$� FӅ�k��ϻ���럴�� �PL��ʿ��pb3ox�ߦebo����Sh �>�R.�0wT{����fx6��P���D��3��#_I\Im;YEe�OԆM�8hxW�=Ete,���dGct\���O$kR�������Xm*���r�o3��D�l�j9���V'�  FAC���|@�ք f?6KARE0�_�~� (Kh��.cf���WpoO�_K�up��a���H/j#�- Eqd/�84���$qu�o��/ o2o?Vo<�7C�)�s��NJԆ�|?�3l\�sy�?�40�?Τwaio�u]?�w58�?�,F�$OJ�
?Ԇ"Iio�!�V��u&A�f�PR�ߩ5, s���v1\  �H552B�Q2�1p0R78�P510.R0 � nel J�614Ҡ/WATUP��d8PW545*�H8R6��9VCAM�q97PCRImP\1tP�UIF�C8Q28  ingsQy0��4P� P63P @P PS�CH��DOCqVڀD �PCSU���08Q0=PqpV�EIOCr��� P5�4Pupd�PR6q9aP���PSET�p�t\hPQ`Qt�8P7�`Q�!MASK���(PPRXY䞓�R7B#POCO�  \pppb3 6���PR�Q��b1Pdy60Q$cJ539.e�Hsb��vLC�H-`(�OPL-Gq\bPQ0]`��P(`HCR��4`�S�aund�PMCISIP`e0aPle5=P9s�p(`DSW� � � qPb0`�aPa��(`P�RQ`Tq�RE`(Poa6901P<cPCM�PHc{R0@q\j23b��V�`E`�S`UPvisP`E` c�`UPc�PRS	a�bJ69�E`sFRDmPsRwMCN:eH931P�HcSNBARa�rHLB�USM�qc�Pvg52�fHTCIP0cTMIL�e"P�`�eJ �PA�PdST�PTX6p967PTEL�p��P�`�`
Q8P8$Q48>a"PP�X�8P95�P`[�9�5qqbUEC-`F;
PUFRmPfa�hQCmP90ZQVCqO�`@PVIP%�w537sQSUIzVsSX�P�SWEBIP��SHTTIPthrFQ62aP�!tPG����cIG؁�`c�P;GS�eIRC%��c'H76�P�e Q�Qr|�Ror��R51P0 s:P�P,t53=P8u)8=Py�C�Q6]`0�b�PI��q52]`sJ56E`s���PDs�CL�qPt5�\r�d�q75UP cR8䀑�u5P sR55 ]`,s� P8s��P�`pCP�PP�SJ77P0\o�6��cRP,P�cR6�ap�`�Q�taT�79P`�64̑Pd87]`�d90�P0c��=P,���5�9,ta�T91P� ��p1P(S���Qpai�P�06=P- C�PF��T	���!aLP PT�S�pL�CAB%�I БIQ` ;�H�UPoPaintPMS�P�a��D�IP|�STY�%�t\patPTO��b�P�PLSR76č`�5�Q��WaNNn�Paic�qNNE`��ORS�`�cR6�81Pint'�FC�B�P(�6x�-W`M��r��!(`OBQ`p�lug�`L�aot �`OPI-���P�SPZ�PPG�Q7v�`73ΒPRQ�ad�RL��(Sp�PS��n�@�E`o�� �PTS-�ǈ W��P�`ap�w�`��P`cFVR��PlcV3D%�l�PsBVI�SAPL�Pwcyc+PAPV1��pa_�CCGIP �- U��L�Prog+PCCR�`�ԁ�B�P �PԁK=�"!L�P��p��(h�<�AP��h�̱�@g�Bـ�
TX�%���CTC�ptp��2��P927"0ҝPs2��Qb��TC-�rmtl;�	`#1ΒTC9`nHcCTE�Perj�]EIPp.p/�E�P��c��I�use��F�ـvrv�F%���T�G�P� CP��%�d u-h�H-�Tra�PgCTI�p��TL� TRS���p�@נ���IP�PTh�M%�l�exsQTMQ`ve#r, �p�SC:���F��Pv\e�PF�IPSV"+�H�$cj�ـ;tr�aCTW-����CPVGF-��SVP=2mPv\fx���pac�b��e��bVP4яfx_m��-��SVsPD-��SVPF�P�_mo�`V� cV֣�t\��LmPov�e4��-�sVPR��\|�tPV�Qe5.W`V6�*u"��P}�po`���`��CVK��2N�IIP��CV�����IPN9�Gene ���D��D�R�D�����  ��f谔�po{s.��inal��n��DeR���`���d�P��omB���o�n,���R�D�R��\���TXf��D$b��o;mp�� "N��P2��m���! ��=�C-f����=FXqU�����g F��<(��Dt II��r4�D��u�� "����Cx_ui X������f2��h	C�rl2��D,r9ui��Ԣ� it2cl�0co��e"�����ا(.)�� ���� ��{� IQnQ ��I[ ��_�= wo��,b{D� ��|�GG� �����4 �e�� vʷ� ���&� 2��Z� uz������� ��TW&q�~q 5�׷&��o? ;0���  �2� ㉻y� ���W&����� ?�3�� A��e�/�> �\�3&T�{�� 77߸ ����� ���ݵ ֵ��&��{8 �l1���S�) ���d� *J� F'{s ~��� 6w:0� ��,���s�- Q�v�� ��� ��,�T �ZBLnx6���6 ��6w���Par ���s>�E��j�6d;sq��F  ����8���ЁDhel���x��ti-S�0� �Ob��Dbcf�OX�����t OFT��P<A�_�V�ZI� �D��V\�qWS��=� dtle�Ean�(bzd��tit)v�Z�z�Ez XWO H6�6����5 H�6H691b�E4܀TofkstF\� Y682�4�`n�f804�E91�g�`30oBkmon_��E��eݱ�� ql]m��0 J�fh��}B�_  ZDTf�L0�f(P7�Ec�klKV� �6|��D8q5��ّ�m\b��p��xo�k�ktq���g2.g���yLbmkLVts��IF��bk������Id #I/f��GR� �han�L��Vy��%��%ere������io�� ac�-� A�n�h���c�uACl�_�^ir���)�g��	.�@�& yG��R630�� �p v�p�&H�f��3un��R57v�O�JavG�`Y��o;wc��-ASF��`O��7���SM������
af��rSafLa�vl�\F c�w a���?V�XpoV �30��NT; "L�FFM��=�@���yh	a�G-�w�� �m2.�,�t�<�̹�6ԯ��sd_�MC'V����qD���fslm��isc.  ?H5522���21&dc.pGR78����0��708J61�4Vip A�TUu�@�OL�54]5ҴINTL�6�t�8 (VCA����sseCcRI��ȑ��UI��n�rt\rL�28gn��NRE��.f,��63!��,�SCH��d Ek�DOCV����p��C,�<�L�0�Q�isp��EIO��xE,�54���ѽ9��2\sl,�S�ET���lр�lt�2�J7�Ռ�MASK��̀OPRXY҇��7��n�OCO��J6l��3�l�� (SV�l�A�H�L�@Օ��5�39Rsv���#�1��LCH���OwPLGf�outl�q0��D��HCR
svg��S@�h��cCSa�!�{�50���D�l�5!�lQ��DS�W��S����̀��OiP����7��PR����L�ұ�(Sgd����PCM���R-0 \s��5P՝��0���n�q� A�J�1��N�q�2��P�RSa���69�� �(AuFRDx�Խ��RMCN����93A�ɐC�SNBA�F9� HLB��� M��4����h�2A�95z�H�TCaԈ�TMIL�6�j95,��85�7.,PA1�it�o��TPTXҴ �JK�TEL��pi�L�� XpL�80�I�)��.�!��P;�J9=5��s "N����H�UEC��7\c�s�FR��<Q��C��57\{VCOXa�,���IP1jH��SUI�	CSX|1�AWEBa���HTTa�8�R6%2��m`��GP%��IG %tutKIgPGSj�| RC1w_me�H76��:7P�ws_+�?�x�R51�\iw0�N���H�53!���wL�8!�h�R66 ��H���Ԡ���@;J56��1���N0���9�j��L���RQ5`%�A|�5q�r�`b,�8 5��{165!�d�@�"5��H84!�C29��0��PJ����n B[�J77!Ԩ�R6�5h3n���2y36P��3R6��-`�;о Ԩ@��ex�eKJ87��#J;90!�stu+�~@n!䬵�k90�kop�B����@!�p�@|BA�g*�n@!Ԍ�Q��06!�@[�F��FaP�6��́,�T�S� NC[�CA�B$iͰl1I��R�7��@q�y�CM]S1�rog+QM��� �� TY$x�CTOa�nv\+��1�t(�,�6�con��~0��15��JNN��%e:��P��9OR�S%x���8A�81]5[�FCBaUnZQ��P!��p{��CMOmB��"G��OL���x�OPI�$\lr"[�SŠ�T	D7�U��oCPRQR9RL���S�V�~`���K�ETS�$1��0��p�3�Ԩ�FVR1�LZQV3D$ ���sBVa�SAPL1�7CLN[�PV��	r�CCGaԙ��CL��3CCRA�n �"W!B�H�CSKQn\0�p��)��0CTPn�ЌQe���p!$bCt�aT80U�pCTC�y�:�RC1�1 (�s���trl,�r��
T�X��TCaerrm�r�MC"�s��#wCTE��nrr�R�Ea�XPj�^��r#mc�^�a"�P�Q�F!$���$p "��rG1�tTG$c�8��QH�$SCTI��! s��CTLqdACK�Rp)��r]La�R82��M��0YPk�.���OF��.���e�{�CN���^�1�"M�^�a�С�Q�`US��!$��M�QW��$m�VGF�$R� MH��P2�� H5� ΐq��ΐ�$�(MH[�VP�uo�Y����$)��D��h�g��VPF��"MCHG̑`e!�+�V/vpcm�N��ՙ�N��$�VPRqd)��CV�x�V� "�X��,�1�($TIa�t\�mh��K��etpK�A%Y�VP%ɠ�!�PN���GeneB�rip����<8��extt���Y�m�"�(�� HB���)��x��������Ȣ�reCs.�yA�ɠn� ���*���p�@M�<_�NĀ6L���8�Ș�yAvL�Xr��Ȉ2��"R;�Ƚ\�ra��	P�� h86��Gu+ʸ�Ͽ��SeLɨm�9�69 �P�Ȩr�Ȩ2�ɹ1��n2�h� �0L�XR}�RI{�e� L�x����c�Ș���N�vpx�L��"��2\r� ]�N�82�d���b@�ɉa��y1��/�k�@8���A��ruk�ʘ �L�sop��H�}�t!s{�����s��9���j965��Scx��h��5 J9��{�
�PL�J	ee�n��t I[
x�c�om��Fh�L�4 �J��fo��D�IF+�6�Q����rGati|��p��1�0&�
R8l߾�M�����P��8� �j�mK�X�HZ����IN�oڠ��3�qf��vi���80�~�l Sl�yQ��#tpk�xb�j�.� @�R�d������,/n(�8�8�0���
:�aO8�<�Q}�CO�ں�PT��O (��.��Xp|�~H���?�7v �wv��8��22�pm���722��j7�^�@ƙ�f��cf�=Yvr���vcu���O�O@�O�O_#_5_7�3Y_΋�wv4{_�_w<�ʈ�ust_�_�cus�_�Z��oo�,o>oPo�io��ngqe��(pLy747�j�WelʨHM47ZKEq {���[m�gMFH�?�(wsK� 8J�n���o���fhl;��wmfD���? :�}(4	<�g J{��II)�̏މw��X�774�kﭏ/7ntˏ݊e�+���se�/�aw���8�ɐ��EX \�!b+: �p��~�00��nh�,:Mo+�xO���1 "K�O��\a��#0��.8���{h�pL?�j+�mon�:2��t�/�st�?-�w�:���)�;��(8=h�;
d Pۻ��{:  ��� X�J0��re�����STD�!treLANG��x�81�\tqd��������rch.�������htw�v�WWָ� R�79��"Lo�51 (�I�W�h�՜��4�aww� r�vy �623c�wh a?�cti�֐�!�X�iؠ�t ��n,�։�����j��"AJP�@�3p�vr{�H�6z��!��- SeT�� E3�) G�J93�4��LoW�4 (�S������ <���9c1 ��8!4�j9�搉�+���y�
��	�b]tN�ite{�R  ��I@Ո�����P��������	 ����Z�vol��X ��9�<�I�Lp���ld*���FՇ864{��?��K��	�k扐�֘1�wmsk��M�q�Xa�e�����p��0RBT�1k�s.OPTNЦqf�U$ RTCamT��y��U��y��U��UlU6 L�T�1Tx����SFq�Ue�6T��U�SP W�b DT�qT2h�T�!/�&+��TX�U\j6�&�U U�UsfdO&�&ȁT����662DP�N�bi��%�Q�%62V��$���%�� �#�(�(6To6e St�%��#5y�$�.)5(To�%tT0�%�5�W6T���%�#�#orc��#I���#���%cct�6ؑ?�{4\W6965"p6}"�#\j536��8�4�"�?kruO O�,Im?Np�C �?tx�0<O�;�e �%����?
;gcJ7 "�AV�?�;avsf`�O__&_8WtpD_DV_0GT�F|_:UcK6�_�_r�O�3e\s��O2^y`O:�mig:xGvgW! m�%��q!�%T�$E A{60�po6��#37N�)5CR5_2E���$0��.�$Ada�Vd���V��?;Tz7�_�e7DD!TF9���#8�`�%���4y�ted� Z@�A}�@�}�04�N�}�}���}�dcH& }����u 6�vp��v1�u1\b�u�$2}���}� R83��u�"}��"}�val!g���Nrh�&��8�J�Y�o�ue��� �j70�v=1��MI=G�uerfa��{�q���E�N�ء��E{YE�ce A�� �񁏯pV�e�A!���2�Յ�Q�%��u1�e�i �@��H�e����J0�� '��b��T��E In�B�  W�|���537g����(KMI�t�Ԇr��ݟ�am���nеvi!g�U -�v J߆�8⹖F���P�y�ac����2���Rɏ jox��2�� djd�<8r}� og\k�0r��g��wmf�wFro/� Eq'�<4"}�3 J8��oni[��ᅩ}���� o� ��ʛ��Im@�R�e��{n�Є��V�o������ w ����裆"POS\����ͯ� menϖ�⑥O�Mo�43��� �(;Coc� An[�t���"e�a\�vp�ֽ.��cflx$�l�e��8�hr�tr�N�T� CF+�x �E/�t	qi�M�ӓx1c��p�f�lx����Z�cx��
0 h�כh8��mo��=� �H���)� (�vSER,���g�0߆0\r�vX�= ��I n� - �ti���H��VC�828b�5��L"�RC��Gn G/���w�P�vy�\v�vm "oƀlϚ�x`��=e�ߠ-�R-3?������v<M [�AX/2�)�.S�rxl�v#�0���h8߷=� RAXB�A�����9�H�GE/Rצ����h߶'"RXk��F�˦;85��2L/�xB�885_�q�Ro�0siA��5\rO�@9�K��v����8���.�n "�v��88��8s�i ?�9 ƀ�/�$�y O�M�S"���&�9R �H74&�`�745��	p��p��ycrI0C�c�hP0� j��-�a%?o��6D950�R7trl��ctlO�APC���j��ui"�L���  �.���^棆!�A�ѪqH��&-^7��� ��6s16C�q�794h����� M�ƔI���99��(���$FEAT_AD�D ?	����Q%P  	�H._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�`�r������� ��������&8 J\n���������TDEM�O fY   WM_� �������/ /%/R/I/[/�//�/ �/�/�/�/�/�/?!? N?E?W?�?{?�?�?�? �?�?�?�?OOJOAO SO�OwO�O�O�O�O�O �O�O__F_=_O_|_ s_�_�_�_�_�_�_�_ ooBo9oKoxooo�o �o�o�o�o�o�o >5Gtk}�� ������:�1� C�p�g�y�������܏ ӏ���	�6�-�?�l� c�u�������؟ϟ� ���2�)�;�h�_�q� ������ԯ˯ݯ��� .�%�7�d�[�m����� ��пǿٿ���*�!� 3�`�W�iϖύϟ��� ��������&��/�\� S�eߒ߉ߛ��߿��� ����"��+�X�O�a� ������������� ��'�T�K�]����� ������������ #PGY�}�� ����L CU�y���� ��/	//H/?/Q/ ~/u/�/�/�/�/�/�/ ???D?;?M?z?q? �?�?�?�?�?�?
OO O@O7OIOvOmOO�O �O�O�O�O_�O_<_ 3_E_r_i_{_�_�_�_ �_�_o�_o8o/oAo noeowo�o�o�o�o�o �o�o4+=ja s������� �0�'�9�f�]�o��� ������ɏ�����,� #�5�b�Y�k������� ��ş����(��1� ^�U�g����������� ����$��-�Z�Q� c������������� � ��)�V�M�_ό� �ϕϯϹ�������� �%�R�I�[߈�ߑ� �ߵ���������!� N�E�W��{���� ���������J�A� S���w����������� ��F=O| s������ B9Kxo� �����/�/ >/5/G/t/k/}/�/�/ �/�/�/?�/?:?1? C?p?g?y?�?�?�?�? �? O�?	O6O-O?OlO cOuO�O�O�O�O�O�O �O_2_)_;_h___q_ �_�_�_�_�_�_�_o .o%o7odo[omo�o�o �o�o�o�o�o�o*! 3`Wi���� ����&��/�\� S�e����������� ���"��+�X�O�a� {����������ߟ� ��'�T�K�]�w��� �������ۯ��� #�P�G�Y�s�}����� ���׿����L� C�U�o�yϦϝϯ��� �����	��H�?�Q� k�uߢߙ߫������� ���D�;�M�g�q� ����������
�� �@�7�I�c�m����� ����������< 3E_i���� ���8/A [e������ ��/4/+/=/W/a/ �/�/�/�/�/�/�/�/ ?0?'?9?S?]?�?�? �?�?�?�?�?�?�?,O #O5OOOYO�O}O�O�O �O�O�O�O�O(__1_ K_U_�_y_�_�_�_�_ �_�_�_$oo-oGoQo ~ouo�o�o�o�o�o�o �o )CMzq �������� �%�?�I�v�m���� �����ُ���;�  2�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ������������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ��������'9   :>Ugy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/� A�S�e�w��������� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/
=C6Yk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ������/�A��$FEAT�_DEMOIN [ E��q��>�}Y�INDEXf��u��Y�ILEC�OMP g�;����t�T����SETUP2 �h������  N ܑ��_A�P2BCK 1i~��  �)B�D��%�C�>��� 1�n�E����)���M� ˯�������<�N�ݯ r������7�̿[�� ϑ�&ϵ�J�ٿWπ� Ϥ�3�����i��ύ� "�4���X���|ߎ�� ��A���e�����0� ��T�f��ߊ����� O���s�����>��� b���o���'���K��� ������:L��p ����5�Y�} �$�H�l~ �1��g�� / 2/�V/�z/	/�/�/ ?/�/c/�/
?�/.?�/ R?d?�/�??�?�?M? �?q?O�?O<O����P� 2�*�.VRCO�O�0*��O�O�3�O�O�5w@P�C�O_�0FR6�:�O=^�Oa_�KT ���_�_&U�_�\h�R_<�_�6*.FzOo"�1	(SoEl�_io�[STM �b�o�^�+P�o�m�0iP�endant POanel�o�[H�o� �g�oYor�ZGIF|��e�Oa��ZJPG �*��e`���z��JJS��ĭ��0@���X�%
�JavaScri3ptُ�CSʏ1���f�ۏ %Ca�scading �Style Sh�eets]��0
A�RGNAME.D)T���<�`\��^����Д៍�АDISP*ן���`$�d���V�e��CLL�B.ZI��=�/`:�\��\�����C?ollabo鯕�	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V����zό�!ߘ�TPEI?NS.XML(�@��:\<����Cus�tom Tool�bar}��PAS�SWORD���>�FRS:\��� �%Passwo�rd Config��?J���C��"O ��3�����i����"� 4���X���|����� A���e�����0�� Tf�����O �s��>�b �[�'�K�� �/�:/L/�p/� �/#/5/�/Y/�/}/�/ $?�/H?�/l?~??�? 1?�?�?g?�?�? O�? �?VO�?zO	OsO�O?O �OcO�O
_�O._�OR_ d_�O�__�_;_M_�_ q_o�_�_<o�_`o�_ �o�o%o�oIo�o�oo �o8�o�on�o� !��W�{�"� �F��j�|����/� ďS�e��������� T��x������=�ҟ a������,���P�ߟ 񟆯���9����o� ���(�:�ɯ^��� ��#���G�ܿk�}�� ��6�ſ/�l������ ����U���y�� ߯� D���h���	ߞ�-����Q߻��߇��,��$�FILE_DGB�CK 1i������� ( �)
SU�MMARY.DG<,���MD:`�����Diag Summary�����
CONSLO�G��y����$����Console �log%���	TPOACCN��%g������TP AccountinF����FR6:IP�KDMP.ZIP�����
��)����E�xception�-����MEMCH�ECK������8�Memory �Data��L�N�)�RIPE����0�%�� Packets LE���$Sn�STAT*#�� %LS�tatus�i	FTP�/�/��:�mment �TBD=/� >�)ETHERN�E�/o�/�/��?EthernU<�?figuraL��~'!DCSVRF1/�/)/B?�0 v�erify alylE?�M(5DIFF:? ?2?�?<F\8diff�?}7|o0CHGD1�?8�?�?LO �?sO~3&�
I2BO)O;O��O bO�O�OG�D3�O�O�OT_ ��O{_
VUPDATES.�P�_��?FRS:\�_�]���Update?s List�_���PSRBWLD.CMo���Ro�_�9�PS_ROBO�WEL^/�/:GI�G��o>_�o�G�igE ��nos�ticW�N�>��)�aHADO�W�o�o�ob�S�hadow Ch�ange��{8+"rNOTI?�=O��Not�ific�"��O��A�PMIO �o��h��f/��o�^7U�*�UI3�E��W��{�UI���� ��B���f��_����� ��O���������>� P�ߟt������9�ί ]�򯁯�(���L�ۯ p������5�ʿܿk�  Ϗ�$�6�ſZ��~� �wϴ�C���g���� ��2���V�h��ό�� ����Q���u�
��� @���d��߈��)�� M���������<�N� ��r����%�����[� ���&��J��n ��3��i� �"�X�| ��A�e�/� 0/�T/f/��//�/�=/�/�/�$�$FI�LE_�PPR�P���� �����(MDON�LY 1i5�  
 �z/Q?�/ u?�/�?�?t/�?^?�? O�?)O�?MO_O�?�O O�O�OHO�OlO_�O _7_�O[_�O_�_ _ �_D_�_�_z_o�_3o Eo�_io�_�oo�o�o Ro�ovo�oA�o ew�*��`�����&�O��*VISBCK,81;3*.VDV�����FR:\o�ION\DATA\���/��Visi�on VD filȅ��&�<�J� 4�n������3�ȟW� �����"���F�՟� |������m�֯e��� ���0���T��x��� ���=�ҿa�s�ϗ� ,�>���b���ϗ� ��K���o��ߥ�:����^����ϔ��*MR�2_GRP 1j�;�C4  ;B�}�	 71�������E�� E��  F@ F��5U������L����M��Jk��Lzp�JP���Fg�f�?ǀ  S����9��Y9}�9���8j
�6̿�6�;��Ag�  ���BH��[B���B���$�������������@UUU#�����Y� D�}�h����������������
C��_C�FG k;T �M���]�N�O :
F�0� � \�RM_�CHKTYP  �0�}�000���OM_MIN�	x���50]X� SSBdl5:0��bx��Y���%TP_D�EF_OW0x�|9�IRCOM���$GENOV_RD_DO*62n�THR* d%�d�_ENB� ��RAVC��mK�� ��՚�/�3�/��/�/�� [�M!OUW s�܋}��ؾ��8�g�;?�/7?Y?�[?  D�C�����(7�?�<B�?B�����2��*9�N SMTT#t[)��X}��C�f�HOSTC�d1ux��\�?�� MCx��;�zOx�  2�7.0�@1�O  e�O�O	__-_;Z �O^_p_�_�_�LN_HS�	anonymous�_�_�_oo1o yO��FhFk�O�_ �o�O�o�o�o�oJ_ '9K]�o�_� ����4o�Xojo G�~�o^�������ŏ �����1�T�� �y����������� ,�>�@�-�t�Q�c�u� ��������ϯ��� (�^��M�_�q����� ܟ� �ݿ��H�%� 7�I�[Ϣ�ϑϣϵ� ���l�2��!�3�E� Wߞ���¿Կ����
� ������/�v�S�e� w����������� ��+�r߄ߖ�s��� ���߻���������� '9K]����� ����4�F�X�j� l>��}���� ��//1/T� �y/�/�/�/�/.D\A�ENT 1v
;� P!J/?  ��/3?"?W??{? >?�?b?�?�?�?�?�? O�?AOOeO(O�OLO ^O�O�O�O�O_�O+_ �O _a_$_�_H_�_l_ �_�_�_o�_'o�_Ko ooo2o{oVo�o�o�o �o�o�o5�oY�.�R�v��z?QUICC0���3��t14��"�����t2��`�r�ӏ!?ROUTERԏ���#�!PCJO�G$���!19�2.168.0.�10��sCAMP�RTt�P�!d�1m�����RT폟������$NAME �!�*!ROBO����S_CFG �1u�) ��Auto-s�tartedFTP&��=?/ ֯s����0�B�� f�x���������S�� ����,�������� �ϼ�ޯ��������� ʿ'�9�K�]�oߒ�� �߷��������� (:~�k�Ϗ��� ���������1�C� f���y����������� �,�>�R�?��c u��`����� (�$M_q� ����� /H %/7/I/[/m/4�/�/ �/�/�/�~/?!?3? E?W?i?����?�/ �?/�?OO/O�/�? eOwO�O�O�?�ORO�O �O__+_r?�?�?�? �O|_�?�_�_�_�_o �O'o9oKo]ooo�_o �o�o�o�o�o�oF_X_ j_~ok�_��� ���o���1�T U��y���������U��)�_ERR w�3�я�PDUSI�Z  g�^�p����>�WRD �?r�Cq�  �guest b�Q�c�u�������"��SCDMNGRPw 2xr�����Cqg�\�b�K�� 	P01.�00 8(q  � �5p�5pz�}5pB  �{� ���H����L��L��L�����O8�����l������a4� x��jȤ�x��8���\�U��)�`�;��#�����d�.��@�R�ɛ_GROU�ېy�����	�ӑ���QUPD � ?u����İT�Yg����TT�P_AUTH 1�z�� <!i?Pendan��-��l���!KAREL:*-�6�H͇KC]�m��U��VISION SET���ϴ�g�G�U� �����R�0��H�B߀��f�x��ߜ߮���C?TRL {�����g�
S�FF�F9E3��AtF�RS:DEFAU�LT;�FAN�UC Web Server;�)�� ��9�K��ܭ����������߄WR_CONFIG |ߛ� ;��IDL_CPU_PCZ��g�B�Dpy� BH_�MINj�)�}�?GNR_IO���g���a�NPT_SOIM_D_������STAL_SCR�N�� ���TPM?ODNTOL������RTY��y����F �ENO���Ѳ]�OLNK 1}��M�������|�eMASTE���ɾeSLAVE �~��c�O_CcFGٱBUO�|O@CYCLEn�>T�_ASG 19ߗ+�
 �� ��//+/=/O/a/�s/�/�/�/�/��N�UM��
@I�PCH�^RTRY_CNZ���@P�������� @kI�+E�z?E��a�P_MEMBE�RS 2�ߙ� 5$���2���ݰ7��?�9a�SDT_I�SOLC  �����$J23_D�SM+�3JOB�PROCN��JOmG��1�+�d8�?��+D�O�/?
�LQ�O __/_�OS_e_w_�_`�O Hm@��E#?>&BPOSREQO��?KANJI_����a[�MON ����b�yN_goyo@�o�o�o�Y�`3�<�� ��e�_ִ��_L����"?`EYLO�GGINLE��������$LANGUAGE ��<T� {q�LeGa2�	�b���g��xP��  �J�g�'��b����>�MC:\RSCH\00\<��XpN_DISP �+G�J��O�O߃gLOCp�Dz����AsOGBOOK �������������X����� Ϗ����a�*��	p�����!�m���!���=p_BUFoF 1�p���2F幟���՟D�� Collaborativǖ��� F�=�O�a�s������� ֯ͯ߯���B�9��K���DCS �>z� =���'�f���?ɿۿ���H@{�I�O 1�� ~?9ü��9�I�[�m� �ϑϣϵ��������� �!�3�E�Y�i�{ߍ�@�߱��������E��TMNd�_B�T�f� x������������ ��,�>�P�b�t���p����L��SEVD0���TYPN�1�$6���QRS�"0&��<2FL 1�"�J0���������GTP�:pOF�NGN�AM1D�mr�tUP�S�GI"5�aO5��_LOADN@G� %�%TI~�pZUZAUN#��(MAXUALR�M�'���(��_P�R"4F0d��1�B�_PNP� V 2��C	MDR�0771ߕ�B�L"8063%�@ ��_#?�ߒ|/�C��z�6��/���/�Po@P 2��+� �ɖ	T 	t  ��/�% W?B?{?�k?�?g?�? �?�?O�?*OONO`O CO�OoO�O�O�O�O�O _�O&_8__\_G_�_ �_u_�_�_�_�_�_o �_4ooXojoMo�oyo �o�o�o�o�o�o0 B%fQ�u�� ������>�)� b�M�����{������� �Տ��:�%�^�p��S�������D_L?DXDISApB��MEMO_AP�jE ?C
 �,�(�:�L�^��p������� 1�C ����4��������4��X���C�_MSTR ����w�SCD 1���L�ƿH��տ� ��2��/�h�Sό�w� �ϛ��Ͽ���
���.� �R�=�v�aߚ߅ߗ� �߻�������<�'� L�r�]������� �������8�#�\�G� ��k������������� ��"F1jUg ������� B-fQ�u����h�MKCFG� ����/�#LT�ARM_��7"0�0N/V$� �METPUᐒ3�ퟎ�ND� ADC�OLp%� {.CMN�T�/ �%� ����.E#>!�/4�%_POSCF�'�.�PRPM�/9ST�� 1��� 4@��<#�
1�5 �?�7{?�?�?�?�?�? �?)OOO_OAOSO�O wO�O�O�O�O_�A�!�SING_CHK�  �/$MODAQ,#����.;U�DEV 	��	�MC:o\HSI�ZEᝢ��;UTA�SK %��%$�12345678�9 �_�U9WTRI�G 1���l3%% ��9o��"ocoFo5#�V�YP�QNe��:SE�M_INF 1��3' `�)AT&FV0�E0po�m)�aE�0V1&A3&B�1&D2&S0&�C1S0=�m)GATZ�o;"tH? g�a[o�xA�� z���� �o>� �o'��K��� ����я:�L�3� p�#�5���Y�k�}�� ����$�[�H���~� 9�����Ưد������ ��ӟ�V�	�z����� ��c�Կ����
��.� ��d��)�;��Ͼ� q�������˿<��� `�G߄ߖ�IϺ�m�� �ϣ����8�J��n� !ߒ�M�������h_�NITOR� G �?�[   	�EXEC1�/�2*5�35�45�55��P�7�75�85�9� 0�Қ�4��@��L� ��X��d��p��|�������2��2���2��2��2��2���2��2��22*3��3��3@�;Q�R_GRP_SVw 1��k (�A��z�4�~�Kａ������K:z�j]�Q_�D��^�PL_N�AME !3%�,�!Defa�ult Pers�onality �(from FD�) �RR2� �1�L6(L�?�,0	l d �������� //(/:/L/^/p/�/��/�/�/�/�/�/ZX2 u?0?B?T?f?x?�?�?�?�?\R<?�?�? O O2ODOVOhOzO�O��O�OZZ`\RD�?�N
�O_\TP�O :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo _)_~o�o�o�o�o�o �o�o 2DVh z�[omo���� 
��.�@�R�d�v����������Џ� �Ef  Fb� �F7���   ��!��d��@� R�6�t������l�๟ʝ�����  ݘ����"�@�F�d����� "𩯹�ݐAG�  ϩU[�$�n�B�E� �� � @oD�  �?��� �?�@��A@�;�f��FH� ;�	}l,�	 |���j�s�d�>�� ��� K(���Kd$2K ���J7w�KY/J˷�ϜJ�	�xܿ�� @I���_f�@�z���f�γ�N�������	Xl��������S��ĽÔ��I �����5���  �����A?oi#��;���� o���l� �π��-���ܛG�G�Ѳ���@n�@a �  �  ���ܟ*�͵	'�� � H�I� �  �Р�n�:�Èl�È�=��̈́�в@�ߚЕ����/������̷NP� � ',���-�@�
�@���?�=�@A���B� � Cj�a�Be�C<i��#�Bи��ee��^^ȹBР��P����0̠�����ADz՟� n�3��C�i�@�R�RиY����  �@�7 ���  ���?�ff������n� ɠ#ѱy9�G
(���I�(�@uP@~����t�t���>�����;�Cd;���.<߈<�g�<F+<L�������,�d�,�̠�?fff?��?&�&��@��@x���@�N�@�?��@T�H�� ��!-�ȹ�|�� 
`�������/ /</'/`/r/]/�/��eF���/�/�/�/@m?��/J?�(E���G�#�� F Y�T?�?P?�?�?�?�? �?O�?/OO?OeOk� �O�IQOG�?�O1?��OmO_0_B_T_������A_�_	_�_P�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�ol�o���W�����o;C�E� q�H�d��؜a@q��e��F�BµWB]��NB2�(A����@�u\?��D�������b�0��|�uR�����
x~�ؽ���Bu*C���$�)`�$ ����GC#����rAU�����1�eG��D�I�mH��� I:�I��6[F���C��I��J�:�\IT�H
~�QF�y��p���*J�/ I8�Y�I��KFjʻCe�o��s��� ��Џ���ߏ�*�� N�9�r�]��������� ���۟���8�#�\� G�����}�����گů ���"���X�C�|� g�����Ŀ������ �	�B�-�f�Qϊ�u� ���ϫ��������,� �P�b�M߆�qߪߕ� �߹�������(��L� 7�p�[����������s($���3:�����$���3���d�,�4��x@�R�wa����l�<~�wa���e����wa4 �{����@��(L:ueP�	P~�A�O�������	���� G2W}h� �����/�� �O�O7/m/[(d=�s/ U/�/�/�/�/�/?�/�1??U?C?y?�=  �2 Ef9gFb-��77�9fB)aa�)`C9A`�&`w`@ -o�?w`e�O)O�?MO�Ow`�?�?�O�O�OD�O9c?�0�A7ht4�w`w`!w`xn
 �O9_K_]_ o_�_�_�_�_�_�_�_��_o#ozzQ ���h��G���$M�R_CABLE �2�h t�a�T� @@�0`�Ae��a�a�a��`ɺ�0�`C�`�aO8��tB�n�d���`�aE�4�GE�#�o�f�#���0��0�DO���By`��Š���bED4E��c,��o�g8 [ ���C�07�d�4
vے�0 ��b��XE��Z&�l�`y`
qCܛp�bHE�
v#=g�5D�Ү�qz
�lҠ`��0�q�p�bw0�
v�%c����b=%	E;h��u/o�c-��4tH� \�?�9�K�]�o�ԏϏ ��
�ɏۏ@���?��eo �a����𪟼��b��� ����"`��( �� ������`����Ӡ���@����_����������� � ���@����*,�� ,�-�\cOM ��ii��3� � �� ��%�% 234567O8901i�{� f�H����������1�����
��`��not sent�3�����;��TESTFECSALGR  e�q�iG�1d.�š
:�� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.x�ml��ֿqta�E��DEFAUL�T-�i4\bGRP ;2�M�  =��a�4��as  �%�Force�s�or checkS  ���b�z��p����h5-[ �ϻ���������ID�%!1s�t cleani�ng of co�nt. v�ilation��}�R��+��[�ߔߦ߸�z��mech�gcal`�����!�0��h5k�@��R�d�v����(�rolle_Ƶ����/���(�:�L���Basic q�uarterly�������,������0�����M��:C@"GpP�a�b`i4�������#AC���M"��{�Pbt���S�uppq�greaCse���?@/&/8/J/\/��C+ �ge��. batBn�y`/��/h5	/ �/�/�/? ?_�ѷen'�v��/�/��/��?�?�?�?�?ѣG=?O�qp"CrB1O��0�/`OrO�O��O�O�t$��Lf�B�C-m��A�O:�OO@$_6_H_Z_l_�t*�cabl�Om���B�S<m��Q�_:�
_ �_�_oo0oo)(Ӂ/�_�_���_�o�o�o��o�o�O@ha�u1�l�2r xm�<qC:��op������ReplaW�fUȼ2�:�._4�F�X�j�|�m�$%���o�������#� ��
��.�@���d��� ŏ׏����П���� U�*�y�����r����� ����	�q��?�߯c� 8�J�\�n���ϯ���� �ڿ)����"�4�F� ��jϹ�˿������� �����[�0�ϑ�f� �ϊߜ߮�����!��� E�W�,�{�P�b�t�� ���߼�����A�� (�:�L�^�������� ������� $s� H������q��� ��9]o�V hz���U�# �G/./@/R/d/� �/�/��//�/�/? ?*?y/N?�/�/�?�/ �?�?�?�?�???Oc? u?JO�?nO�O�O�O�O+J�r	 H�O�O_ _6M2_@OBE:_p_>_ P_�_�_�_�_�_ o�_ �_oHoo(oZo�o^o po�o�o�o�o�o �o� :z �bA?�w  @�q _ ���Fw�� ��H* �**  @q>v�p2T�f�x�:�p������ҏ��eO ^C7�Տ#�5�G�	�k� }���ُ���c���� �W��C�U�g���ß )�����ӯ���	�� -�w�����9��������m�Ͽ��=�O�E�	A�$MR_HI_ST 2�>uN��� 
 \�$Force� sensor �check  1�23456789�0q�3����ß��N}SB�� -319.8 �hours RU�N 9.�Y�!1�st clean�ing of c�ont. ven�tilation 0ÄϖϨ�O�*�<� � Or߄ߖ�M�_߹� ���ߧ����8�J�� n�%���[������ ���"���F�X��|��3�����i�����:�S�KCFMAP  ]>uQ��r�5�������ON�REL  .��3���EXCFEN��:
��Q�FNCXJJOG_OVLIM8dN�\� ��KEY8�=�_PAN7�P���������SFSPDTYP8xC��SIG�:>��T1MOT�G���_CE_GRoP 1�>u\�D�����/� ���/�/U// y/0/n/�/f/�/�/�/ 	?�/???�/c??\? �?P?�?�?�?�?�?O�)OOMO,���QZ_�EDIT5 )T�COM_CFG 1���[�O�O�O� 
�ASI ��y3�
__+[_O_��>O�_bH�T_ARC_U�.Ń	T_MN_M�ODE5�	U?AP_CPL�_g�NOCHECK {?�� �� o.o@oRodovo�o �o�o�o�o�o�o�*!NO_WAI�T_L4~GiNTƑA���EUwT_7ERRs2���3���ƱJ�����X>_)��|MO�s��}�x:Ov���8�?����� l��r_PARAM�r�����j���5�<5�G� =  r�b� t�s�X�������������֟�0�����b�t�����SUM_?RSPACE������Aѯۤ�$ODR�DSP�S7cOF�FSET_CAR8t@�_�DIS���PEN_FILE�:�7�AF�PTION_IO��q��M_PRG %���%$*����M�W�ORK �yf ��춍��"��������	 ������gT���RG_DSBL'  ��C�{u���RIENTTO�7 ��C� A� �UT_SIM�_Dy���V~�LCT ��}�{B �٭��_PEX��P=��RAT�W �dc��UP S���`���e߰w�]ߛߩ��$�2�r�L6(L�?���	l d ������&�8�J�\� n��������������"�4�F�X���2 �߈�������������*�<w�Tf x�������8J`�ˣ@G���Tz�Pg ������/"/ 4/F/X/j/|/�/�/�/ ���/�/??0?B? T?f?x?�?�?�?�?�? �?�?�/�/,O>OPObO tO�O�O�O�O�O�O�O�__(_:_��O�!�y_�]2ӆ��_�^ �_�_�W^]^]��/ooSog�Hgrohozo �o�o�o�o�oF`�|#|`�A�  9y�����OK�1��k������<�EA��nq @D�  Ђq����nq?��C���s�q1� ;�	}l��	 |�Q��s�r�q>���u �sF`H<z�H~�H3k7�GL�zHpG�99l7�k_B�LT�F`C4��k�H����t��-�Ae��¾k�����s���  �ሏ�����EeBVT���d}Z�����ڏ ���q-�Fk��y�{FbU����n@6�  ����z�Fo��Be	�'� � ���I� �  y�:p܋=���ڟ웆�@���B�,���B���g�Ag9N����  '|����g��B��p�B�ӀC׏����@  �#�Bu�&�e{e�^^މB:p2���>�m�6p�Z���Dz?o}�܏�� ����׿������Ǒ���� f�  � ��M���*�?�faf�_8�J�ܿ 3pϑ�ñ8�Чϵʖq$.·�(����P��ɐ'��s�tL�>��/�;��Cd;��.<�߈<�g�<F+<L ��^o�iΚrd@��r6p?f7ff?�?&�п��@��@x���@�N�@���@T싶�Z���� �tމ�u�߈w	�x��t i�>�)�b�M��q�� ������������:� %�^�������W���S�E�  G�aF�� Fk����� ����1U@yd ������q��	 ��{�A��h�����a��ird��A{/w/J/5/n/
vA��A���":t�/� C^/�/Z/ ލ?���/�/1??��K�W����g��p�E� ~1�?04�80
1�1@IӀ���BµWB]�N�B2�(A���@�u\?����������b�0��|�uR�����
�>�ؽ����Bu*C���$�)`�? ����GC#����rAU�����1�eG����I�mH��� I:�I�6[F���C4O�I��J�:\�IT�H
~Q�F�y�Ol@��*J�/ I8Y��I��KFj��C��-?�O�O__ >_)_b_M_�_�_�_�_ �_�_�_o�_(oo%o ^oIo�omo�o�o�o�o �o �o$H3l W�{����� ��2��V�h�S��� w�����ԏ������� .��R�=�v�a����� ��П����ߟ��<� '�`�K�]��������� ޯɯ��&�8�#�\�z�3(J���3:a�������J�3��pc4���������<���1����ڿ��1���e���14 �{2�2�r�`Ϡ�τϺϨ��%PR�P���!�h�!�K�x6�o�Z�����u� |ߵߠ���������� 3��W�B�{�f�4���������d�A���� !��1�3�E�{�i��������������  2� Ef�7Fb�7��6B�!�!� KC9� �� �0@�/ `r������#x��+=�3Q?, V�8v��0��0��0�.
 D����� //%/7/I/[/m//��/�:� ��ֻ��G���$PAR�AM_MENU �?2���  DE�FPULSE�+�	WAITTMO{UT�+RCV?� SHELL�_WRK.$CU�R_STYL� �4<OPTJJ?P�TB_?Y2C/?R_DECSN 0�Ű< �?�?�?�?�?OO?O :OLO^O�O�O�O�O�O��!SSREL_IOD  .�����E�USE_PROG %�*%�O0_�CCCR0�B���#CW�_HOST !F�*!HT�_=ZT��O_�Sh_zQ�S�_<[_TIME
2�FXU�� GDEBUG��@�+�CGINP_�FLMSKo5iT�RDo5gPGAb` 2%l�tkCHCo4h�TYPE�,�  �O�O�o#0Bk fx������ ���C�>�P�b��� ������ӏΏ���� �(�:�c�^�p������7eWORD ?	��+
 	RS�c`��PNS���C4�JOv1��TyE�P�COL��h��2��gLP 3������OjTRACECTL 1�2Ż�! �� �Қ�q�_DT Q�2�Ǡ���D � :m����Ԡ�Ԡ��}�hׯ���;�4� �4��4���;�u:�Pq:���;�8�	8�U
8�8�8�8�E8�8��@:�8�8���� ���*ٱ޴���ؿ �$�6���
�l�~�@� R�dϞϰ��������� 
��V�h�zߌߞ߰� ��������
�,�>�P��*�<�v��*� +�8� (��)��* ����������)�;� M�_�q����������� ����%,�>�P� b�t������������ С�*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6@ubt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀�V�߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h?�z?�?�?�?�?�1�$�PGTRACEL�EN  �1  ���0���6_UP �/���A@�1�@�1_CFG7 �E�3�1U
@�<D�0<D�ZO<C�0uO$BDEF�SPD �/L��1�0��0H_C�ONFIG �\E�3 �0�05d�D��2 �1�AaPpDsA�A�0��0�IN'@TRL ɽ/MOA8pEQPEv�E��G�A�<D�AILID(C��/M	bTGRP 1}ýI l�1�B  ������1A�33FC�� F8� E�� @eN	�A�AsA�Y��Y�A�@� 	 �vO�Fg�_ ´8cokB;`baBo,o�>oxobo�o�1>о�?B/�o�o~��o =%<��
C@yd ��"������  Dz@�I�@A 0�q� �������ˏ�� �ڏ���7�"�4�m��X���|���Ú)ґ�
V7.10be�ta1HF @�����Aq�ܢQ  �?�� �BܠP�p �C���&�B�EQ�A���Q�P�Q�� @ß[�m����<CA���0�b�@���f�������ҡ�R�ܣ�R����1�i������t<B!CeQ�KNOW_M  �lE7FbTSV ĽJ�BoC_�b� t�������������1��]aSM�SŽK ���	NB�0����ĿK���-�bb��A�R� �P����0�Ŗ��bQ+MR�S��T�iN�`��d���V]ST�Q�1 1�K
 4aMU�iǨj� K� ]�oߠߓߥ߷����� ��2��#�h�G�Y�� }�������
������,�27�I��1�#<t�H��P3^�p�����,�4���������,�5(:,�6 Wi{�,�7����,�8�!3n,�MAD�6 F�,�OVLD  �KD�xO.�PAR?NUM  �MC\/%�SCH� E�
9'!G)�3Y%UP�D/��E�/P�_C�MP_��0@�0'�7E�$ER_CH�K�%5H�&�/�+RqS���bQ_MO��+?=5_'?O�_RES_G6��:�I�o �?�?�?�?O�?O7O *O[ONOOrO�O�O�{4]��<�?�Oz5�� �O__|3 #_B_G_ |3V b_�_�_|3� �_ �_�_|3� �_�_o|3�Oo>oCo|2V 1��:�k1!�@c?��=2THR_IN�Rc0i!}�o5d�fM�ASS�o Z�gM�N�o�cMON_QUEUE �:ը"�j0��O�N� U�1Nv�+DpEND8Fqd?`yEXEo`uƅ BEnpPAsOP�TIOMwm;DpPR�OGRAM %�$z%Cp}o(/BrT�ASK_I��~O?CFG �$���K�DATA��&T���j12/ď ֏������+�=�O� a����������͟���INFO�͘�� 3t��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����
�Θ� '��FJ�a K_N��T��˶�ENBg ڽw1��2���GN�2�ڻ� P(O�=�{��]ϸ�@���v� �u�uɡd�Ʒ_EDIT ��T�����G�WER�FL�x�c)�RGA�DJ Ҷ�A�  $�?j00��a��Dqձӆ5'�?��ʨ�<u�)�%e������FӨ�2Y�R��	H;pl�G��b_�>�pAodɻt$�*�/� **:�j0�$�@�5Y�T���^��q�߈b~�L��\� n���������� �����4�F�t�j�|� ������������b LBT�x�� ��:��$, �Pb���/� ���/~/(/:/h/ ^/p/�/�/�/�/�/�/ V? ??@?6?H?�?l? ~?�?�?�?.O�?�?O O O�ODOVO�OzO�O _�O�O�O�O�Or__ ._\_R_d_�_�_�_�_�_�_�f	g�io�pWo �o{d�o�~o�ozo�B�PREF S�Rږp�p
�?IORITY�w[�}��MPDSP�q���pwUT6����OoDUCT3������OG��_T�G��8��ʯrTOE�NT 1׶� �(!AF_IN�E�p,�7�!t�cp7�_�!u�dN���!ic�mv��ޯrXYK��v����q)� ,�����p��&�	� �R�9�v�]�o����� П������*��N�`�*�sK��9}�ߢ�\��Ư ,�/6�H�������خ�At�?,  �Hp���P�b�t����u�w�HANCE �R��:�wd��连�2s��9Ks��POR_T_NUM�s�p����_CAR�TREP{p�Ω�SoKSTA�w dʷLGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_a_seiban�o \��olߒ�}߶ߡ��� ������"���X�C� |�g���������� ���	�B�-�f�Q��� u������������� ,<bM�q� ������(|L�VERSIyp��w} di�sabledWS�AVE ߾z	�2600H76%8S?�!ؿ����/ 	5(�r)og+^/y�e{/�/�/��/�/�*�,/? ��p���_�p 1��Ћ� ������Wh?z?�W*pURGE��B�p}vgu6,�WF�0DO�vƲ©vW%��4(�C�WR�UP_DELAY� �\κ5R_HOT %Nf�q׿�GO�5R_NORM�AL&H�r6O�OZGS�EMIjO�O�O(qQ/SKIPF3��W3x=_98_J_\_] �_�_{_�_�_�_�_�_ �_	o/oAoSoowoeo �o�o�o�o�o�o�o +=aOq�� ������'���7�]�K�������)E�7$RA{���K/��zĀÁ_PARA�M�A3��K @�.�@`�61�2C�<��y��C��6$�BÀBTIF��4`�RCVTMO�Uu�c��ÀD�CRF3��I ��+Q;/�CC�SeD�#�1�=h�-0�t�]�/��ޅ��{���1�0��_���k_���Cd;���.<߈<��g�<F+<L����Ѱ��d�u� L�������ϯ�����)�;�M�_���RD�IO_TYPE � M=U�k�EFP�OS1 1�\�
 x4/����� +�$/<��$υ�pϩ� D���h��ό��'��� ���o�
ߓ�.ߤ�R� ��������5���Y� ��i��*�<�v���r� ��������U�@�y� ���8���\������������?��c����2 1�KԿX��T�x��3 1����nY�>S4 1�'9�K�/�'/�S5 1���/�/��/�/:/S6 1� Q/c/u/�/-??Q?�/S7 1��/�/
?�D?�?�?�?d?S8 1�{?�?�?�?WOBO�{O�?SMASK �1L��O�D�GX�NO���F&�^��M�OTEZ�Ż��Q_�ǁ�%]pA݂��P?L_RANG!Q]��_QOWER ��ŵ�P1VSM_D�RYPRG %�ź%"O�_�UTAR�T �^�ZUME_PRO�_�_4o���_EXEC_E�NB  J�e�GSPD`O`WhՅjbgTDBro�jRM�o��hINGVERS�ION Ź�#o�)I_AIR7PURhP �O(.�MMT_�@T�P#_�ÀOBOT_I/SOLC�NTV@Az'qhuNAME�l���o�JOB_OR�D_NUM ?��X#qH7�68  j1Zc�@�r
�rV��s��r�?��r?�r�pÀP?C_TIMEu�a��xÀS232>R1��� LT�EACH PEN�DANw�:GX��!O Main�tenance /Consj2�����"��No UseB�׏������p1�C�y�V�NPO�P\@�YQ�cS�oCH_L`�%^� �	ő��!U�D1:럒�R�@VGAIL�q@�Ӏ�J��QSPACE1 ;2�ż ��YR s�i�@Ct�YRԀ'{~��8�?�� ˯����"���7�2� c�u�����G���߯ѿ 򿵿�(��u�AC� c�u�����Ͻ�߿�� �ϵ��(��=�_�q� �ϕ�C߹������߱� �$��9�[�m�ߑ� ��Q������߭��� � ��	�W�i�{���M� ������5���. S�e�w�����I���� ���*?a s��E���� �/&//;/]o� �����/2/�/? "?�/7?Y/k/}/�/�/ O?�/�/�?�?�?O0O�OKA��*SY�PpM*�8.30�261 yB5/2�1/2018 gA �WPfG|�H��_TX`� !$�COMME��$USAp �$ENABLE=DԀ$INN`QpgIOR�B�@RY�E?_SIGN_�`�A�P�AIT�C�BWR�K�BD<�_TYP<�CRINDXS�@�W�@%VFRI{�_�GRPԀ$UF�RAM�rSRTOO}L\VMYHOL�A�$LENGTH�_VTEBTIRS�T�T  $S�ECLP�XUFIN�V_POS�@�$MARGI�A�$WAIT�`�ZX�2�\�VG2�GG1��AI�@�S�Q	g�`_�WR�BNO_USE�_DI�BuQ_RE�Q�BC�C]S$CUR_TCQP�R"a�^f �GP_ST�ATUS�A @� �A3`�BLk�HE$zc1�h�P@���@}_�FX �@�E_MLT_CTf�CH_�J�`CO�@�OL�E�CGQQ$�W�@w�b#tDE�ADLOCKuD�ELAY_CNT��a3qGt�a$wf _2 R1[�1$X<�2[2�{3[3$Zwy�q%Y�y�q`%V�@�c�@�b$V�`�RV�UV3oh>b�@ � �d�0ar'MSKJ�LgWaZ��C`NRK�PS_RATE�0$���S
`�Q�TAC��PRDH���e�S*��a4�b�  �DG�A 08�P�flp bquS�2ppI�#`
`�P� 
�S\` � �A�R_ENB�Q �$RUNNER_AXI��<`ALPL�Q�RU�T�HICQ$FL�IP7��DTFER�EN��R�IF_C	HSU�IW��%V)�CG1����$PřA�Q��Pݖ_JF�P�R_P�	�RV_�DATA�A � $�ETIM|���$VALU$��	�OP_  � �A  2� �SC*��	� �$IT�P_!�SQ]PNPOU�}�o�TOTL�o�D�SP��JOGLI�b��PE_PKpc�O�f�i��PX]PTA�S�$KEPT_GMIR��¤"`M�b&�APq�aE�@��y�q�g@١c�q�PG�BRK6�x���L�I��  ?�SJ��q�P�ADEz�ܠB�SOCz�MOTN�v�DUMMY16�Ӂ$SV�`DE�_OP��SFSP�D_OVR
��f�@LD����OR��[TP8�LE��F��l����OV��SF��F����bF�d�ƣ&c�)�fQc�LCHDL}Y��RECOV���`��W�PM��gŢ�#RO������_F�?�� @v�S �NVsER�@�`OFS�PC,�CSWDٱc�ձ����B����TRG�|š�`E_FDO���MB_CM}���B��BLQ�¢	�Q�̄Vza�BUP�g��G
��AM���@`�KՊ�e�_M!�d�A�Mf�Q��T$CAԕ���DF���HB�Kd�v���IOU2��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�y3A��ATIO�0��͠��US����WaAB��R+c�`t��`DؾA��_AUX~w�SUBCPUP���S�`����3Եжc8���3�FLA�B�HW_Cwp"�Ns&��]sAa��$UN�ITS�M�F�AT�TRIz�Z�CY{CL�CNECA����FLTR_2_�FI��TARTU�PJp����A��LPx������_SCT*cF_F�F_P���b��FS��+�K�CHA�/Q��*�d�RS�D��Q����Q���_TH�PROr���հGEMPJ���G�T�� �Q�D�I�@y�RAILAiC/�bMX�LOf�xS��ځ���拁��V��PR#�S`appz�C� 	���FUNC���RI�N`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ngDAQ�B�rkLD�र&q�M�K���TI���j���$�@RIA_[SW��AF��Pñ#��%%�p9r1���MOIQ���DF_l~P(�PD"LM-�{FA�PHRDY�DORG�H; _QP|�s%MULSE~P�z���*�� J��J�ײ��FAN_A�LMLVG��!WR=N�%HARDP���UcO�� K2$SHADOW]�kp�a802��� STOf�+�Y_^�w�AU{`R<��eP_SBR�z5����:F�� �3MPINF?�\�4�λ3REGV/1DG��+cVm �C�CFL4(��?�DAiP���Z`�� �����Z�g	 �P(Q$�A$Z�Q V�@�[��
� ��EG0߀o���kAAR�����2�axG��AX�E��ROB��RE%D��W�QD�_�Mh�CSYA��AF��FS�G�WRI�P~F&�ST�R����E�˰EH�H)��D�a\2kPB6P��=V��Dv�OTOr�1)���ARYL�`tR�v�3���FI&�~ͣ$LINKb!�\��Q�_3S��8�E��QXYZ2�Z�5�VOFF���R��R�XxPB��`ds�G�cFI�0�3g�������_J��'�ɲ�S&qR0LT2V[6���aTBja�"2�bC���DU�F]7�TUR� X���e�Q�2XP�ЊgFL�E���x@�`�U9Zy8���� 1	)�%K��Mw��F9���8������ORQj��G;W3���#�Ґd ����uz����1�tOV	E�q_�M��ё?C�u EC�uKB�v'0�x-�w H��t���& `��q ڠ�B�ё�u�q�wh�0ECh����ER��K�	�EP����AT�K�6e9e�W���AXs�'��v� /�R ����!��  ��P��`��`�3p�Yp�1�p�� � � �� (�� 8�� H� � X�� h�� x�� �������DEBU��$%3�I��·RA!B���ٱ�sV��� 
d�J、��@� ����������Q���a ���a��3q��Yq+$�`�%"<�cLAB0b8�u�'�GRO���b<��B_s��"T ҳ*`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Q`θuݸ��PNT0~���SERVE �NZ@ $`EAV�!�PO�����nP!�P@�$!Y@�  $>�TREQ�b
=��BG�K��%"2\��� _ � l��5�D6ESRRVb(�I��V0`�;���TOQ:�7�L��@
�R��e G�%ĩQ�� <�50F� �,�`�z�>�RA~� 2 d!�2����S�  M�`�pxU ����OCu�G�  ��C�OUNT6Q��FZ�N_CFGF� 4#��6��TG4�_��=�����Î�VC ���M �"��$06��q ��FA E� &��X�@������$�A����AP��P@�HEL�0��� 5b`B_BA�S��RSR�6"�CSH����1�Ǌ�U2��3��4��5��6��7��8��}�R�OO����P�PNL�EA�cAB)ë ��A[CKu�INO�T���(B$UR0� =�_cPU��!0��OU+�Pd�8j��� V���TPFWD_KA1R��� ��RE(ĉ qP�P�>QUE�:�RO�p�`r0P1I � x�j�P�f��6�Q�SEM��0��� An��STYL�SO j�DIX�&������S!_TMCMANsRQ��PENDIt�$KEYSWI�TCH���kH}E�`BEATM83PE{@LE��>]�J�U��F��Sp�DO_HOM# Ol�@�EF�pPRaPB�A#PY�C� O�!<���OV_M|b<0 IOCM�dFQ���h�HKYA# D�Q�7��UF2���M���p�cFOR�C�3WAR�"�O}M|@  @S�T#o0U)SP�@1�U2&3&4E���*T�O��L���8OUNLOv�D4K$�EDU1  �S�Y�HDDNF� �M�BLOB  �p�SNPX_;AS�� 0@�0|��81$SIZ�1�$VA{���MU/LTIP-��# �A� � A$��� /4`�BS���0�C���&FRIF�BO�S���3� N=F�ODBUP߰��%@3;9(��ҋ�Z@� x��SI��TE�s�r�cSGL�1T�Rp&�Н3B��@�0OSTMTq�3Pg@�VBW�p�4SHO�W�5@�SV��_�G�� 3p$PC�J�PИ���FB�PHSP AW�EP@�VD�0WC� ���A00��PB �XG XG XG$ XG5�VI6VI7VI8VI9
VIAVIBVI�XG�YF�0XGFVH��XbIU1oI1|I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1Y1Y2UI2bIU2oI2|I2�I2�I@�`�X�I2p�X�I2�IU2�I2�I2�I2Y�2Y�p�hbI3oI3�|I3�I3�I3�I3��I3�I3�I3�I3��I3�I3�I3Y3�Y4�i4bI4oI4�|I4�I4�I4�I4��I4�I4�I4�I4��I4�I4�I4Y4�Y5�i5bI5oI5�|I5�I5�I5�I5��I5�I5�I5�I5��I5�I5�I5Y5�Y6�i6bI6oI6�|I6�I6�I6�I6��I6�I6�I6�I6��I6�I6�I6Y6�Y7�i7bI7oI7�|I7�I7�I7�I7��I7�I7�I7�I7��I7�I7�I7Y7ZTҁVP� UD�#y"ՠ��
<A62���t�R��CSMD� ��M5�Rv�,]��Q_h�R���pe����<�YSL��>�  � �%\2 ��+4�'��W�BVALU��b��'�z��FH�ID_L����HI��I���LcE_��㴦�$0�RD�SAC�! �h �VE_B�LCK��1%�D_CPU5ɧ 5ɛ ������C�� ��R �" � PW�j��#0��LA�1�SBћì���RUN_FLG�Ś�����@� ����������H����Х���TBC2���# � @ B ��e �S�8=�F'TDC����V���3d�Q�THF�����R�L�ESERCVE9��F��3�2��E��Н�X -$��LEN9��F���f�RA��W"G�WI_5�b�1��д2�MO-�T%S60U�I�k�0�ܱF����[�DyEk�21LACEi�0�CCS#0�� _M�A� j��z��TCV����z�T�������.Bi�'A�z�'AJ$h�#EM5���J��@@Ri�V�z���2Q `�0&@o�h��JK��VK9��{���щ�J0����JJ��JJ��AAL���������4��5�ӕ NA1������.�LD�i_�1�CF�"�% `�GROUP���1�AN4�C�#~m REQUIR�ҎEBU�#��6�$Tk�2$���z�я #�& \�A�PPR� C� 0�
�$OPEN�CLOS�St��	i�
��&' �M�fЩ���W"-_MG�7CB@�A����BBRK@NOL�D@�0RTMO_�5ӆp1J��P ��������������6��1�@ ��Р�#�(�# �����'��+#PATH''@!6# @!�<#� � '��1�SCA���6I�N��UCJ�[1� C0@UM�(Y ��#�"������*���*��� P�AYLOA~J2=LؠR_AN^�3�L��91�)1AR?_F2LSHg2B4LO4�!F7�#T7�#ACRL_�%�0ȏ'�$��H��.�$yHA�2FLEX�u�J!�) P��2�D߽߫�v �2��* :����z�FG�]D����z���%�F1]A�E�G4�F�X�j�|���BE������ ������(��X�T*� A���@�XI�[�m�\At�T$g�QX<�=�� 2TX���emX������ ������������t+	
"J>+ �-�`K]o|�٠AT�F�4�ELFPѪs��J� *� JEmC3TR�!�ATN�v�zHAND_VB�.��1��$, $�8`F2Av���S�Wu�-� $$M*0.�]�W�lg��PZ����A@��� 1����:AK��]AkAz��LTN�]DkDzPZ G��C�ST_K�lK�N}DY��� A ����0��<7]A<7W1@�'��d�@g`�P� ������"�J"�. M�2D%"�H����ASYM$j%0�� j&-��-W1�/_�{8� �$������/�/�/�/ 3J�<�:9�/�89�D_�VI�v����V_UNI�ӛ��cD1J����╴�W<��n5 Ŵ�w=4��9��?�?$<�uc�4�3�
!%�H���/�j��0��DIzuO�Ķ8
!k�>0 �`��I��A��#���@ģ����@��HQl� �1 � /�MEB.Qp��9�ơT}�PT�;pG �+ GtA� ���'��T��0 $DUM�MY1��$PSm_�@RF�@  G �b�'FLA@ Y�P(c|��$GLB_TP�ŗ���p9 P�q��2 X� �z!ST9�� S�BRM M21_V��T$SV_ERb*0O�p����CL�����AGPO��f�GLv~�EW>�3 4H ��$YrZrW@�x�A1+�A���"jк �U&�4 8`N�Z�"�$GI�p}$&� -� �Y��>�5 LH {��}�$F�E��NEA�R(PN�CF��%PT�ANC�B;�JOG܌@� 6.@$JOINTwa?pd��MSET>�7  "x�E��HQtpS{r��|up>�8� �p�U.Q?�� LOC�K_FOV06���B�GLV�sGLt�T?EST_XM� 3�'EMP����Ҏ_�$U&@%�w`24� Y��5��2�d���3��CE- ����_ $KAR�QM��TPDRA)������VECn@��IUھ�6��HEf�TO�OL�C2V�DREN IS3ER6�N�@ACH� 7?1Ox �Q�29Z�H �I�  @$R�AIL_BOXEzwa�ROBO���?��HOWWA�R�1�_�zROLMj��:qw�jq� ��@ O_Fkp!� d�l>�9�� +�R O8B: �@d�;�"�OU�	;�Һ�3ơ�r�q_�_$PIP��N&`�H�l�@��#@CORDEDd�p >�f�fpO�� < 7D ��OB⁴s d���Kӕ���qwSYS�ADR�q�f��TCHt� 7= ,8`ENo��1Ak�_{�-$Cq_��f�VWVA��>� �  &��P�REV_RT��$EDITr&VSHWRkq�֑ &RJ:�v�D��JA�$~�a$HEAD�h6�� �z#KE:�E�CPSPD�&JKMP�L~��0R*PF��?��1%&I��5S�rC�pNE; �q��wTICK�C��M��13�3HN��@� @� 1Gu�!_GqPp6��0STY'"xLO��:�2l2?�_A t 
m G3%S%$R!{�=��S�`!$��w`���ճ�r��Pˠp6SQU��x�E��u�TERC��0��TSUtB ����hw&`gw�Q)b�pO����@IZ��4{��^�PR�kј�B1XPU���E_�DO��, XS�KN~�AXI�@���UR�pGS�r� ^0�d&��p_) �ET�BQPm��o��0Fo�2�0A|���Rԍ���a;�SR�Cl>@P��b_�yU r��Y��yU��yS��yS ���UЇ�U���U���U �]��Ul[��Y�bXk�]Cm�����YR�SC�� D h��DS~0��Q�SPL���eATހ���A�]0,2N�ADDRE�S<B} SHIF�{s��_2CH�pr�I��=q�TVsrI��E"���a�Ce�
��
c�VW�A��'F \��q��0l|\A@�rC�_B"R{z�p�ҩq�TXSCWREE�Gv��1TINA���t{��c��A�b?�H T 1�ЂB�����I��Ap��BE�y RRO������� B���4�UE�4I �g�!p�S���RSM]0�GU�NEX(@~Ƴ�j�S_S�ӆ��Á։񇣣��ACY�0� 2-H�pUE;�J���\��@GMT��Lֱ��A��O	�BBL�_| W8���K �Լ0s�OM��LE�/r��� TO!�s�RwIGH��BRD
�%qCKGR8л�T�EX�@����WIDTH�� �B[�|�<���I_��Hi� OL 8K���_�!=r���R:�_���Y�SC�O6q�M�g0紐U��h�Rm��LUMh��FpGERVw �P����`�N��&�GEKUR��FP)�)� �LP��(RE%@�a)�ק�a�!��f �5*�6�7�8Ǣ#B@�É@���tP�fW��S@M�USR�&�O <����U8�Qs�FOC)��PRI;Qm� :����TRIP�m�SUN����Pv��0���f%��'���@�0 �Q����AG ��0T� �a>q�OS�%�RPo���8�R/�A�H�L4����	U¡�SU�g��¢�5��OFF���T��}�O�� 1�R�����S�GU�N��6�B_S�UB?���,�SRT�N�`TUg2��mCO9R| D�RAUrPE�yTZ�#'�VCC���	3V AC36�MFB1�%d�PG� �W (#��ASTEM�����0�PE��T3G�X y�\ ��MOVEz�A��AN�� ���|M���LIM_X�� 2��2��7�,�����0ı�
�BVF�`EӐ��~��04Y��IQB�7���5S��_Rp� 2��� WİGp+@��}СP��>3�Zx ����3���A�ݠCZ�DRID���ѡVy08�90� De�MY_UBYd���6��@��!��X��GP_S��3��L�K�BM,�$+0DE�Y(#EX`�����U/M_MU� X����ȀUS�� ���G0`PACI���а@ ��:��:,�:����CRE/�3qL�+���:[��TARG"��P�r��R<��\ d`��A��$�	4��AR��SW2 ��-��@Oz�%qA(7p�yREU�U�01�Z,�HK�2]g0��qP� N� �E9AM0GWOR��ާMRCV3�^ U���O�0M�C�s�	���|�REF _���x(�+T� �� �������3_RCH4(a�P�Ѐ��hrj�NA�5��0�_ ��2����L@��n�@@OU~7w6���Z��a2[��R1E�p�@;0\�c�a�'2K�@SUL��]2��C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��PQ5I�]7q�}�Tg`�4D`�0.`0�APg_HUC�5SA��CMPz�F�6�5�5
�0_�aR��a�1I�\!X�9��VGFS���ad ��M8��0p�UF_x��B� �ʼ,RO��Q��'l����UR�3GR�`.�3IDp���)��D�;��A��~�IN"��H{D���V@AJ���S͓UWmi`=�����TYLO*��5�D����b�t +�cPA�= �cCACH�vR��UvQ��Y��p�#CZF�I0sFR�XT����Vn+$HO��� �P!A3�XBf�(1 ���$�`VPy� ^bO_SZ313he6K3he12J�eh chG�6chWA�UMP�j���IMG9uPAD<�iiIMRE�$�b/_SIZ�$P�����0 ��ASYNBU=F��VRTD)u5t�qΓOLE_2DPJ�Qu5R��C��U���vPQuECCUlVEMV �U�r�W�VIRC�aIuVTPG���rv1s��5qFMPLAqa��v����0�cm� CKLAS�	�Q�"���d  �ѧ%ӑӠ@�}¾�$�Q���Ue A|�0!�rSr�T�# 0! �r�iI��ml�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f �� >֦3�@Sp�SgLOW>�RO��ACCE���!� 9��VR�#���p:���A1D�����PAV�j��� D����M_B8"���^�JMPG ���g:�#E$SSC@��F�vPq��hݲ�vQS�`qVN��L;EXc�i T`�s�r���Q�FLD �DEsFI�3�0p2���:��VP2�V�j� �A��V|�4[`MV_PIs���t���A�@��F	I��|�Z��Ȥ����`�A���A��~�GAߥ�1 LOO��1 JC�B���Xc��^`�#P�LANE��R��1F@�c�����pr�M� [`�噴��S����f� ���Af��R�Aw�״t9U��pRKE��d��VANC�OO��V���� k����ϲ�R_AA� l��2� ��p�#HĎ��m h�@��O K��$������kЍ0O)U&A�"A�
p�p�SK�TM@FVIEM 2l ��P=���n <<��dK�/UMMYK1P���`D��AC�U��#AU��o �$��TIT�g$PR����OP���VSHIF�r�p`J�Qs�ؙ�fOxE$� _R�`U�#����s��q ������G�"G�޵'�9T�$�SCO{D7�CNTQ i�l�>a� -�a�;�a�H�a�V����1�+�2u1��D�����  � S�MO�Uq��a�J,Q�����a_�R[�ir�n�*@LIQ��AA/`�XVR��s��n�TL���ZABC�t�t�c�]
AZIP��u撖��LVbcLn"�^��MPCFx�v:��$�� ���DMY_LN�������@y�w Ђ(a�u� �MCM�@CbcCA�RT_�DPN� �$J71D ��=NGg0Sg0�B�UXW� ��UXE#UL|ByX@���	��|!Z��x 	���m��YH�Db  y �80���0EIGH��3n�?(� H����$z ���|������$B� Kd'��_X��L3�RVS�F`���OVC�2' �$|�>P&��
q����5D�TR�@ �V:�1O�SPHX��!�{ ,� *<��$R�B2 2 ����C!�  �@ V+| b*c%g!H�b)g"��`V*�,8�?�V+�/V.�/�/ ?�/�/V(7%3@/R/ d/v/�/6?�/�/�?�?@�?O4OOION;4]? o?�?�?�?SO�?�?�O�_�O0_Q_8_f_N;5 zO�O�O�O�Op_�O_ o8o�_MonoUo�oN;6�_�_�_�_�_�oo %o4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8����� Ǐ=�_�n���R���şx��ڟN;G � џ�
�� ����W�i�{����� ��ï�.�������A��dW�<�N�|� ������Ŀֿ�ޯ� ��0�B�_�R�d�� �϶������������ �*�L�^��rτ�
� �����������&�p8�J�l�~� `ҟ @�з��������-����&�,� ��9�{�����a��� ������������A 'Y����� ����a#�1�
��N;_MO�DE  ��S ��[�Y�AB���
/\/*	|/��/R4CWORK_{AD�	��T1/R  ���� ��/� _INTVA�L�+$��R_O�PTION6 ��q@V_DAT�A_GRP 2,7���D��P�/~? �/�?�9��?�?�?�? OO;O)OKOMO_O�O �O�O�O�O�O_�O_ 7_%_[_I__m_�_�_ �_�_�_�_�_!ooEo 3oioWoyo�o�o�o�o �o�o�o/e S�w����� ��+��O�=�s�a� ������͏���ߏ� �9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_T�IM����ΑR� ��Ƙ/��5�;#�U!P"�Z����  �?E�W�i�{�����.��ïկ�����'(~�T"2F���dR�I�Y��2�o+@a얿����)�u���� k0ϴ��_ ��  T� � ��2�D�)�T D��Q�zόϞϰ����� ����
��.�@�R�d��v߈ߚ�/V凷�����߽��B�_;�o �W��p��
�t���Diz$� �0 � �T"%!��� ������������ ��*�<�N�`�r��� ������������ &8J\n��� �����"4FX ��࿁�� �����/`4� =/O/a/s/�/�/�/�/ �/�/�!!/ �0޲k� ݵu�0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ ok$o6oHoZo lo~o�o�o�o�o1/�o �o 2DVhz �/5?������ ��&�8�J�\�n��� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-��?�Q�c�u��� �� ��`Ò�ϯ���� )�;�M�_�q������� ��˿ݿ� ����\3� ���&2,���	12345�678v�h!B_!��2�Ch���0�ϵ����� �����!�3�9ѻ�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� h�K߰���������
� �.�@�R�d�v����� ���������* <N`r���� ���&��J \n������ ��/"/4/F/X/j/ |/;�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�/�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_�? L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o=_�o�o�o�o�o �o 2DVhz@�����h��� ���u�o.�@�R���Cz  B��_   ���2&�_ � _�
����  	�_�2��Տ����_�p������ďi�{� ������ß՟���� �/�A�S�e�w����� ����N������+� =�O�a�s��������� Ϳ߿���'�9�K�"_������<v�_���$SCR_GR�P 1
� ��� t ���� ��	 �����������������_������)�a�����&�DE� D�W8���l�&�G��CR-35iA �90123456�7890��M-�20��8��CRg35 ��:�
��D�������������:֦�Ӧ�G���&������	��]�o������:���H���>��������@���&���ݯ:���j����g������B��t����������A����  @�`��s@� ( ?�=���Ht�P
��F@ F�`z�y� ����� �$ H��Gs^p��B��7�� /�0//-/f/Q/�/ u/�/�/�/8���P�� 7%?����"?W?-2<?<���]? �H�1�?t�ȭ7@�������?-4A, ��&E@�<�@G�B-1 3OZOlO-:HA��H�O�O|O P��B(�B�O�O_��E�L_DEFAUL�T  �����`SHO�TSTR#]A7RM�IPOWERFL�  i�/UYTW7FDO$V /UR�RVENT 1�����NU L�!DUM_EI�P_-8�j!AF_INE#P�_-4O!FT�_->�_r;o!��`o �*o��o!RPC_M'AIN�ojh�vo�oN�cVIS�oii��o�!TPpPU��Ydk!
P�MON_PROX	Yl�VeZ�2r���]f��!RD�M_SRV��Yg�O�!R��k��XYh>���!
�`M���\i���!RL�SYNC�-98|֏3�!ROS�_�-<�4"��!
C}E4pMTCOM����Vkn�˟!	��C'ONS̟�Wl����!��WASRCd��Vm�c�!��'USBd��XnR��� Noӯ�������!���E��i�0���WRV�ICE_KL ?�%�[ (%S?VCPRG1��-:"Ƶ2ܿ�˰3�	�"˰4,�1�˰5T�Y�"˰6|ρ�˰7�ϩϐ˰�����9���� ȴf�!�˱οI�˱�� q�˱ϙ�˱F���˱ n���˱���˱��9� ˱��a�˱߉��7� ���_������� ��)����Q����y� �'���O����w� �������� ˰��İd�c��� ���=(a s^������ /�/9/$/]/H/�/ l/�/�/�/�/�/�/�/ #??G?2?k?V?}?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O��O�O�O	_�O-_��_�DEV �Y��MC:5Xd��GTGRP 2�SVK ��bx 	�� 
 ,�PK 5_�_�T�_�_�_ o�_'o9o o]oDo�o hozo�o�o�o�o�o �o5{�_g�� �������� ?�&�c�u�\������� Ϗ���J\)���M� 4�q���j�����˟ݟ ğ��%���[�B� �f������ٯ���� ���3��W�i�P��� t���ÿ���ο�� �A�(�e�L�ί��R� ���ϸ������ �� O�6�s�Zߗߩߐ��� �������'�~ϐ�]� ��h�������� �����5��Y�@�R� ��v���������@�	 ��?&cu\� ������� ;M4qX���� ���/�%//I/ [/B//f/�/�/�/�/ �/�/�/�/3??W?� L?�?D?�?�?�?�?�? O�?/OAO(OeOLO�O �O�O�O�O�O�O�O_�iV �NLy�6� * 		S=>��+c"_VU@T�n_Y_B���B��2�J�j~Q��~_g_�_�Q%J?OGGING�_�^�7T(?VjZ�R{f��Y���/e�_%o7e�Tt�]/o�o {m�_�o�m?Qi�o�o�;)Kq%� �o�}os���� ��9�{`��)��� %���ɏ���ۏ�S� 8�w��k�Y���}��� ş���+��O�ٟC� 1�g�U���y������ �'����	�?�-�c� Q���ɯ����w���s� ���;�)�_ϡ��� ſOϹϧ�������� �7�y�^ߝ�'ߑ�� �ߣ��������Q�6� u���i�W��{��� ���=��M���A�/� e�S���w�������� ����=+aO ������u�� �9']��� M������/ 5/w\/�%/�/}/�/ �/�/�/�/=/"?4?�/ ?�/U?�?y?�?�?�? ?�?9?�?-OO=O?O QO�OuO�O�?�OO�O _�O)__9_;_M_�_ �O�_�Os_�_�_o�_ %oo5o�_�_�o�_[o �o�o�o�o�o�o!co H�o{��� ���; �_�S� A�w�e�������я� ��7���+��O�=�s� a������П���� �'��K�9�o����� ��_���[�ɯ���#� �G���n���7����� ����ſ����a�F� ���y�gϝϋϭϯ� ����9��]���Q�?� u�cߙ߇ߩ���%��� 5���)��M�;�q�_� ���߼��߅������ %��I�7�m������ ]�����������! E��l��5��� ����_D� we����� %
//���=/s/ a/�/�/�/��/!/�/ ??%?'?9?o?]?�? �/�?�/�?�?�?O�? !O#O5OkO�?�O�?[O �O�O�O�O_�O_sO �Oj_�OC_�_�_�_�_ �_�_	oK_0oo_�_co �_so�o�o�o�o�o#o Go�o;)_Mo ����o��� �7�%�[�I�k���� ������ُ���3� !�W���~���G�i�C� ���՟���/�q�V� �����w�������� ѯ�I�.�m���a�O� ��s�������߿!�� E�Ͽ9�'�]�Kρ�o� ������Ϸ���� 5�#�Y�G�}߿Ϥ��� m���i������1�� U��|��E����� ����	���-�o�T��� ���u����������� G�,k���_M� q����� ��%[Im� ��	���// !/W/E/{/��/�k/ �/�/�/�/	???S? �/z?�/C?�?�?�?�? �?�?O[?�?RO�?+O �OsO�O�O�O�O�O3O _WO�OK_�O[_�_o_ �_�_�__�_/_�_#o oGo5oWo}oko�o�_ �oo�o�o�oC 1Sy�o��oi� ����	�?��f� x�/�Q�+���Ϗ��� ��Y�>�}��q�_� ������˟���1�� U�ߟI�7�m�[�}�� ��ǯ	��-���!�� E�3�i�W�y�ϯ��ƿ ��������A�/� eϧ���˿UϿ�Q��� ������=��dߣ� -ߗ߅߻ߩ������� �W�<�{��o�]�� ��������/��S� ��G�5�k�Y���}��� ������������C 1gU������{ ����	?-c ���S���� ��/;/}b/�+/ �/�/�/�/�/�/�/C/ i/:?y/?m?[?�?? �?�?�?? O??�?3O �?COiOWO�O{O�O�? �OO�O_�O/__?_ e_S_�_�O�_�Oy_�_ �_o�_+oo;oao�_ �o�_Qo�o�o�o�o �o'ioN`9 ������A&� e�Y�G�i�k�}��� ��׏���=�Ǐ1�� U�C�e�g�y����֟ ���	���-��Q�?� a���ݟ��퟇��ϯ ��)��M���t��� =���9���ݿ˿�� %�g�Lϋ���mϣ� �ϳ�������?�$�c� ��W�E�{�iߟߍ߯� �����;���/��S� A�w�e��������� �����+��O�=�s� �����c��������� ��'K��r��; �������# eJ�}k�� ���+Q"/a� U/C/y/g/�/�/�// �/'/�/?�/+?Q??? u?c?�?�/�?�/�?�? �?OO'OMO;OqO�? �O�?aO�O�O�O�O_ _#_I_�Op_�O9_�_ �_�_�_�_�_oQ_6o Ho�_!o�_io�o�o�o �o�o)oMo�oA/ QSe�����%{,p�$SER�V_MAIL  �+u!��+q�O�UTPUT��$�@�RV 2��v  $� (�q�}��SAVE�7�(�TOP10 �2W� d O6 *_�π(_� �����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u�����`����Ͽݷ��YP���'�FZN_CFGw �u$��~����GRP �2�D� ,B�   A[�+qD;� B\��  �B4~�RB2�1��HELL�!�u��j�k�2���>��%RSR���� ���
�C�.�g�Rߋ� v߈��߬�����	����-�?�Q��  �_�%Q���_�슨�,p����)ޖ�g�2,pd��ﾆ�HK 1�� ��E�@�R�d��� �������������� *<e`r���?OMM ������FTOV_EN�B�_���HOW_?REG_UI�(��IMIOFWDL� �^�)WAIT���$V1��^�NTIM���VA�_)_UNIT�����LCTRY�B�
�MB_HDD�N 2W�  2�:%0 �pQ/�qL/ ^/�/�/�/�/�/�/�/��"!ON_ALI_AS ?e�	f�he�A?S?e?w?�: /?�?�?�?�?�?OO &O8OJO�?nO�O�O�O �OaO�O�O�O_"_�O F_X_j_|_'_�_�_�_ �_�_�_oo0oBoTo �_xo�o�o�o�oko�o �o,�oPbt �1������ �(�:�L�^�	����� ����ʏu�� ��$� Ϗ5�Z�l�~���;��� Ɵ؟����� �2�D� V�h��������¯ԯ ���
��.�ٯR�d� v�����E���п��� ϱ�*�<�N�`�r�� �ϨϺ���w����� &�8���\�n߀ߒߤ� O�����������4� F�X�j�|�'����� �������0�B��� f�x�������Y����� ����>Pbt ������ (:L�p�� ��c�� //$/ �H/Z/l/~/)/�/�/ �/�/�/�/? ?2?D?�V?]3�$SMON�_DEFPRO ����1� *S�YSTEM*0�m6RECALL �?}9 ( ��}
xyzrat�e 11 >14�7.87.149�.40:1253�2 =�=3148y �1�95172]?lO+M}�561�>��?�?�?�O�O4G�66��?ZOlO~O_!_4G|?O�E2896 �O��O_�_�_8Ctp?disc 0I_[P�\_n_�_o#o6Etpconn 0�M �_�_�_�o�o�O�4Jo \ono�o#6_H_Z_ �o�o���o�?Xj |��2D��� ������T�f�x�	� �.�@�ҏ������ ,���P�b�t����)� <�Ο��������:A�8copy fr�s:orderf�il.dat v�irt:\tmpback\I�[�y��
��/L/��mdb:*.*ԯ���ؒ���7D3x��:\ H�ɰZ�[�s����(�
;@4��aǿٿV��� ϗϩϼ�ίW�r��� �'�:���^���ߓ� �߸�K�]���#� 6�����l��ߏ�ﴟ �AJ�\�n���#�6�H�844 ����� ������J�\�n���#6OHO02[�������99����I [y
/0?�� R
���8�H����Vt�/)/ }5 ?����/�/�/� �Xs�/?(?;�/ _�/?�?�?�L/^/ ��?O$O7/�?�?m/ �?�O�O�/�/P?�/}O _ _3?E?�Oi?�O�_ �_�?�?VO�?y_
oo /OAO�_eO�_+o�o�� ��Qocouo�o*=O	192^��o����B�$SNPX�_ASG 2�����q�� P 0 '�%R[1]@g1.1��y?��s%�!��E�(�:�{� ^�������Տ��ʏ� ��A�$�e�H�Z��� ~���џ����؟�+� �5�a�D���h�z��� ��ů�ԯ���
�K� .�U���d�������ۿ ������5��*�k� N�uϡτ��ϨϺ��� ���1��U�8�Jߋ� nߕ��ߤ�������� ��%�Q�4�u�X�j�� ������������;� �E�q�T���x����� ������%[ >e�t���� ��!E(:{ ^������/ �/A/$/e/H/Z/�/ ~/�/�/�/�/�/�/+? ?5?a?D?�?h?z?�? �?�?�?�?O�?
OKO .OUO�OdO�O�O�O�O �O�O_�O5__*_k_ N_u_�_�_�_�_�_�_ �_o1ooUo8oJo�o�no�o�o�d�tPAR�AM �u��q �	��jP��d9p�ht���pOFT_KB_?CFG  �c�u��sOPIN_SI/M  �{vn���p�pRVQS�TP_DSBW~�r"t�HtSR }Zy � &!p�INGS EL_O5SEM���v�TOP_ON_ERR  uCy8��PTN Zu^k�A4�R��_PR�D��`V�CNT_GP 2�Zuq�!px 	 r��ɍ���׏��w�VD��RP 1�i p�y��K�]� o���������ɟ۟� ���#�5�G�Y���}� ������ůׯ���� �F�C�U�g�y����� ����ӿ��	��-� ?�Q�c�uχϙϫ��� ��������)�;�M� _�qߘߕߧ߹����� ����%�7�^�[�m� ������������ $�!�3�E�W�i�{��� ������������ /ASew��� ����+= Ovs����� ��//</9/K/]/ o/�/�/�/�/�/�/? �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O�O)�PRG_CO7UNT8v�k�GuNKBENB��FEMpC�:t}O_UPD 1}�{T  
4O r�O�O�O__!_3_ \_W_i_{_�_�_�_�_ �_�_�_o4o/oAoSo |owo�o�o�o�o�o�o +TOas �������� ,�'�9�K�t�o����� ����ɏۏ����#� L�G�Y�k��������� ܟן���$��1�C� l�g�y���������ӯ ����	��D�?�Q�c� ��������ԿϿ�� ��)�;�d�_�q�=L�_INFO 1޵E�@ �2@���������� ��ٽ`y*�d��h'��¬߾�=`y;MYS�DEBUGU@�@���d�If�SP_PwASSUEB?xۿLOG  ��ʠC��*ؑ�  ���A��UD1�:\�ԘΥ�_MPAC�ݵE&�8�A���V� �A�SAV �!�������X����SVZ�TEM�_TIME 1"����@ 0  [X��X�X�����$T1SVGgUNS�@VE'�E���ASK_OPTIONU@�E�A�A+�_DI��qOG��BC2_GRP �2#�I�����@��  C���<Ko�C�FG %z��� q�����`�� 	�.>dO�s �������* N9r]��� ����/�8/#/ \/n/��Z+�/Z/�/�/ H/�/?�/'??K?]� k?=�@0s?�?�?�?�? �?�?O�?OO)O_O MO�OqO�O�O�O�O�O _�O%__I_7_m_[_ }__�_�_�X� �_�_ oo/o�_SoAoco�o wo�o�o�o�o�o�o =+MOa�� �������9� '�]�K���o������� ��ɏ���#��_;�M� k�}��������ß� ן��1���U�C�y� g�������������� �	�?�-�c�Q�s��� �������Ͽ��� �)�_�Mσ�9��ϭ� ������m���#�I� 7�m�ߑ�_ߵߣ��� ��������!�W�E� {�i���������� ����A�/�e�S�u� w������������� +=O��sa�� �����9 ']Kmo��� ����#//3/Y/ G/}/k/�/�/�/�/�/ �/�/??C?��[?m? �?�?�?-?�?�?�?	O �?-O?OQOOuOcO�O �O�O�O�O�O�O__ ;_)___M_�_q_�_�_ �_�_�_o�_%oo5o 7oIoomo�oY?�o�o �o�o�o3!Ci W������ ���-�/�A�w�e� ���������я�� �=�+�a�O���s��� ����ߟ͟��o�-� K�]�o�ퟓ�����ɯ��צ��$TB�CSG_GRP �2&ץ��  �� 
 ?�  6�H�2� l�V���z���ƿ��������(�d׊E+�?�	 �HC���>���G����C�  �A�.�e�q�C��N>ǳ33��S�/]���Y��=Ȑ� C\�  Bȹ��B���>����P���KB�Y�z��L�H�0�$����J�\�n�����@�Ҿ����� ����=�Z�%�7��鈴�?3�����	�V3.00.�	�cr35��	*����
�������Ƈ� 3��4�  7 {�CT�v�,}��J2�)��������CFG +�ץ'� *�������I����.<
�<b M�q����� ��(L7p[ ������/ �6/!/Z/E/W/�/{/ �/�/�/�/.�H��/? ?�/L?7?\?�?m?�? �?�?�?�? OO$O�? HO3OlOWO|O�O��� �Oӯ�O�O�O!__E_ 3_i_W_�_{_�_�_�_ �_�_o�_/oo?oAo So�owo�o�o�o�o�o �o+O=s� E���Y���� �9�'�]�K�m����� ��u�Ǐɏۏ���5� G�Y�k�%���}����� ßşן���1��U� C�y�g�������ӯ�� ����	�+�-�?�u� c����������Ͽ� ��/�A�S�����q� �ϕϧ��������%� 7�I�[���mߣߑ� �������߷��3�!� W�E�{�i����� ��������A�/�e� S�u������������� ��+aO� s��e����� 'K9o]� ������#// G/5/k/}/�/�/[/�/ �/�/�/�/??C?1? g?U?�?y?�?�?�?�? �?	O�?-OOQO?OaO �OuO�O�O�O�O�O�O ___M_�e_w_�_ 3_�_�_�_�_�_oo 7o%o[omoo�oOo�o �o�o�o�o!3�o �oiW�{��� ����/��S�A� w�e�������я���� ���=�+�M�s�a� ��������ߟ�_	� ��_ן]�K���o��� ����ۯɯ���#�� �Y�G�}�k�����ſ ׿��������U� C�y�gϝϋ��ϯ��� �����	�?�-�c�Q� s�u߇߽߫������ ��)��9�_�M���� /����i������%� �I�7�m�[������� ������������E Wi{5���� ����A/e S�w����� /�+//O/=/_/a/ s/�/�/�/�/�/�/? '?��??Q?c??�?�? �?�?�?�?�?O�?5O GOYOkO)O�O}O�O�O��O�N  �@S� V_R�$T�BJOP_GRP� 2,�E�  ?�Vi	-R4S.;\��@�|u0{SPU �>��UT� @�@LR	 ��C� �Vf  �C���ULQLQ>�33�U�R�����U�Y?�@=�Z�C��P��ͥR�>�P  B��W$o�/gC��@g�d�Db�^����eeao�P&ff�e=��7LC/kaB� o�o�P��P�ef�b-C�p��^�g`�d�o�PL�Pt<�eVC\  �Q�@�'p�`�  �A�oL`�_wC�BrD�S�^��]�_�S�`<P�B��P�anaa`C�;�`L�w�aQo�xp�x�p:���XB$'tMP@�PCAHS��n���=�P𥅡�trd<M�g E�2pb����X�	� �1��)�W���c�� ����������󟭟�7�Q�;�I�w���;d��Vɡ�U	V3�.00RScr35QT*�QT�A��� E�'�E�i�FV#�F"wqF>���FZ� Fv�R�F�~MF����F���F��=�F���F�ъ�F��3F����F�{G
�GdG��G#
�D���E'
EMK�E���E����E�ۘE����E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F���vF�u�<#�_
<t���ٵ�=�_��V� �R�p�V9� ]E_STPARtp�H�FP*SHR\�ABL/E 1/;[%�S�G�� �W�G�BG�G� WQG�	G�E
G�GȖ�QG��G�G�ܱv�RD	I~�EQ�ϧϹ�������W�O_�q�{ߍߐ�߱���w�S]�CS  !ڄ���������� ��&�8�J�\�n��� ���������� ]\�`� ��	��(�:������
��.�@�w�NUoM  �EEQ�P	P ۰ܰw�_CFG 0���)r-PIMEBF_TTb��CSo�,GVERڳ-B,�R 11;[ 8I��R�@� �@&  ����� ��//)/;/M/_/ q/�/�/�/�/�/?�/ ?J?%?7?M?[?m?> �@�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_l�_�Y@cY�M�I_CHAN8 �c cDBGLVĂ�:cX�	`ET�HERAD ?*f�\`��?�_�uo�oQ�	`ROUT6V!	
!�d�o~�lSNMASKQh|cba255.u�ߣ'9ߣY�OOLOFS_DIb���U;iORQCT�RL 2		�Ϸ~T����� #�5�G�Y�k�}����� ��ŏ׏�����.���R�V�PE_DE�TAI/h|zPGL�_CONFIG �8�	���/�cell/$CID$/grp1V�@̟ޟ����Ӏ�o ?�Q�c�u�����(��� ϯ������;�M� _�q�����$�6�˿ݿ ���%ϴ�I�[�m� ϑϣ�2��������� �!߰���W�i�{ߍ��߱�%}F�������/�A�C�i�H� Eߞ����������?� �.�@�R�d�v���� ������������* <N`r��� ����&8J \n��!��� ��/�4/F/X/j/ |/�//�/�/�/�/�/ ??�/B?T?f?x?�? �?+?�?�?�?�?OO �?>OPObOtO�O�O�O����User� View ��}�}1234567890�O�O�O_#_`5_=T�P��]_���I2�I:O�_�_�_�_�_�_X_j_�B3�_GoYo�ko}o�o�o o�op^4 6o�o1CU�ovp^5�o���� �	�h*�p^6�c� u����������ޏp^7R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3� �OM�_�q��������y  e��Yz���	�� -�?�Q���uχϙ�俀����������>�� e�5i��c�u߇ߙ߫� ��d������P�)�;� M�_�q��*�<��i� ��������)���M� _�q������������ ����<�û��=Oa s��>����* '9K]f� Q�������/ �%/7/I/�m//�/ �/�/�/n<��^/? %?7?I?[?m?/�?�? �? ?�?�?�?O!O3O �/<׹��?O�O�O�O �O�O�?�O_!_lOE_�W_i_{_�_�_FOXG9 +_�_�_oo(o:o�O Kopo�o)_�o�o�o�oP�o ��	g�0�o M_q���No� ���o�%�7�I�[� m�&l�n��Ə؏ ���� ��D�V�h� ��������ԟ柍� g�ڻ}�2�D�V�h�z� ��3���¯ԯ���
� �.�@�R���3uF�� ����¿Կ������ .�@ϋ�d�vψϚϬ� ��e�w���U�
��.� @�R�d�ψߚ߬��� ��������*���w� ��v������� w�����c�<�N�`� r�����=�w��-��� ��*<��`r ����������  ��1C Ugy�����<��    -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_��  
��(  }�%( 	 y_ �_�_�_�_�_�_o	o +o-o?ouoco�o�o�o:�Z* �Q &�J\n�� ����o���9� (�:�L�^�p������ ���܏� ��$�6� }�Z�l�~�ŏ����Ɵ ؟���C�U�2�D�V� ��z�������¯ԯ� ��
��c�@�R�d�v� ����᯾�п�)�� �*�<�N�`ϧ����� �Ϻ��������&� 8��\�n߀��Ϥ߶� ��������E�"�4�F� ��j�|������� �����e�B�T�f� x�������������+� ,>Pb��� ������� (o�^p��� ���� /G$/6/ H/�l/~/�/�/�/�/ /�/�/?U/2?D?V?�h?z?�?�/�`@  �2�?�?�?�3�7�P���!frh:\�tpgl\rob�ots\m20i�a\cr35ia.xml�?;OMO_O qO�O�O�O�O�O�O�O ���O_(_:_L_ ^_p_�_�_�_�_�_�_ �O�_o$o6oHoZolo ~o�o�o�o�o�o�_�o  2DVhz� �����o�
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ �ݟ��&�8�J�\� n���������ȯߟٯ ���"�4�F�X�j�|�@������Ŀ־�8.1� �?@88�?�ֻ�ֿ� 3�5�G�iϓ�}ϟ��� ���������5��A��k�U�wߡ߿��$T�PGL_OUTP�UT ;�!�!/ ������ ��,�>�P�b�t�� ������������ (�:�L�^�p�������������2345678901������ ���"��BT fx��4�����
}$L^ p��,>���  //$/�2/Z/l/~/ �/�/:/�/�/�/�/?  ?�/�/V?h?z?�?�? �?H?�?�?�?
OO.O �?<OdOvO�O�O�ODO VO�O�O__*_<_�O J_r_�_�_�_�_R_�_ �_oo&o8o�_�_no �o�o�o�o�o`o�o�o "4F�oT|� ���\��}���@��0�B�T�e�@�������� ( 	 ��Џ����� �<�*�L�N�`����� ����ޟ̟���8� &�\�J���n�������@��ȯ���"������ �*�X�j�F�����|� ¿Կ��C���ϱ�3� E�#�i�{�忇ϱ�S� ���������/ߙ�S� e�߉ߛ�y߿���;� ������=�O�-�s� ���ߩ��]������� �'����]�o���� ��������E����� 5G%W}����� �g���1� Ug	w�{�� =O	//�?/Q/// u/�/��/�/_/�/�/ �/�/)?;?�/_?q?? �?�?�?�?�?G?�?O �?OIO[O9OO�O�? �O�OiO�O�O�O!_3_ �O_i_{__�_�_�_��_�_�R�$TPOFF_LIM >�|op:��mq�bN_SV`  �l�jP_MOoN <6�d�opop2l�aST�RTCHK =�6�f� bVTCOMPAT-h�af�VWVAR >rMm�h1d �o� �oop`ba_�DEFPROG �%|j%ZER�O ZUZAUN�	�j_DISPL�AY`|n"rINST_MSK  t|� ^zINUSsER�odtLCK�|�}{QUICKMExJp�"rSCRE�p�6��btpscdt�q��b*��_.�ST�jiRA�CE_CFG U?Mi�d`	�d�
?�u�HNL �2@|i����k  r͏ߏ���'�9��K�]�w�ITEM �2A�� �%$�12345678�90����  =<�П��  !���p��=��c�� ^����������.� ��R��v�"�H�ί�� Я������*�ֿ�� �r�2ϖ�����4�޿ �ϰ���&���J�\�n� ��@ߤ�d�v��ς��� ���4���X��*�� @�����ߨ��� ����T���x���� ��l��������,�>� P�������FX��d ������:� p"��o��� ��F6HZt~ ��N/t/�/��//  /2/�/V/?(?:?�/ F?�/�/�/j?�??�? �?R?�?v?�?QO�?lO �?�O�OO�O*O|O_ `O _�O0_V_h_�Ot_ �O__�_8_�_
oo �_@o�_�_�_Lodo�_ �o�o4o�oXojo3�o N�or��o���s�S�B���zψ  h��z 8��C�:y
 P�v��]����UD1:�\�����qR_G�RP 1C��?� 	 @Cp� ��$��H�6�l�Z��|�����f���˟��<�ڕ?�  
�� �<�*�`�N���r��� ����ޯ̯��&��0J�8�Z���	�u������sSCB 2D� ����π(�:�L�^�pς��|V�_CONFIG E���@����ϖ��OUTPUT yF������� 6�H�Z�l�~ߐߢߴ� �����������#�6� H�Z�l�~������ ��������2�D�V� h�z������������� ��
�.@Rdv ������� )<N`r�� �����//% 8/J/\/n/�/�/�/�/ �/�/�/�/?!/4?F? X?j?|?�?�?�?�?�? �?�?OO/?BOTOfO xO�O�O�O�O�O�O�O __+O>_P_b_t_�_ �_�_�_�_�_�_oo '_:oLo^opo�o�o�o �o�o�o�o $�� ��!�bt���� �����(�:�-o ^�p���������ʏ܏ � ��$�6�G�Z�l� ~�������Ɵ؟��� � �2�D�U�h�z��� ����¯ԯ���
�� .�@�Q�d�v������� ��п�����*�<� M�`�rτϖϨϺ��� ������&�8�J�[� n߀ߒߤ߶������� ���"�4�F�W�j�|� ������������� �0�B�S�f�x����� ����������, >Pa�t���� ���(:L>/x���k} gV�K���/ /&/8/J/\/n/�/�/ �/W�/�/�/�/?"? 4?F?X?j?|?�?�?�? �/�?�?�?OO0OBO TOfOxO�O�O�O�?�O �O�O__,_>_P_b_ t_�_�_�_�O�_�_�_ oo(o:oLo^opo�o �o�o�o�_�o�o  $6HZl~�� ��o���� �2� D�V�h�z�������� ԏ���
��.�@�R� d�v���������Ϗ� ����*�<�N�`�r� ��������˟ޯ�� �&�8�J�\�n����������Ż�$TX_�SCREEN 1}Gg��}ipnl/���gen.htm�ſ�*�<�N�`Ͻ�Panel soetupd�}�d�@�Ϸ����������� ��6�H�Z�l�~ߐ�� ��+�������� �2� �߻�h�z������ 9�g�]�
��.�@�R� d������������� ��}���<N`r ��;1�� &8�\��������QȾUA�LRM_MSG k?��� � Ȫ-/?/p/c/�/�/�/ �/�/�/�/??6?)?�Z?%SEV  �-�6"ECFoG I���  ȥ@�  }A�1   B�Ȥ
 [?ϣ��?O O%O7OIO[OmOO�O��O�G�1GRP 2�J�; 0Ȧ	 ��?�O I_BB�L_NOTE �K�:T��#lϢ�ѡ�0R�DEFPRO %+ (%N?u_Ѡ c_�_�_�_�_�_�_o �_o>o)oboMo�o\�INUSER  �R]�O�oI_ME�NHIST 1L��9  (�0� ��)/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,1133,1�oDV�hz~�� }9361�����r �$�6�H�Z�l�~�� ����Ə؏����� � 2�D�V�h�z�	����� ԟ���
���.�@� R�d�v��������Я �����9Rq��B� T�f�x���������ҿ ����ϩ�>�P�b� tφϘ�'�9������� ��(߷�L�^�p߂� �ߦ�5������� �� $����Z�l�~��� ��C�������� �2� �/�h�z��������� ������
.@�� dv�����_ �*<N�r �����[�/ /&/8/J/\/��/�/ �/�/�/�/i/�/?"? 4?F?X?C�U��?�?�? �?�?�?�/OO0OBO TOfO�?�O�O�O�O�O �O�O�O_,_>_P_b_ t__�_�_�_�_�_�_ �_o(o:oLo^opo�o o�o�o�o�o�o �o $6HZl~i?{? ������2� D�V�h�z����-� ԏ���
����@�R� d�v�����)���П� ��������N�`�r� ������7�̯ޯ�� �&���J�\�n�����������$UI_�PANEDATA 1N���ڱ�  	�}�����!�3�E�W� )Y�}�7�뿨� ���������i�&�� J�\�C߀�gߤߋ��� ��������"�4��X�.7�� �q}�� ����������B�� ��%�I�[�m������ 
�����������! E,i{b������l�ܳ7� <N`r���� -���//&/8/� \/n/U/�/y/�/�/�/ �/�/?�/4?F?-?j? Q?�?�?%�?�?�? OO0O�?TO�xO�O �O�O�O�O�OKO_�O ,__P_b_I_�_m_�_ �_�_�_�_oo�_:o �?�?po�o�o�o�o�o o�o sO$6HZ l~�o����� �� �2��V�=�z� ��s�����ԏGoYo �.�@�R�d�v�ɏ�� ��П������ <�N�5�r�Y������� ̯���ׯ�&��J� 1�n�������ȿڿ ����c�4ϧ�X�j� |ώϠϲ���+����� ���0�B�)�f�Mߊ� �߃��ߧ�������� ����P�b�t���� ������S���(�:� L�^����i������� ���� ��6Z�lS�w�'�9�}���"4FX)�}��l��� ��/j'//K/2/ D/�/h/�/�/�/�/�/ �/�/#?5??Y?��C��=��$UI_PO�STYPE  �C�� 	� e?�?�2QUI�CKMEN  �;�?�?�0RESTORE 1OC��  �L?��6OCC1O��maO�O�O�O�O�O uO�O__,_>_�Ob_ t_�_�_�_UO�_�_�_ M_o(o:oLo^oo�o �o�o�o�o�oo  $6H�_Ugy�o ������ �2� D�V�h�������� ԏ����w�)�R� d�v�����=���П� �����*�<�N�`�r� �������ޯ�� �&�ɯJ�\�n����� ��G�ȿڿ�����7oSCRE�0?�=u1sc+@Wu2K�3K�4K�U5K�6K�7K�8K��2USER-�2�D�SksMì�3��4��U5��6��7��8����0NDO_CFG� P�;� ��0P�DATE ���None�2���_INFO 1eQC�@��10%� [���Iߊ�m߮��ߣ� ���������>�P�3��t��i���<-�OFFSET T�=�ﲳ$@������ 1�^�U�g��������� ��������$-Z@Qcu���?�
�����UFRAME�  ����*�R�TOL_ABRT8	(�!ENB*?GRP 1UI�1Cz  A�� ~��~�����!���0UJ�~9MSK  M�@�;N%8�%x��/�2VCCM�³V�ͣ#RG�#Y��9���/����D��BH�p71Ce���3711?�C06�$MRf2_�*S��Ҵ�	���~XC56 *�?d�6���1$�5��m�A@3C��.' ��8�?���OOKOx1FOsO�5��51��_O�O��? B����A2 �DWO�O7O_�O8_#_ \_G_�_k_}_�__�_ �_�_�_"o�OFoXo�%TCC�#`mI1�i������� GF�S��2aZ; ��| 2345678901�o�b���� �o��!5a�4Bw�B�`56 311:�o=L�Br5v1�1 ~1�2��}/��o�a� �#�GYk}� p�������ُ� 1�C�U�6�H���5�~� ��ߏ���	���4�dSELEC)M!v1�b3�VIRTS7YNC�� ����%�SIONTMOiU������F���#bU��U��(u FRk:\H�\�A\��� �� MCLOG��   oUD1��EX�����' B@ ����̡m��̡_  OBCL�1��H� �  =�	 1- n?6  -�������[�,S�A�`=�̩͗��ˢ��TRAIN⯞b�a1�l�
0d�$j�T2cZ; (aE2ϖ� i��;�)�_�M�g�q� �ϕϧ��������	���F�STAT 	dm~2@�zߌ�*jq$i߾��_GE�#�eZ;�`0�
�� 02��HOMI�N� fU��U�� ~�����БC��g�X���JMPE�RR 2gZ;
  ��*jl�V�7��� ������������
��@2�@�q�d�v�B�_ߠ�RE� hWޠ$LE�X��iZ;�a1-e���VMPHASE'  5��c&��!�OFF/�F�P2*n�j�0�㜳E1@��0ϒE1!1�?s33�����a k/�kxk䜣!W�m[�䦲�[���p�o3;�  [i{��� �/�O�?/M/ _/q/��/��//�/ '/9/�/=?7?I?s?�/ �?�/�/�?�??Om? O%O3OEO�?�?�O�? �O�O�?�O�O�O__ gO\_�OE_�O�_�O�O /_�_�_�_oQ_Fou_ �_|o�o�_�oo�o�o �o�o;oMo?qof- �oI����� 7�[P����� ����ˏ��!�3�(� :�i�[�ŏg�}�������TD_FILTuEW�n�� �ֲ:���@���+�=� O�a�s��������� ֯�����0�B�T��f�x���SHIFTMENU 1o[�<��%��ֿ���� ڿ����I� �2�� V�hώ��Ϟϰ��������3�
�	LIV�E/SNAP'�?vsfliv��E�����ION �* Ub�h�menu ~߃�����ߣ���p���	����E�.�50�s�P�@j� ��AɠB8z��z��}��x�~�P�� ���KMEb���<�0���MO��q����z�WAITDI/NEND�������OK1�OUT����SD��TIM.����o�G��� #���C���b������RELEASE�������TM�������_ACT[������_DATA 	r��%L����x�RDISb�E��$XVR�s����$ZABC_GR�P 1t�Q�,�#�0�2���ZIP�u'�&�����[MPCF_G' 1v�Q�0�/�� w�ɤ�� 	�Z/  8�5�/�/H/�/l$?��+�/�/�/?�/�/�???r?�?  �D0�?�?�?�?�?�;����x�]hY�LIND֑y�� ��� ,(  *VOgM.�SO�OwO�O�M i?�O�O^ PO1_�OU_<_N_�_�O �_�_�__�_�_x_-o oQo8o�_�o�oY&#s2z� �� �oC�e?a?>N|�o�q����qA�$DS�PHERE 2{6M��_�;o��� !�io|W�i��_��,� �Ï���Ώ@��/� v���e�؏��p�����`�����ZZ�� �N