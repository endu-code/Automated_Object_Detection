��   ʇ�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DCSS_C�PC_T� �$COMMENT� $ENA�BLE 6 MO�DJGRP_NU�MKL\  ?$UFRM\] ?_VTX 6 � �  $Y�Z�1K $Z2�STOP_TYPK�DSBIO�ID�XKENBL_C�ALMD�USE_PREDIC? � &S. �c 8J\TC�~u
SPD_LI_0���SOL�&|Y0  � 1CHG_SIZO$APGESDIS��G�!C����Jp 	�J�� &�"��))$'2_SE��� XPANIN�� �STAT�/ D $F�P_BASE �$_ K�$!� �&_V�.H�#u h$J- ��ZAXS\UPRJLW7Se���&� | 
�/�/�/D&?8?z�h$ELEM/ �T ��2�"NOxG�0�3UTOOiƤ2HAD�� $oDATA"�%e0  @@p:�0� 2 
&PNp% � p!U*.n   �FS�CzH�B� �B(�F�D(��RUC�DROBOT��H�CqBo�E�F$CUR_2Rh$�SETU�	 l|� �P_MGN�INP_ASS� 0"@�� �3�8B7gP�@U�^V�Sp!�h$T1�
`B|8�8�TM �0 6P�+ Ke�1V�RFY�8
dD5F1ȕ ��W��1$�R�8SPH/ ({ �CA�CA�CA�3�BOX/ 8�0������b�'oEjTUIR�0 � ,{ FR`E}R�02 $�`o �a_S�b��gZN/ 0# {9F0� -a0rZ_0�_0�u0  @Q�Yv	�o~:o �$$CLLP  ����q���Q��Q�pVER�SION�x�M@�5�qIRT�UAL��q' 2� �xQ   ��Double� Parts SGide�� �0�p����#PD � DM-�N���  �@k���Ŀ� �����0��q��/�A�S��^���
�y�DJ@� D�p+����� �򫏽�r��a�W�u� ���ٟ�Z��~��� Ɵ��F�{������� � 2�h�����/���S� ¯ԯ毛�
���ѿ@� ��d�v���=Ϭ�a�s� ⿗ς��*���N�� ߄�%�Kߺ��ρ��� �߷�N�8���\�n�#� ��G�Y�k��ߏ���� ��4������|�1��� ��9���w�������� B�T���x�
?Q�� u����,���� b���_�� ��(:L/p %/7/�[/F/���/ /�/�/H/�/?~/�/ E?�/i?{??�/�? ? 2?�?V?OO/O�?SO �?�?�O�?�O�O�O@O �OdOvO�O�O;_a_s_ �O�___N_<_�_o o�_9o�_�_�_�opo �o�o&o�oJo\ono# �oGY�o}�o�o �4��j�
�� �g���������ӏ B�T�	�x�-�?�֏�� u�������ϟ�� b������M���q��� �����(�:���^��� %�7���[�ʯܯ� � ��ǿٿH���l�~����E�4�i�{���$D�CSS_CSC �2!���?Q  D���� ���*ƶ������A� �S�4߉�X߭�|��� �����������<�a� 0�B��f������ ���'���K��o�>� P���t��������� ��5Y(}L^���'ɘ�GRPw 2�� ��,�	Z�?*cN� r������/ )//M/8/q/\/�/�/ �/�/�/�/?�/�/7? "?[?F??j?�?�?�? �?�?�?�?!OOEO0O iOTO�O�O�O|O�O�O �O�O�O/__S_>_w_ �_�_f_�_�_�_�_�_ oo=o(oaoso�oPo �o�o�o�o�o�o�o' K]o:�~� ������5���_GSTAT 2���1�,8��?�  �?����Ǚg�8�(����� ,��Ǫ�4� ���y�Dr*@�m�aDC��$�8�t����z�1�/�/��4���Ux������ĀZC�����/����t��~��8z���?�D���<:z?����̉B��Y��"�DE:�=�����|�@?�|�:z�+�����ު�|�:�z(�=��B���a�נ�D�j���|�<�=��D�̉��A��bD�\�������2��m�:����(C��4���ſ&x���v� ����ȑ������ � F�X�6�|�����͐'� ��%�ęį�د��$� �0�Z�D�V���z��� ����n�����>�P� .�tφϠ�ڿ��� ���������:�<� N�pߚ߄ߦ����� � �d�6�H�&�l�~�\� ̟ޟ������ҏ��� ��,�>�P�b�t��� �����������> ��.t�d���� ������(R <^�r���� ���6/H/&/l/~/ \/�/�/�/�/��/ ?�/ ?J?4?F?�?j? |?�?�?�?�?�?�/.O @O�/dOvOTO�O�O�� ����������&� 8���\�n�t_������ �������O�O"\ono �O~o�o�o�o�o�/�/ O�?"L6X� l������� $���of��oV����� ��ҏ��o8���� D�.�P�z�d������� ���П���ď^� p�N�������ʯܯ�O ,o>o�O_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
o����Ro�Ϟ� �����ϲ���
���� 4�>�0�R�T�f߈߲� �߾���������*� T�F�����Ϧ���� ����.�h�>�D�J� t�^������������� �� "L6�� ��~����J� \�n�,�>�P�b�t��� ������ο��<�� (�:�$6H��/�/ �/�/?�/(?:? �Z d?np?�?�?�?�?�? �?�?�?O$ONO8OZO �Ov�O�O?�O�O�O  _2_L?vO\_�OX_z_ |_�_�_�_�_�_o�_ oFo0oRo|o�O�o�o _�o�o�o*z/ �/�/\n���� ����/"/4/F/ X/^�Tf�/��� ܏"�4��X�j�P_�o ��fo��ʟ��֟ �� �6� �2�l�V�h��� ��J����ԯ�,�
� P�b�|�����ʯ��¿ �����������*� L�v�`ςϬ�ү���� @��$��H�Z�D�� ��z������ 0�
��.�@�R�d�v� �����ߖ�Џj��n� ,�R�0�B��������� ����������0 <fPr���� �z�&J\: ��������� ��(//4/^/H/Z/ �/~/�/�/�/r?? �/B?T?2?x?�?t��� ��߼��������� (�:�L�ROp���� ����?�? �:_L_f? p_�_`_�_�_��/�/ �/�/ o*oo6o`oJo lo�o�o�o�o�o�o �/�_D�_TzXj ���_��o�"� �.�X�B�d���x��� ď��Џ��䏢<�N��,�r���b������q��$DCSS_JP�C 2�u�Q ( D���#�� �@� G��(�}�L�^�p�ů ��ӯ���ܯ1� �U� $�6�x���l�~�ӿ�� ��ƿ��?��c�2� ��Vϫ�zό��ϰ��� ��)���7��q�@ߕ� d߹߈ߚ�������� 7���*��N��r� �����������E� �&�8���\������� ����������@e 4F�j|��� �+�OsB T�x����� �9//]/,/�/P/b/ �/�/�/�/�/�/�/�/ G??k?:?�?^?�?�? �?�?�?O�?�? OUOP$OcO"�ԕSݐ�@NO�OrODO�O�O_ �O?__$_u_H_Z_l_ �_�_�_�_�_�_�_;o o o^o�oVoho�o�o �o�o�o�o7
E .Rd���� ���3���*�{� N�`���Ï������̏ ���A��&�w�J��� n���������ȟڟ� =��"�s�F�X�j��� ����ޯ�֯�9�� ]�0���T�f�����ſ ����ҿ�5���,� }�P�bϳφϘϪ��� �����C��(�y�L� ��p��ߔߦ������ ��?��$�u�H�Z�H�MODEL 2ΟKxp�e�
 �<��c��  g���l���� �R�)�;�M�_�q��� ���������� %7�[m��� ����a�J�� !�	w���� /��B//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?t?K?]?�? EW�?�?O?�?�? LO#O5O�OYOkO�O�O �O�O _�O�O6___ l_C_U_g_�_�_�_�_ �_�_ o�?�?�?oo �_couo�o�o�o�o�o �o�o)vM_ �������*� ��`�7�I�[�1o�� Uo����k�ُ�8�� !�n�E�W�i�{����� �ß՟"�����/� A�S���w���֯���� ѯ��0�ˏ���x�O� a�������俻�Ϳ߿ ,���b�9�KϘ�o� �ϓ��Ϸ�������� L�#�5�G����A�o� ��������$����� 1�C�U��y����� ��������	�V�-�?� ��c�u����������� ������d;M� q������ N%7I[m ���/���/ !/3/	�/-[/m/�/ �/�/?�/�/?X?/? A?�?e?w?�?�?�?�? O�?�?BOO+OxOOO aOsO�O�O�O/�/�/ �O�OP_�O9_K_]_o_ �_�_�_�_o�_�_�_ o#o5o�oYoko�o�o �o�o�o�o�o6 l__GY�A� ����D��-�z� Q�c�u���������Ϗ �.���)�;�M�_� �������}���ϟ <���%�7���[�m��� �����ǯٯ�8�� !�n�E�W���{����� �ÿտ"����X�� ��E�W�-ϛϭ��� ����0���+�=�O� a߮߅ߗ��߻����� ����b�9�K��o� ���i���ϻ���� �#�p�G�Y���}��� ��������$��Z 1CUgy��� ���	��h� 1C������ /�//d/;/M/�/ q/�/�/�/�/�/?�/ ?N?%?7?�?[?m?? U�?y�?�?&O�?O \O3OEOWOiO{O�O�O �O�O_�O�O__/_ A_�_e_w_�_�_�_�_��_�_�_�:�$DC�SS_PSTAT ���_a�Q    �po~j no A(�o�o�o�o�o | �```q�`7o0B�9*c_elpa��~PdSETUP ;	_iB�"d�3��1�tKiT1SC� 2
�zp�1C�z�3��+��uCP� R�|��0D �?v����?����Џ�� ����<�N�`�/� ����e���̟ޟ��� �&���J�\�n�=��� ������گ��>d�!� 3���W�i�{�J����� ÿ������ڿ/�A� �"�wω�XϭϿ��� ��������=�O�a� 0߅ߗ��������f� ��'���K�]�o�>� ������������ #�5��Y�k�}�L��� ������������1 C�߼�y��� ���	�?Q c2��hz�� �//)/�M/_/q/ @/�/�/�/�/�/�/V h%?7?�/[?m??N? �?�?�?�?�?�?O�? 3OEOO&O{O�O\O�O �O�O�O�O__�OA_ S_e_4_�_�_??�_ �_j_oo+o�_Ooao soBo�o�o�o�o�o�o �o�o'9]o� P������� �5�G��_�_}���� ��ŏ׏������� C�U�g�6�����l�~� ӟ埴�	��-���Q� c�u�D���������� �Z�l�)�;�¯_�q� ��R�����˿���� ��7�I��*�ϑ� `ϵ����Ϩ����!� ��E�W�i�8ߍߟ߯���$DCSS_T�CPMAP  �������Q @ z�Jz�z�z���z�Uz�z�z�	�W  z�z�z�Uz�z�z�z�Uz�z�z�zЕz�z�z�z��z�z�z�z��z�z� z�!z�"�z�#z�$z�%z�&�z�'z�(z�)z�*�z�+z�,z�-z�.�z�/z�0z�1z�2�z�3z�4z�5z�6�z�7z�8z�9z�:�z�;z�<z�=z�>�z�?z�@��UIR�O 2����� ���0�B�T� f�x����������������,>Py� �y������ �	-?Qcu �����Z�~ �)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?�?
/�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O��Or?_��UIZNw 2��	 �����L_^_p_u�G_�_ �_�_�_�_�_o�_,o >oPooto�o�ogo�o �o�o�o�o(�oL ^p�E���� � ���6�H�Z�)� ~�����e�Ə؏ꏹ� � �2���V�h�z�I� ����ԟ����
�ٟ�.�@�R�_��UFRwM R����8}ߪ���{���ͯ �(��L�^�9����� o���ʿ��� �ۿ$� 6��G�l�~ϕ��ϴ� S�������� ���D� V�1�zߌ�g߰��ߝ� ����
���.�@��d� v�Ϛ��K������ ����<�N�)�_��� ��q����������� &8\n��� C����"� FX3|�i�� ����/0//T/ f/}t/�/�/�/�/�/ �/??�/>?P?+?t? �?a?�?�?�?�?�?�? O(OOLO^Ou/�/�O �OEO�O�O�O __�O 6_H_#_l_~_Y_�_�_ �_�_�_�_�_ o2oo VohoO�o�o=o�o�o �o�o
�o.@d vQ������ ��*��N�`�wo�� ��5���̏�����ݏ �8�J�%�n���[��� ����ڟ�ǟ�"��� F�X�2�