��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ��5/IRTU�AL-9LOO�R G��DD?8�?�������k,  1 <DwH8G�����D��82 ��-��Z�Z]/o/@�/S/�/�/�-_ �/��/�/;�$MNUR>AP"�� 8���=��?{���<�i��t-����D	?x
 �?tt>2qn�>|l��F���9������0���+?��&������S�R��ǿ����Ѯ���w<S����ʢ�Č��C��-b{5��3��?��;�[��?��7J�j�:>�e:>�@��0���ã�AzD���#��
{5��x?��o;'��7ue��'�&�0���0�<�i8��/�ȭO����^��{5�?}�z�B��>d����O0f>>����@�>��?y�BB��hį%"�=%&C*/ fO��_O�O�O�O�O�O��E��?���A�H
T����������1��<H�)��ʠ Č�� C���%7N_UM  ��>�� "5TOOL/?4 
E3�O�_��O�_�_  ¢�����ZDCF���_�_e?�+����YC�;���_o=e�1#B�1�CG��)o�;o�V���zC���aoso�o �_�o�o�o�o/�l�����33C�@:RW1(fTIVyWV#