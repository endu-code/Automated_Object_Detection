��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S�ETHOST�� NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!�N� D� $PRIMA�R_IG !$ALTERN1�<WAIT_TI�A �� FT�{ @� LOG_8	�CMO>$D?NLD_FI:��SUBDIRCA�P�����8 .� 4� H�AD_DRTYP�H �NGTH��tY�z +LS�&$ROBOT2�PEER2� MA�SK4MRU~O�MGDEV�6�� �RCM+ ;$Z ��QSIZ�X�� �TATUSWMA�ILSERV �$PLAN� <�$LIN<$C�LU���<$TO��P$CC�&FR\�&�JEC�!�%�ENB � ALkARl!B�TP��3�V8 S��$�VAR9M ONx
6��
6APPL
6�PA� 5B 	7PO�R��#_�!�"AL�ERT�&�2URL� }�3ATT�AC��0ERR_oTHRO�3US�9z!�800CH- Y�4�MAXNS_�1;�AMOD�A�I� $B� (�APWD  � L�A �0�NDAT{RYQFDELA_Cx@y'>AERSI��A�'ROtICLK�HMR0�'� XML|+ :3SGFRM�3�T� XOU�3PIgNG_�_COPA1�Fe3�A�'C�25�B_AU�� k 6R,2�COU�!H!UMM�Y1RW2?�RD�M*� $DI}Sc �SMB��	"�BCJ@"CI�2AIP6E�XPS�!�PAR��TCL�
 �<(C�0�SPT9M�E� PWR��Xx�X�Qo l5Ȥ�!�"%�7�ICC"�%� kfR�0le=P� _DLV��Y)No3 <oNb�X_�P~#Z_INsDE
C�`OFF� ~UR�iD��c� �  t ��!�`MON�%sD\�&rHOU�#EWA�,vSq;vSqJvLOC�A� Y$N�0H�_HE���@I�"/ 3 $AR�Pz&�1F�W_�\ �I!F�`;FAp�Dk01#�HO_� oINFO�sEL	%G P K  !�k0WO` $oACCE� LVtZk�2H#ICE�>L�  �$�s# O���k���
���
`�K`SQi�  �5|�I�0ALh�z�'0 V��
���F��������܅�$� 2ċ$b�w��@����� č��!r��Z���4���Ċ!�147.87.?224.20h�S���96����܁܁�3�_{p_  �ċ� bfh.ch̟�1�C�U�g� y���������ӯ^�� _FLTR  ���π �����B���n�nxč2n���rSH�PD 1�ĉ  P!
�robstatison֯՚!k�.�Q�ſ������� �޿?��c�&χ�J� �Ͻπ��Ϥ����)� ��M��"߃�Fߧ�j� �ߎ��߲���%���I� �m�0��T��x�� ������3���W�� {���P���t������� ������Sw: �^�������= a$Zׯ$� _L�A1��x!1.�ğP��1�Q255.�%�S���2 ��E �//*/<&3F/�� l/~/�/�/<&4�/�50�/�/??<&56?��0\?n?�?�?<&6�?�%@�?��?�?
O1�?P���MY� MY���c��� OQ� �VN<�O �O_�O+_=_O_"_s_�_NPd_�_�_�_�_ �_o!o3o�_Woio{oVNLoM��o�l�o�Ao
.@U}�iRConnec�t: irc\t//alertsE ����Pu�����1�C�UуP_R8�d��H�~��� ����Ə؏���� �2�D�V�S$���8�(p����o͟ߟ���QA8��d�A�@�B4��j�h9�Q+�n�@DM_�A+�~�SMB 	X��8%ğVO��߯���_CLNT 2
X� 4C�ɯ0��l �c�B�T���x���Ͽ ������)�;��_��q�Pϕ��MTP_CTRL ��%���ϙdc���ߋ�@�?�*�c߳l��N����@{�Vߵ�Ƥ�������ѓC���USTOM d{���}�@ }��DTCPIPu��{��h�E�TELҮ{��A���H!�Ta�t�çr�oblolr�  ����!KCL����F��!C�RT��������?!CONS&�����n+���