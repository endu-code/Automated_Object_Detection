��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP������8 . 4� H�ADDR�TYP�H NG#TH���z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�� RCM�+ ;$xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAXNS�_�1�AMOiD�AI� $B�� (APWD � � LA �0�N�DATRYQFDE�LA_C@y'>AERcSI�A�'ROtICLK�HMR0�'� �XML+ :3SGF�RM�3T� XOU>�3PING_�_C�OPA1�Fe3�A�'C8�25�B_AU�� 8k 6R,2COU�!H!_UMMY1RW2?��RDM*� �$DIS�̌ S�MB�	"�BC�J@"CI2AI<P6EXPS�!��PAR�te�RC�L�
 <(C<�0�SPTM�E� �PWR��X�VV!S=Mo l5�d�!�"%�7�ICC��%� kfR�0leP� _DLV��U�Q)No3 <oNb�X_�P~#Z_INsDE
C�`OFF� ~UR�iD��c� �  t ��!�`MON�%sD\�&rHOU�#EWA�,vSq;vSqJvLOC�A� Y$N�0H�_HE���@I�"/ 3 $AR�Pz&�1F�W_�\ �I!F�`;FAp�Dk01#�HO_� oINFO�sEL	%G P K  !�k0WO` $oACCE� LVtZk�2H#ICE��L���$�s# �S��k���
��
`��K`SQi�_  �5|�I�0�ALh�z�'0 ��
���F��������܅�$� 2ċ��w������� č��!r�Z����4���Ċ!1�47.87.22O4.20h�S����96����܁܁3�_�{p_  ċ�� bfh.ch ̟�1�C�U�g�y����������ӯx�� _F�LTR  ��π� ���������n�nxč2n��rS�H�PD 1ĉ�  P!
ro�bstation\֯՚!k�.� Q�ſ��������޿ ?��c�&χ�JϫϽ� ���Ϥ����)���M� �"߃�Fߧ�j��ߎ� �߲���%���I��m� 0��T��x����� ���3���W��{��� P���t��������� ����Sw:�^ ������=� a$Zׯ$ _�L�A1��x!C1.�ğP�1�>Q255.%�&S���2��@E �//*/<&3F/��� l/~/�/�/<&4 �/�50�/�/??<&56?��0\?n?�?�?<&6�?�%@�?�?�?�
O1�?P��MY�� MY���c��� Q� �VN<�O�O_ �O+_=_O_"_s_�_NPd_�_�_�_�_�_o�!o3o�_Woio{oVN LoM��o�l�oAo
�.@U}iR�Connect:� irc\t//alertsE�� ��Pu����(1�C�UуP_R8�d��H�~������� Ə؏���� �2�D�DV�S$���8�(p�����o͟ߟ��Q$A8��d�A�B4���j�h9�Q+��@D�M_�A+��SMB 	X�8%ğ�VO��߯���_CL�NT 2
X� 4C�ɯ0��l�c� B�T���x���Ͽ���� ��)�;��_�q�P�����MTP_CT_RL ��%�� �ϙdc���ߋ��?ߐ*�c߳l��N���@�{�Vߵ�Ƥ��������ѓC��US?TOM {��љ}�@ }�DT�CPIPu�{���h�E�TEL��{��A���H!T�a�t�çrob7lolr�  ���?!KCL�����F��!CRT���������!�CONS&����n+���