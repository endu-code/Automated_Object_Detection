��  ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCTD_�DATA_T � �<$SW�_DIR  � BCONST�IFDABS � ^SdIII�gCTCH iS�N��KEI_D�gT1D_f$�NUM��� �MN�COMa ��]AI  �M�
�o �SA (FS�ZZ*TFSOrO*FSU9U*�OPM ��OR�DRM~'$II� �F�� �_SIP���EMJ�SN�"!S&����B"1$�CT�ZU(�X%H=&KP��~$�~"��$�'IR����"1$�^%�#l#�DO#�#�$�M�(0�&2�$0S�F� / B3w<�MENW ��MCMF_C�/1T4EN�U3T�W�U3FDB]8C�j9FGgTOOL_� �~4IU4I�0�_FR�1�1TR�QGAI� O$TDC�1� J�$>�2$DSR�2AWEV "G A�A�L_TI�1$MOVE_L�#�WG��TRN@Y�,A 44PAR��   ��T0PEEa �6�BKB�JD,E�D �CK�KK�ID_M�I�@�K@�J3�J�J1P�IFP�Sk" 44SU��0  L�$LIMIT�2� $INSER�TE@$�@A
E{NUyRSRBP�Y�P�W41I3�bH;NX0~P��RBC@�WTE��Th6f�QALx4bAE�WFV�3c�c�2|QZGbU�XUN%hV�P�T\4neUwhGRA�Px!�TRETRY�f�g1�l2gEC�_DDE#�a�gA�_POf �bANP�0�eFT]DL#KALRCT%`�3V/2,-p�VCvb=p�bK$�bA�<pL�}Pl#HD_RAPXfuD�yq�kq�w�UR$p�B��tVA_SWMb�p�3�q��p5E�A�PLE��smM�OR]CPH$�FSDF]@�2F_LpR�4CP�� P%a�W@TN_Vi CuNM@F�MIN�p��Eq_ML_LM>�VEL_CU �s�$AUT_RV�h�t�qp� 
CEPT�H�a���a^�X�DA�MP_�3UA��Y0O�RCSTOP_TH3REfȄAV��h0����t�RA%q�M��� І�AZ@��OSC_GD� �s0��)��$FORCE_O�@{PMOL1b�!�HOP�4R�U�P�T���ROT�PCx!�PC�RED{P����CH1G`��tєDP�ғ�V�����R�a3qINISH�3��1OF�_��t��d��u��F�χ`�OCITY(p�`��NsPD�`�t0���$���A �ScTk_}_�_�_�W�05� ($WO�R�A 2$�\A ' /�C2[R���ST̀ ���CH�r�_�#RVd�Ln�N�E_��F�_�AC��_�C`]q�2}��ck�_M���DC�$_�V�3k�V�����W������d�8��d���RTN��i��T�A����ALGwO_S~�$P�a���x�REV_I�T!��MU�t�`C!COF�Q>���X���wGAM�PAS��v��_O�NTR��YFѐ��TR�V�CNPL��E���*�rtCNC`+1"�ѐ-O�CHW�L�_��F-�r�;�d�OVMb/�QR�!֢�IO���D���hע�JTH�l#d�PA�����P�DA  i��DSP�VsCNMONLS@��*�w$8�RC��V��P�KPGRI�j�R�Gfu�˔x��u�O���g�T��O�Ae�R�vb����V�13��PyD���AGWA֗��THӃ%��q3�M0��E����VRYac�� �g�M��g���OVK���� /յ�;֌���VL^�!���T1CO���_�TR�/1u�MG�sI�o��.xy@%a8INDEsq�ϐTM9�זZCC���ZRGCUSP�F>����qp��T�WD�Ʊɖ�SR���7t���OL�&�?��q<NSK�܀P`��sAXCP�_P�r+R�(SR��-DI7�-E��$�J,E�RTY�L�UFFIXE�sR�EG�1�����F���Ѐ1sM���CgNFC��EN�0��V��E�RT�V*TMU�RG` �4 Z��4 DU?B-'TS Y(**�@Ss��z%PQz$|z%IP�/�4 AP���(�!V�]C2"N,�0PM`���!�н�#RC�(P!8'�@QPY0H5&@B4��_sC3���r.[R�_p�d`U��@VAD>CMVROU
b�1�PERIO�sF1P���2D-��3%T��1_D��2�Ĥ�3��T����K�9K��K�7CL���0�gADJ����_Udr;[PAUX�@�_	 4�@C�P?a$� A�&�n@ ~qUX_AXS��PJF�� 
 h�D�rӠ�Cd� �C�t�C�F�@�H�G1P��FOXp4XAXISU� Tj��D͡ȹq�E��AP@M@ �	BQ܀HR
$I�DX\PRV�QSa�GR�T�L $FN�E_Uנ���TTOOL�R�p;�A���p�y1DOf` �\��0R_PKG��RQ BQ �NR�PBQS�P[Q 2	hQ�P��S�P2�Q�Qdba	�1a~d�$VFLw03IM�,�LT�r��:a��Tc�6Tb����O$DYG��C$d0
JgGUg	�d�4�d�c�MPSWP  �$� @��  ��i��a�@&�@ &�`VERSION�h�  ��5�aIRTUAL��o�avS?�h&?�  �aL| J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x���a+u|P11 2�9{\�@p��� ֓Ә�� � ?�a @x�@����A�  � ����#����3��-��?�Q�?�g�U�����  D  Bp�  =��Ϳ�?333?�a�̠��̤@��ߥA ��/�  & G�P �?fffˡ>��ߥ�������0�ܙ D���̤ˡ��k�C� Z�[��`�0�����ӿٲ��B�ђI@ɟK��ÿ��;���F@� K���������Dz ��l�W�I��ٺ��ܑ�P`��w���ēV��'�9�K�]�o�5� ����_�q�ۿ���� ���#�9�G�y�7�I� j�߳�����������a��!���y�3�� ��ϋ�9�K�]�oρ� �ϙ���x���D���� �������,>� b������� ����ɤ����ȗ�Đؓ��� �2/d���L����^/\�Ϣ�]�ĐW��"�@
�"��'B��������8�/"  $đƚ�$1>B,4_��(�ā��1?��?�?�8>����ā�//@/ �?T/f/?O�/�/�/�/ �/�/�O??,?>?P? b?;_�?__�?�?�?�? �?OO(O�_o^OpO �O�O�O�O�O�O�O _ _$_�oH_Z_3~_�W@��fx���2�� ���	���o2�2-�V�h�z������� ԏ��������Dq dd�����l��ߩߩ�b �����o����ğ���cd�p(������qT�@� a>Ho�
}p��[��c|�>LŠ��_v���<#�
�Qsbp|��X��o�C��� a?e?a��3�T`��@ �G_� 
�T���_����x�2bo%{Bta�������@1��U�g�k�`>X��ؤ����ϑ�It$� ��$$�>�٢
���A��߭�'��ϼ��4�+���s�.����Ճa$�=���(4$ܛ�S��e�;��.��>���H�Ճa5�����8M�Y��;�=@���3��a�B�	9� R�=�v�a�ߡ����������m����  �b\'��� ���`k�S�K�X�,�w��������/�����C���Q�??333�;�s�<��saD/ � C``G�P ?fff/a>$���? _	W�_��0��_g� ;�5c?�4'e���u�j� F�@ ��[�� DzI ���w5����y ܃�� ���/���/�/7 I�_I/[/m//�/�/ �/�?�?�?�/?!?3? E?W?i?{?�?kO}O�?�?�L�Oq�O�� �����O���O�O �_
__._@_R_d_o �_�_,o�_o�_�_o obo%`&/ $.(��?��>�"� �o����}��o��E+ ̰�B��+��ȴC�� 8�����{j4�~gĠ{t ��"�������$�3t�7�q�����>���3t�cu�� ��������)� W���_�q��������� ��ݏ�ȯ�%�7�I� k�%����j���ǟٟ ���Ϳ3�E�W�i� {�a�������կ�L�o 0��������2Q/ߐA�S�e�v�Uώ�2 �߲����������� 0�B�T�[Ru���� �����7M;	;	/�DO *GT�V� �M�D�i���Op�����Ѱ�
���A>�a��f��28�BH���>L! xH���g�<#�
�ϲp��w�E�v������A��7������@\A�b�f� �D?B,��7J���_���Bб���Z{� p��N���>�4�_�U�/��It$ Z//$��>�5
/a'A��a/	/�/-/?&ސ�+����%.�����%��$敕�%(4$��%�/�+�;��.#5>��yH/5��5��?5O8M�YK5��=  g5��8�x?�+	�/�? �?�?�7?�?O$O6O�HOZO�o�GnlG  ;¸`�X ���E�E��A��O�O@�O	_�2 _^����`y=�e?333����B�����D/  �C��G�P ?fff��>���e�Y �Q�iȌOVb�m��� �W�i�]ooo�o��k���_wo�o�`F@� uawU�`Dz �P$to�o�jn���� ��_�_oo 'o�KoU�)��o�o ﯥ�����1� ��"�Y�k�}����� ��ŏ׏�ǟٟX�1��̸k��oC��o '9KQ���0�B��� f�x���������z�� �����l�>�P�b�t� ��lu�ς\�nπϊx�O�������4� ����C�<���R( ����c�$�C�  ���׺��ڷ  �Ę��~Jk���_V�؏���/�?�Q�]�>�����]��������� �+��O�a�s߅߳� U������������� 9�K�$o������ �������#�5�G� u�k�)���������� ����1ǼZό�/0/B/X%2�l�/�/H�/�/�-��"2�/ ? ?2?D?V?h?z?�? �?�?�d�n�>�GY GZ<���Y�Y����� ��ijO|O�O�O�FK �GLO^Ib!W�#�> �'_����4U>L}PdQ�<.B�<#�
K+�p4_�B�t�FB�����SU�RkU@��lT��o�δ ���ζ��0o��eB,TUPo�o�o�o�o��P>a�T�Ox�OrICIt$ �-$�&>��R
k�wAHD�e���v�@�+���+�.��y�7��A$敕G��(4$�S���;���.�>��H����A5����8'M�Y���==dPÅ�B�ԏ�{	�
��� .��g�Y�n�������ඟ%o�=��ȗ  B��R�T_b�P #��J��X/�A�S��e��|�j�B�	�<�S��?333�E+���D7IcaD/  C�G�P ?fff�A>�Q8D���� O=X蟲��M�O� ��o��˿���?Y��ӿ-�Kl�F@ `_�k�ӥbl�Dz� ��k�]�/��~!^/P) �;�M�_�q��� Iߧ���s߅���K ��%�7�M�[ߍ�K� ]�~����������� !�3�u�#�5����Sl���)ϟ�M�_�qσ� �ϧϭ�GR����X�� ������
�@R �v��������/�ϸ����ȫ�� viڗ�N. k_=C��/o�㢄`s� ��U�"�d�Q�f�PcE ci3�/6|P3$�ښ@�$E>�Us��(���)o�<�?�8>��� ��:/-/?/Q/c/u/ �/`O�/�/�/�/?�O ?)?;?M?_?q?J_�? �?�_�?�?�?O#O�_ 7OIO"omOO�O�O�O �O�o�O�O_!_3_o W_i_B�_{���z���u2	����$�.�F�2A�j� |�������ď֏��� ��
�-�Xqxd���� �l�����b������Ɵ؟���!�wd��p<������qh�T�_a>\��}z�o� s��>L٠�� o���y<#�
�Q�bp���/�l��o.�c���_aSeWa��G�h`ǥ@�Ȥ[s��T���_�V�ꌿFbo9{B �a�����3�E�(�i�{�.k�>l������ϥ�It$ ��$�8�>��
���A������;�����H�+���̇�.������G�$敕��(�4$ܯ�g�y�;�{�.��>��H���G�5����8M�Y�O�=���G��a0�V�	M�f�Q�� u��ߵ������� �����'��$�  �bp;������ g�_�l�@���������PC�����c��e��S?333O���P�|��ñD/  Ct`�G�P ?fffO�>8���Ss	k�_ !xD�s{�O�Iw S�'H;e#��/x��j� F@ �0�/o�� Dz] �����I�q��y ܗ�����/ /�/�/K]�_]/ o/�/�/�/�/�/�?�? �??#?5?G?Y?k?}?��?�?O�OO�?g|� #O��O����� /	_���O�O�__0_ B_T_f_x_2o�_�_@o �_$o�_oo,ovo$%�t:/&8B(� OPp\cҹ6��o�~ǯ ���o��E?��BPp ?��ܴW���L����� �jH��gؠ�tPq6�#� �����8�GtK߅�x��	��>���Gt �w������ ����+�=�k��s� ��������͏���� ܯ'�9�K�]��9��� ��~�ɟ۟���-�#� �G�Y�k�}���u��� ů���lD�������2eC�U�g�y���iϢ�2������ ����� �2�D�V�h� of���Դ������ KMO	O	C�XO>Gh�j@"�4�a�X�}�Ӵ�@���������p�>�a��z��B�B\���>L5 \���{�O<#�
��p������E,ϊ������p������İ#@ pA$�b�z�B�SB@�@KJ���s���B� n�������t >�Hs�i�*/^�It$ C/$��K>�I
#/u'A ��u//�/A/S&��+�{���%.����%ޣ�$敕�%(4�$�5�/�+;��=.75>��HC5���5��S58M�	Y_5��= {5��L��?�+	�/�?�?�?�7 ?O&O8OJO\OnO}K��$CCSCH_�GRP12 2�����A?&� \��Xo>��  O��` �lt �E�E���A �__,_>_�2U_C^ʿ���`Q�e?3�33��R����#D�/  CаG�P_ ?fff��>� ��e�Y�Q�}��Ojb �m����W�i��o�o �o���2o�o�E`F@ 8uDa�U�E`Dz�PYtDo6p�j6��� �o &o8oJo\o"��o�L� ^��o�o����� &�4�f�$�6�W����� ��ď֏����N������f����x� &8J\n����� e�w�1�������ѯ� �����+���O���s� �������u�Ϸ���ϵϿxȄ���ٳ .��i�'�#��x�q� H��R<L������8 �W� ����� 4 ����J���sLV�����/�t���>����Ē���� �*�<�N�`�9��ߖ� �ߺ��ߊ�����&� 8�J�#n��Y��� �������"��F� X�j�|�����^���� �����0B/f������S/e/w/�%2@�l�/�/�/�/=�22?C?U?g?y?�? �?�?�?�?�?�d�nN 1!Q|Y|Zqȝ�Y�Y �՟����i�O�O�O�O�FP� W�O�I(�!AW-3�>5�\_��S�H��iU>L�P�Q�cB�<#�	
�`pi_RE��V<B���,0�U bA�U@푡T4� Lo��В�fȚeo��Ba�U�o�o�BT�P>�Ea�T�O�O�~CItk$ �$6>��R	
��wA}D���x��v!P+���`��.���l� Q$�{��|�(4$܈��@�R�;��.��>���H�� Q5�=�Ѕ8M�Y܅(M�=�P�� R�	�/�	 &�?�*�c�N������� ��ǟٟ�Zo Mؾ��  �I�b �T�b�PX�@�8JE�h d�v����������<B��>��S,�?33�3(U`�)TlI�aD/�  CMG�P /?fff(Q>amD ,�L�D�����L� TM(_"�P�,� �!π�?���bπ��F@ �Š��Hb��Dz6��Ġ���d�"�8�!�/�) �p��� ������~�ܿ�Ϩߺ� $�6π6�H�Z�l߂� ���߀��������  �2�D�V�h��X�j���������^����� �Ϧϸ�������|R�� �����	-?Q u����� �O��M/���/����) 5�i ���.�_nC��/�� ��`��) e�"�d0a �f%`�E�ih!?k�P h$)!��$z>�U��8� $$�^o�<�?�8>��� $�:P/b/t/ �/�/�/�/�O�/�/? ?D?�OL?^?p?�?�? �?_�?�?�_ OO$O 6OXOolO~OWo�O�O �O�O_�O�o _2_D_ V_h_No�_�_w�_l@�/����u2>� �.�@�R�c�B{�2v�����ÏՏ��� ��/�A�H�?�b��q �dةت�l$�(�(�r 1��AC����:�1�V��d�pq�ݟ��q����Ia>���S}p���5sť>L����5o��Ty<#�
�Q�bpůd���c�����Ia�e�a�|��`��@I������ Sd,�o۶$���{bLon{B�a��G�h�@z�]Ϟϰ�ckM�>���!�L�B��ړIt$� �$m�>�"�
��N�AٔN���p�߼,�}�+��̼�.������|�$�=���(4$��՜�ޮ�;��.�>���H�|�5���,�8M�Y8儝=@��T�|�%qe��	�� �������������#�5�G���\�4Y�  (r�p�E� �M���������u����������x�������*��?333�����ș��D/ � C�`G�P ?fff��>m�ɔ� �	��_Vxy�C��� ��~���J\}pe�X��d��j� F�@ ��d��� Dz� $���~���y ���� �/8B/??� ��_�/�/�/�/�/�/ ?�?�?OF?X?j?|? �?�?�?�?O�O�OEOO�L�XO�0_�� //&/8/>_آ_/_ �_S_e_w_�_�_�_go �_�_uooYo+o=oOo ao�oY%�o/I[mw(�<O�p�c�k� !�~��Γ0)� Ut �R�pt�P�Č�0� �������j}��g��t �qk�X�֎L�m�|t��ߺ�,�>�J�>���|tJ����� ����<�N�`�r� ��B�����̏ޏ��� ۯ&�8��\�n����� ��n�ȟڟ�����"� 4�b�X��|������� į��������p�G y��/�E�2�xߐ�ߜ߮߿�����2 ������1�C�U�g� y��������	� 4	4
)̀M�	�	xO sG�ϟW�i��������8���9�K�O���
�� Q>�a��R8 R��!>Lj Qx����<#�
8��p!���EaϿ����� Q��@���X@�AY�b�� w��Bu�7�Jײ����B�A=��� ��/��� >�}����_/6�It$ Zx/$��>�~
X/�'A5��/R/�/v/�&���+���5.����$5��$敕45(4$�@5�/
;�;��.l5>��yHx5��5���5O8M�Y�5��=Q  �5����?�+	�/�? �?OGT?FO[OmOO��O�O��n�G  ��p��L � U�E���A�_._@@_R_�2i_W^����`y��e?333���R��$�XD/  �C�G�P ?fff��>�-��ei �Q<����O�b}��� �Wy��o�o�o̵���Fo�o8�Y`F@� LuXa�U Y`Dz �PmtXoJ�jk�K�=� �(o:oLo^o po6��o�`�r��o�o 8�� ��$�:�H�z� 8�J�k�����Ə؏� ��� �b��"���z�4������:L^ p����4y���E� ����ӯ���	�ÿ-� ?�ѿc����������� ϵu���Ϸ����xȘ����c�G}� ;�X&�υ�\��Rq `������m���  P�P ���#�i  �����J��2�`V������/����>����Ħ���,�>�P� b�t�M��ߪ߼����� ����(�:�L�^�7 ���m��������� �$�6�Z�l�~��� ����r������  DV//z�����g/y/�/�%2�l�/�/H�/
?=�322.? W?i?{?�?�?�?�?�? �?�? t�nNE!e�Y �Z�ܝ�Y�Y��ϗ ��i�O�O�O�OVd� )W�O�I�!UWA3L>I�p_-g�\��}U>L�P�Q�<wB)<#�
�t�p}_RY��VPB��L@D�U4bU�U@��TH�`o/� ���fܚyo3&+Bu�U�o�o 2Vh`>Ya�T_x�O��CIt$ �-$%6>��R
��A�D��(���v5P�+���t�.��y���4Q$敕���(4$ܜ�T�f�;���.ȅ>��H�ԅ4Q5���8'M�Y��<M=�P�4R��C�	:�S�>� w�b�������ɟ۟����noM��  �]�(b�T�b` l�T�LJY�-hx��������0�ů��PB�R�<�S@�?333<Ut��=T�I�aD/  C�aG�P ?fff<Q>%a�D@�`�X� �(1���`�hM<_6� d�@��5�(O����vϔ��F@ `�Ŵ��\b��DzJ� �Ĵ���x�6��!�/�) ܄�������̿ ����ϼ���8�Jϔ J�\�n߀ߖߤ��ߔ� �������"�4�F�X� j�|��l�~��������r����ϨϺ��� �������R����� /ASe�� -���c��a/'�//%//����= I�i#���. �_~C��/��,��`�� = ,e2�dDa�f9`�E �i|5?�P|$=!#�@4�>e��%84$8��ro�<�?H>��� 4$Jd/v/�/�/�/�/ �/�O�/??*?X?�O `?r?�?�?�?�?�_�? �?�_O&O8OJOlO&o �O�Oko�O�O�O�O_ _�o4_F_X_j_|_bo �_�_��_(l�1/����u2R�0�B�T�$f�w�V��2���� ŏ׏�����1�C� U�\�S�v��q�d�� �l8�<�<�0rE�+�U�W��!�N�E�j��d��p���������]a>�̯g}���Is٥>L"�	�IoӒ�hy<#�
�Q�bp�ٯx���w�����]a�e�a�����`�@]�����g/d@�-o�8�տ�b`o�{B �a����[�|ώ�qϲ���wka�>��5�`�V����It$ 0�$���>�6�
�b�A��b�
߄�.�@֑�+������.�����Ր�$敕��(�4$��հ���;�{�.$�>��H0�ސ�5��@�8M�YL嘝=	�h吢9qy��	�߯���� ������%�7�I�[��j��$CCSCH�_GRP13 2������&� \�~|E�y  <r ���Y��a������� ����+��B�0����>��?333����ܙ��D/  C�`GÿP ?fff��> ��ᔜ�	��_jx�� W�ĝ������ ���el����j2F@ %%1���2Dz� F$1#/���#���y � %7I?mw/ 9?K?���_�/�/�/ �/?!?S?O#ODO{? �?�?�?�?�?�?�?;O �O�OzOSO\��O� e_/%/7/I/[/m/s_ �R_d_o�_�_�_�_ �_�_�ooo�o<o�o `oro�o�o�o�%��/0~���(�qO�p �cɠ�V��ޓe ^�5U�)�9R�p���� %Ġ�Dƕ����j�� �g!��t�q�����`�9���t��οa�s��>����t�� ���)�;�M�&�q� ������Տw�ݏ�� �%�7��[�m�F��� ����ǟ韣����� 3�E�W�i�����Kϱ� ïկ���߿�/�� S���|�@�R�d�zՁ2��߿����������2�0�B�T�f� x���������� ���>�i	i
^̵M�	 �	���O�G�������������=�m�n�P����.�ڱ>"q�I��@R5R��V>�L� �ƿP���<#�
m�M�pV��2U8����)���ڱ� �u.��@�A� !r9�Ϭ��B��l�JR�ݿ��BN�vr ��/�//A/��� �>2������/k�I�t$ �/$��>��
�/�'Aj��/�/�?�/�& +��̞M5.���Y5$�敕i5(4$�xu5-??;;��.�5�>��H�55{���58M�Y�5�=� �5���?;	?,OOPO;G�?{O �O�O�O�O�OG���n>�G  ��6p ��� EU-U%�2Q Q_c_u_�_	B�_�^�)��+p�u?3�33MRY��D�/  C:�G�P_ ?fff>� Z�u9i1aq���
_�b 9}A�g=y/�o�o ���{o�oOmʎ`F@ �u�a�U5�`Dz#`�t�oQpz�р�r� �]o oo�o�o�ok��o��� ��#m�#�5�G�Y� o�}���m����׏� ����1�C�U���E�W�֟��i���K�� o�����ϯi ����z������,� >���b�t�Ϙ�꿼� ο��<��u:� ���������͟�"� ��G��pލW��Ϻ� ��b�����Ң ����U��X� � U���J��g���V���?K������>������=�O� a�s߅ߗߩ߂����� ���1���9�K�]�o� ���l�������� �#�E��Y�k�D�� ����������� 1CU;y�d/����
ߜ/�/�/�%2@+|	??-???P=//h22c?�?�?�?�?�? �?�?
OO.O5t,~ON z!��Y�Z��ii 	"��./0y�O�O'__CV�� ^W�O�I(�!�Wv3��>~��_�@-����"#�U>L��P�Q"�BA)<#�	
��p�_QR���PV�B����uy�Uib��U@6��T}� �o@/��f��oh9[+B��U�o4�UgJ��P:`>��ad9_/_��CItk$ 	�$Z6>�b	
�;�A�D;��]�x��jP+��̩��.�����iQ$�{��Ņ(4$�х�����;��.��>���H	�iQ5�=��8M�Y%�qM�=�PA�iR!R�x�	 o���s������ן� ���"�4��oIM!�F�  "��]b 2d�b:`�����J��bh ����ѯ�e���讅B����cu�?33�3qU��rT�I�aD/�  C�G�P /?fffqQ>Za�D uŕ����C(f�0� �Mq_k���u7�I�jπ]EO׿Qϫ���F@ ���Q��b�Dz�����ϭ�k�8�!�/�) ܹ�˿ ݿ����%�/���� m���ߑߣߵ��� ���������3�E�W� i�{���������2�����E����� ������%�+�R
 �@Rdv�� T��b�F* <N�FՖ/\�6/H/Z/d��)�r ~�i X�/�.�_�C/?�� a�p��r ae=2�dya vn`�E�i�j?��P �$r!X�E4�>9e�Z8�i$m��oL+O7H>���i$7J�/�/�/ �/�/�/?�O)?;?M? _?�?/_�?�?�?�?�? �?�_O%O�_IO[OmO O�O[o�O�O�o�O�O _!_O_E_i_{_�_ �_�_�o�_�_�o]l@4/f/�
��2�2�� e�w��������Ă2�������0�B� T�f�x����ĈΫ��q �d!�!�|m�q�q�er z�`����D�V���z����d%���&�8�<��҃��>���}p����~s�>LW��>�~o��y<#�
%arp�����N��������e�a-�Ų�`E�@��F��� �ddu�bo$�m�
��b�o�{Bq.�*ϐϱ�@�Ϧ����Ϭk��>��j�����L�#�It$� e�$��>�k�
Eߗ�A"���?߹�c߼u�Ơ+����.�����š$�=�!�(4$�-������;��.Y�>���He�š5���u�8M�Y��͝=@>���Ţnq����	�� �������A�3�H�Z��l�~�������}��  qr����� 9�����ݚ��	�-?��VD����s��?333�ͥΤ�E�D/ � C�`G�P ?fff͡>���� �	�)o�x������ ͯ���ϓ���e���3�/%zFF�@ 9%E��FDz� Z$E7/	/�X�8�*� �'9 K]#?��/M?_?� �%o�/�/�/?'?5? g?%O7OXO�?�?�?�? �?�?�?OOO�O_�OgO!\��O/y_'/9/ K/]/o/�/�_!�f_x_ 2o�_�_�_�_�_�_�o o,o�oPo�oto�o�o �o�o�%��/����(ȅO�p�cPɴ� j(�E��yr�IU� ^�MR�p����Z�ձy� ʰ=�=�zƏwV�� �q�������M���t����u�����>����t�����+� =�O�a�:��������� 鏋����'�9�K� $�o���Z�����ɟ۟ �����#���G�Y�k� }�����_�ůׯ��� ��1�C��g���� �T�f�xߎ�2��ߐ��������� �2 �D�V�h�z���� ���������2�R� }	}
r��M�	�	���O �G�������������Q���������B
.�9�>6q]��TR8IR��j>L� �xڿd���<#�
��a�pj	FU��=���9�-�1��!B��@�A�5rM�� ���B����Jf ���Bb����// /C/U/�� >F�������/�It$ Z�/$�>��
�/�'A~��/�/?�/�&�" +���a5.����m5!$敕}5(4$܉5A?S;�;��.�5>��yH�5!5���5O8M�Y�5)�=�  �5!��
O0;	'?@O +OdOOG�?�O�O�O�O��O�O[��n�G  ��Jp�� � YUAU9�FQe_w_@�_�_B�_�^=��?py�-u?333)�aR*m��D/  �CN�G�P ?fff)>n�-uMi Ea����_�bM}U�) #gQy-/�o"�����o	c�ʢ`F@� �u�a	eI�`Dz 7`�t�o�e#z�є��� �qo�o�o�o �o��o�����%7 ��7�I�[�m�����Ï ����������!�3� E�W�i���Y�k��ß}����_կ��� ����}¯ԯ�� ��
��.�@�R��v� ��Ϭ���п���� P��uN���� �����*�6ìW�� �ޡk����ߥ�b� ��*��Ҷ1�& ���i�"�lǲ i�*рZ��{���V�!��%?_������>���!���Q�c�u߇ߙ� �߽ߖ�������E� ��M�_�q���� ������%�7�Y� m��X�������� ���!3EWi O��x/�����/�/�/�%2?|?/?HA?S?d=C/|22w? �?�?�?�?�?�?OO 0OBOIt@~cN�!��Y �Z�%�)i)i"2�� B/Dy�O_;_2_WV�� rW�O�I�!�W�3J>���_T-����6#�U>L`�Q6<�BU)<#�
���p�_eR��/dV�B��J���U}b��U@J��T�©oT/ -��f%��o|Mo+B��U�oHi{^��dN`>�a"dM_xC_��CIt$ �-$n6>�#b
�O�A�DO��q��-�~P�+��̽�.��y�Ʌ}Q$敕م�(4$�兝���;���.�>��H��}Q5��-�8'M�Y9��M=�PU�}R&!f���	������ ������� ��$�6��H�W��$CCSC�H_GRP14 �2���y��&� \�m.2�p)   )"��qbFd�bN`֥�� �Jávh�����y�(/���B���+c��?333�Uޢ�T�I��aD/  C�G�P ?fff�Q>na�D��ʹ±�W( ��D©ͱM�_���ɉ l�~ϟ�qYOφ���<��F@ �����b�Dz��3�����Ϡ�1�/�) �� ��$�6���Z� d�&�8�ϴ������ ���� ��@����1� h�z����������@(�����g�@����z� ��R ��$�6�H�Z� `�R?Qu�� ������) {M_q��{ժ/`��k/}/�/���^� � �y��C/>�_�C R/K?"��p&� ue r2t�a1v�`�E�i� �?�`�$�!��z4�>Me&��8�$���oNL<`OlH>����$lJ �/�/�/??(?:?_ ^?p?�?�?�?d_�?�? �? OO$O�_HOZO3o ~O�O�O�O�O�o�O�O �o _2_D_V_�_z_8 �_�_�_�_�_�o
oo �@o�li/�/-�?�Q�g�2�̚�����Џ�	���2��/�A� S�e�w����������� �����+tV�V�K|�� �����r�������y� ������Ԧ*tZ�易[�m�q����a>�!6��}-"�sC��>L��s��o=��y<'#�
Za:rpC��p������a@u
qb���pz�@�� {�"&���d��oY� ��?��b�o�{B;qc� _����������.��k˰>���ʯ����X��It$ ��$�>%���
z���AW����t��ߘߪ���+��=�:�.���F����$敕V�(4$��b��,�;��.���>��H����5�����8M�Y���=s������q��	�	 ���=�(�v� h�}���������4�ڝ|���  �r # �ôn�˰2� �>Pbt���y�� ��%?333�:�F�z��D/  C'pGÿP ?fff�> �G�%&^o�x�� �&-.���*)�� ���e֟h�</Zz{F@ n%z�"�{Dz�$zl/�>/���m�_� � J\n��X?��/ �?�?�/Zo?"?4? F?\?j?�?ZOlO�O�? �?�?�?OO0OBO�O 2_D_�O�OV\��O8/ �_\/n/�/�/�/�/�_ V��_�_go�_�_�_o o+o�oOoao�o�o�o �o�o�o�o)�%'��/0����(ȺO� s�����]�z�H�� ��~U����R��΂ ��
�����r�r�Bz�� Ew��B����քT�ʵ���t��8Ϫ���Ș>����tȚ*� <�N�`�r�����o��� ̏ޏ�����&�8�J� \�n���Y�������ڟ ����2��F�X�1� |��������֯���� ��0�B�(�f�x�Q� ������ߛ߭��Ձ2,����,�=��U�2P�y���� ��������	��"$. <�gчĲ	�
���M ��_�G�)����0����K��P����wc�#�>kq��-݉R~Rӟ>�L� �ϙ�.�<#�
����p�>{U8��=r���#�b� f��Vw��@#Q� jr�-���R��J�U�&�H�B���� !/B/T/7/x/�/=�'�>{�&�/��I�t$ �/$G�>��
�/(7A��(?�/�J?�/6W +��̞�5.����5V$�敕�5(4$�x�5v?�;;��.�5�>��H�5V5{��E8M�YE^�=� .EV��?Oe;	\?uO`O�O�G�?�O �O�O�O_!_�6�~>3W  �p J�'�UvUn�{Q O�_�_�_�_RB�_�^�r��tpbu?3�33^�R_���D�/  C��G�P_ ?fff^>G ��bu�iza��0�S_r �}��^Xg�yb/$6 WJ�2��o>����`F@ �u�a>e~�`Dzl`�t�o��pXz���߻� ܦo �o�o�o�o���ޏ ��Zl��l�~����� ��Ə����ȟ� �2� D�V�h�z�����������������2��
� ���� ���� ��	�ÿ-�?�Q�c�u� ��Aϫ���O��3�� �)�;υ�3���I�#�5�G�Q���_�k� �EW�Ϲ����
�� ڥNb�ޢ_�N*�� f
&[�����W�� � ��_�EZ2��&�VG�V�Z?���$�>���V�$��ߘ� �߼����������(� :�L�z������ ���� ���6�H� Z�l���H������� ����<2�Vh z������/��J!�S��/�/	?52@t|R?d?v?�?�=x/�22�?�?�?�?OO /OAOSOeOwO~tu~�N �!�ij,Z�^i^i R"g�M�w/yy1_C_p_g_�V�0�W_%Y()1�W�3>���_��-�ڢk#�U>L�D`+ak�B�)<#�	
�p�_�Rץ;/�V�B����e�b�2e@�3d�� �o�/Qb�OvZ��o���+B�e}��������`>��aWd�_x_9�SItk$ R�$�6>�Xb	
2���AT��,���xP�b��P+�����.������Q$�{���(4$���ҏ�;��.F�>���HR��Q5�=�b�8M�Yn��M�=+`���R[!����	 ��џ������.� �5� G�Y�k�}��o�MjΏ�  ^"���b {d&r�`�ҥ�Jס�h ����,���C�1��B����`c��?33�3�U�T�I2qD/�  C�G�P /?fff�Q>�a�D ��޹ֱ�(��y��� �M�_���ɾ�ϒϳπ��O Ϛ���*3�F@ &�2����b3�DzȰG�2�$��ϴ�8E1%?9 ��� &�8�J��n�x�:�L� ������������� "�T��$�E�|��� ����������<�����{�T������f� &�8�J�\�n�tbS e������ ��=�as ������/��/�/�/���r�� �=y ��W/>2o�Cf/_?6 ��Kp:� �e�2Gt�a fv�`*U*y��?�C` �$�!���4N�e:��8��$���obLtO�H>����$�J�/�/? ?*?<?N?'_r?�?�? �?�?x_�?�?OO&O 8Oo\OnOGo�O�O�O �O�O�o�O_�o4_F_ X_j_�_�_L�_�_�_ �_�_�oo0o	�To�l@}/�/A�S�e�{�2�� ����ҏ�����2�1�C�U�g�y��� ������ӟ������� ?tj�j�_|�������r ������ɍ���̯ï�>tn��o�����/���a>#!J��}pA6�sW�>L������oQ��y<#�
naNrpW���3���*����auqv��/p��@��"":� ��d��omƶ�S�r�o �BOqw�s�����@���0�B��k߰>3�೴ޯԯ��l�It$� ��$��>���
����Ak��߈��߼���+���N�.����Z��$�=�j�(4$�v�.��@�;��.��>���H���5�����8M�Y���=@������q���	� -��Q�<���|������������H�����  �r7 �״ ��߰F.&�3�R�dv�
��*���, ��%?333��N�Z���D/ � C;pG�P ?fff�>��[�% :2ro�x�:-B� �>)���/u��|�P/nz�F�@ �%��6Dz$�$��/R/*����s� �^p� ��l?��/�?�?/ $/no$?6?H?Z?p?~? �?nO�O�O�?�?�?O  O2ODOVO�OF_X_�O�Oj\��OL/�_p/�/ �/�/�/�/�_j��_�_ {o�_�_	oo-o?o�o couo�o�o�o�o�o �o=�%;�?���	8��O�#s���� �q���`�����U ���R��₣���� �����Vz�Yw��V� ����h�޵������LϾ�Пܘ>����ܚ>�P�b�t� ��������Ώ���� 2�ԯ:�L�^�p����� m���ʟ��� ��$� F� �Z�l�Eϐ����� Ư��ꯨ�� �2�D� V�<�z���e߰��� ��߯�����2,,
��.�@�Q�0�i�2 d������������ ��/�6$-.P�{ћ� �	�
��]
�_ W/�1)����(D����_�����ы
w�7�>q�AݝR8�R#ӳ>L� �x#ϭ�B�<#�
ʱ��p�R�U��Q����7�v�z��j���@7Q�~r�A� 	�R��Z�i�:�\�B����5/V/h/ K/�/�/Q�;>��:0�/��It$ Z
?$[�>�
�/<7A��<?�/^??6�k +��̪5.�����5j$敕�5(4$��5�?�;�;��.�5>��yH
Ej5��EO8M�Y&Er�=�  BEj�SOy;	p?�O tO�O�G�?�O�O�O_�#_5_D[�$CCS�CH_GRP15 2���fQ�&� �\Z�]�  ғp^3�;�U �U���Qc�_�_�_oPfBo
n����pvu?333r�Rs|���D/  C���G�P ?fffr>[��vu�i�aο D؈_1r�}��r�g�y v/Yk�^�F��osx���pF@ �u0qse�pDz�` �����z������ ��o�o�o#� GQ��%���ʿ�� ��ŏ׏���-���� �U�g�y����������ӟ�ïկT�-�笸 g��?����#�5� G�M��,�>���b�t� ��������v���� �h�:�L�^�pϺ�h����~�X�j�|߆�� K��Р��zW0���� ��?�8���b ��� b_��z&o��� �ʌ���� �Ԕ�zZg� ��:f|��n?�x;�M�Y�>����� Y�����������'�  K�]�o���Q�� ����������5�G�  k�}�������}�� ���1Cqg %/������� 	�/-V߈�?,?>?T52�|�?�?�?�?�=�/�22�?
OO .O@OROdOvO�O�O�O �t�~�N�!$CiCj8, ���i�i�"�����/�y@f_x_�_�_�V$G0@�WH_ZY^1g�3�>��#o�-���#0e>Ly``a�*R�)O<#�
G'"p0o��R�p/�VR������Oe�b ge@ ��hd���/����@Fv��,���+B(! PeL����	����`>q�d�_�_n�^ESIt$ ��$�6K>��b
g���ADT���a�ۏ�����P+�{��'�.���3���Q$敕C�(4�$�O���;��=.{�>��H���Q�5����8M�	Y���M=``���R�!П��	���*�� c�U�j�|�������!��M��ħ   �"��b�d[r�`�� �J��h+�=�O�a��(x�f�R���c��?333�U'��T3Y�gqD/  C G�P ?fff�Q>�a4T����K�( 䯮��]�_��� ��������OU���)�<G*h�F@ [�g�ϵrh�Dz��|�g��Y�+���z1Z?L9 �7�I�[�m��E�� ��o������G��� !�3�I�W��G�Y�z� ������������/�@q�1����C��� %ߛI�[�m�ߑߣ� �Cb��T��� ��<N�r �����/��?`�ߴ/�/�/��ȧ� � �ry֧�/J>go1S �/�?k߲�po� �e �2|t�a�v�`_U_y/* �?2'x`/4�!֪�4AN�eo��8�$�%�L<�O�H>����$�J ?)?;?M?_?q?�?\_ �?�?�?�?O�_O%O 7OIO[OmOFo�O�O|o �O�O�O�O_�o3_E_ i_{_�_�_�_�_� �_�_oo/oSoeo >��o�l�/�/v�������2������*�		�B�2=�f�x��� ������ҟ����� �)�T�tt�����|�� ���r�����
�¯ ԯ����st��8��������d�P�q>�X!��vk�s���>Lհ���o���<'#�
�a�rp��+�ph�*�_���q@OuSq��C�dpõ@ ĴW"o���d���o�� ����Br5�B�q�� ���/�A�$�e�w�*{�>h���	��ߡ��It$ ��$4�>%��
���A�����7�����D�+��=̃�.�����C��$敕��(4$�ܫ�c�u�;��.���>��H��C�5�����8M�Y��K�=���C��q,�R�	I�b�M���q��� ����������}�#�|�   �r l 7�ķ��{c[� h<ȇ���?����_��a �O%?333K��L������D/  CppGÿP ?fffK�> 4���O%og�o�@ 
"o-w�K�Es)O�/ #/D/7u��+/�/�z�F@ �%�+k��DzY�$��/��/E*ց���� � ������?�	? �?�?G/Y/�oY?k?}? �?�?�?�?�O�O�OO O1OCOUOgOyO�O�O {_�__�O�\�_�/ �_�/�/�/�/�/�/o ���_�_�oo,o>oPo boto.�o�o<�o  �o(r 5p�6?0�"�4�>8�_L� Xs��2���ÿ��� ���U;���RL�;�� ��S���H����ɋzD� �w԰��L�2
�����4�C�G�����>���C��s� ��������͏ߏ��� �'�9�g�	�o����� ����ɟ�����ؿ#� 5�G�Y�{�5Ϗ���z� ůׯ���)����C� U�g�y���qϯ����� �7��@��������2a,?�Q�c�u��eߞ�2���������� 
��.�@�R�d�k$b. �������	�
��G]K K?�T_:Wd�f)0]Ty���Д P	����l�>�q��v��R�RX��>�L1X���w�<#�
����p���U8(߆����l��� �����@lQ  �r�v�>�OR<��GZ���oϑ�B��/ j/�/�/�/�/�/��p�>�Doe&?��I�t$ ??$��>�E
?q7A��q??�?=?O6� +��̞�5.����5�$�敕�5(4$�xE�?�;;��.3E�>��H?E�5{��OE8M�Y[E��=wE�HшO�;	�?�O�O�O�GO_ "_4_F_X_j_��W~>|W  K��p �h"p�U�U���Q ��_�_oo�B0onʻ���pM�u?3�33��R���!D�/  C��G�P_ ?fff�>� ���u�i�a�y؜_fr �}����g�y�/m ���{����� pF@ �q�e� pDz�`4���p�z2��� ��o %7��[e�'� 9�������Ǐُ� ��A����2�i�{� ������ß՟�)�ׯ�h�A����{��S� ��%�7�I�[�a�� @�R��v��������� п����Ϙ�*�|�N� `�rτ���|��ߒ�l�~ߐߚ��_��д� *)�WD����S�L� #��b8 '��Зs�4$ �S&�)�ʠ��� 0�ԨюZ{���o'f����?�O�a�m�>�����m����� ����)�;�_�q� �����e������� �%��I�[�4��� ������������! 3EW�{9/�� �����/A��jߜ�.?@?R?h52@�|�?�?�?�?�=�/�22�?O0OBOTOfO xO�O�O�O�O�t�~�N 1,$WiWjL,���i�i �"�����/�yz_�_�_�_�V+$[0�W\_nY(r1gC�>�7o��-.�#��#De>L��`ta�>R�)<#�	
[;"pDo�R ��/�VR���%!ce�b {e@ȡ|d� '�/����Zv��@���+B<!de`������/���`>� q�d�_�_��YSItk$ ��$�6>��b	
{�͇AXT͏u��x�����P+���;��.���G��Q$�{��W�(4$�c���-�;��.��>���H���Q5�=���8M�Y��]�=t`ӕ�R�!�
�	 ���>�)�w�i�~� ������Ư5�M��ا  �"$��b �dor�`3��Z ��h ?�Q�c�u�����z�R����c�?33�3e;�dGY{qD/�  C( G�P /?fffa>�aHT �'��_�(����'� /]o��+�������π��Oi���=�[*|�F@ o�{��#r|�Dz���{�m�?���8�1n?`9 �K�]� oρϓ�Y���߃�� ���[�#�5�G�]� k��[�m��������� ����1�C���3E����W���9߯]� o߁ߓߥ߷߽Wb� �h���, �Pb����� ��*/��(?���/�/�/��Ȼ�0#�y ꧠ/^>{oES�/�? �p�0�e�2�tq �v psUsyC*�?F'�` C41��4UN�e���8��$��9�L�O�H>����$�J+?=?O? a?s?�?�?p_�?�?�? �?O�_'O9OKO]OoO �OZo�O�O�o�O�O�O _3_�oG_Y_2}_�_ �_�_�_�_��_oo 1oCo)goyoR��o�l@�/�/������ą2� ��	��-�>��V�2Q�z�������ԟ ���
��#��=�h� �t�����|�����r ����֯���1��t��L���ʩ΁x�d�$q>l!��.�p����>L��б��/�<#�
�a�rp��?�|�>�s���$qcugq��W�xp׵@$شk"�� .��d�o������Vr'I�B�q����"�C�@U�8�yߋ�>{(�>|����'���ߵ�It$� ��$H�>���
��)�A��)���K��߼�X�+��̗�.������W�$�=���(4$ܿ�w�މ�;��.��>���H��W�5����8M�Y�_�=@а/�W� �@�f�	]� v�a����������������"1�$CC�SCH_GRP1�6 2����S&� �\G�/J�  �� K� ���(� ��o��Pȼ����S�	�s��u <�c%?333_���`�����D/  C��pG�P ?fff_�>H���c%�� �o1�u"�-��_�z �)c�F/X/y/Ku3���`/�/�z�F@ `�%�`��Dz� 4��/�/z*�ʏ�� �����/ �?4/>? OO|/�/�o �?�?�?�?�?�?O�O �O_BOTOfOxO�O�O �O�O_�_�_A__�\�T_�/,o�/�/�/? "?4?:o��o+o�oOo aoso�o�o�oc�o�o qU'9K]��U5��k?E�W�i�s8�8_���s��g�ێ ׿��,�%��Up�� b ��O�L���g��\�ϥ ���zy��w�����g
@T�Ҟ'� i�x�[���(�:�F�>��� x�F�����̏ޏ��� ��8�J�\�n���>� ����ȟڟ���׿"� 4��X�j�|�����j� į֯������0�^� T��x����������� ������l�C�u���+�A�2�,t���$�������2���� 	��-�?�Q�c�u��� ���$�.�����00 %�|]��t҉_oW�߀�)Se�����4��5G	K������>�q��b�R��>LfM�����<#�
4��p���U]߻����������<���T@�QU�r /��sĄR�q�3&|Z/�¤���B �=9/�/�/�/�/�/?�˥>�y���[?2It$ t?$���>�z
T?�7A�1�?N?�?r?�6� +����E.���� E�$敕0E(�4$�<E�?K;�{�.hE>��HtE��5���E8M�Y�E��=M�E�}ѽO�;	�?�O�O_ WPOB_W_i_{_�_�_�/���~�W  ���p��H"�e �U���Q�o*o<oNoP�BeoSn����p��u?333�b�| 	T!D/  C��G�P ?fff�>�!�u y�a8� ���_�r ���g� �/����Ű�B�x�4�UpF@ H�0Tq�e�UpDz�`i��TF���zg�G�9� �$6HZl2� ���\�n���4�� ��� �6�D�v�4�F� g�����ԟ���
���^�����v�0�� �����6�H�Z�l�~� ����0u���Aϫ��� Ͽ��Ͽ�)�;��� _ϱσϕϧϹ�߱���Ǐ�߳���ψ� ������_)�Wy�7�T �߁�X��bm \��� ���i$��&�LL) ����e����Z�� .��\f�����?/x������>����� ����(�:�L�^�p� I�������� � �$�6�H�Z�3~��� i���������  2/Vhz��� n/���
/@ R+?v�����c?u?�?�52�|�?�?�?OM�//B2*OSOeO wO�O�O�O�O�O�O�O �t�~^A1a$�i�j�, ح�i�i�"�˧�/�y@�_�_�_�_
f`$�0@%g�_�Y�1Qg=C�>E�lo=c�X��#ye>L�`�a�sR9O<#�
�p"pyo�bU��/fLR����<%@!�e0rQ �e@ ���dD�\?���@�vتu/" /";Bq! �e���.��R�d�+p>Uq�d o�_��^�SIt$ Џ$!FK>��b
���A�T����$�Ώ��1`+�{��p�.���|��0a$敕��(4�$ܘ�P�b�;��=.ĕ>��HЕ0a�5����8M�	Y�8]=�`�0b�!�?�	6�O�:�s�^� ������ůׯ���j�]���   �"Y�$r�d�rph�P� HZU�)xt�������,�(����LR�N��c<�?3338ep�9d|Y��qD/  C] G�P ?fff8a>!q}T<�\�T��
8 -���\�d]8o2�`�<� ���1�$%_���r�<�*��F@ �հ��Xr��DzF��԰����t�2��1�?�9 ܀ϒϤ϶��ώ��� �߸���4�FߐF�X� j�|���������� ����0�B�T�f�x�@��hz������ n���ߤ߶������� ��b���+ =Oa/��)/� /��//_/�]?`#��/?!?+���� 90E#�y��/�>�ozS �/�?�(��p�90(u B�t@q�v5p�U�yx* 1O{'�`x491�D�N u��!H044�n�L<�O�H>���04�J `?r?�?�?�?�?�?�_ �?OO&OTO�_\OnO �O�O�O�O�o�O�O�o _"_4_F_h_"|_�_ g�_�_�_�_oo� 0oBoTofoxo^�o�o ���o$|�/-?��я���2N�,�>�P�b�s�	R���2������ӟ ���	��-�?�Q�X� O�r����t���|4 8�8�,�A'Q�S�� �J�A�f��t쀁����������Yq>��!ȿc���E�յ�>L��EϢd�<'#�
�a�rpտt�p��s�����Yq@�u�q���­p�@Y Ġ"��c�+t<)�� 4
�ϋr\~�B�q�� ��W�xߊ�m߮���s{]�>��1�\�R��꣯It$ ,�$}�>%�2�
�^�A�^����*�<捰+��=���.����匱�$敕��(4$������;��.� �>��H,���5���<�8M�YH���=�d���5�u���	���������� ��!3EW��l�|D.i  8� � ��U� �]����� ������������� :Ø%?333�����ة��D/  C�pGÿP ?fff��> }�٤�%���of�� S"�-������)��Z/ l/�/�uh��t/�/�z F@  5!t�� Dz�!4/�/��/�*���� � �� //$/�?H/R? O&O�/�/�o�?�?�? �?�?�?.O�O�O_VO hOzO�O�O�O�O�O_ �_�_U_._�\�h_�/ @o�/ ??$?6?H?No �-o?o�ocouo�o�o �o�ow�o�o�i ;M_q�i5��?0Y�k�}��8�L_�� �s�{1���֣@� 9�e�%�b����`� !Ԝ�@֑����z�� �w�Ԅ��{
h��\�}�������<�N�Z�>�����Z��� Ώ�����(��L� ^�p�����R���ʟܟ � ���6�H�!�l� ~�����į~�د��� � �2�D�r�h�&ߌ� ����¿Կ����
��� .π�W����-�?�U�2�,�����������2����/�A� S�e�w��������$�. �����DD9ܐ]� ��ҝ_�W�߯)gy����H��IP[	_�	����>�q�$��bb��1>�Lza��+��<#�
H�(�p1�e8q�������� ��P�	�h@�Qi �r/�߇ĘR��G&�Z-/�¸���B)�QM/ �/�/�/�/
??�˹�>!���o?FI�t$ �?$��>��
h?�7AE�?b?��?�?�6� +��̞(E.���4E�$�敕DE(4$�xPEOK;��.|E�>��H�E�5{���E8M�Y�E��=a�E����O�;	�?_�O+_WdOV_ k_}_�_�_�_"/���~>�W  ��� ��\"� ee 
a �,o>oPobo�Byogn�����u?3�33�(b�4	h!D�/  C�G�P_ ?fff�>� 5�uyqL����_�r ���g��/�� �����V�*�H�ipF@ \�hq�e"ipDz�`}�hZ�,�p�z{�[�M� �8 J\n�F����p� ����H����"�4� J�X���H�Z�{���ğ ֟�����0�r� �2�����D��į&��� J�\�n���������D ����UϿ�ѿ���� ���=�O���s��ϗ� �ϻ����Ņ�ۏ�������Ȩ����� s)�W��K�h2�ߕ� l��b� p������}$ ��&�``)0���3� y0����Z��B��pf�����?&/������>����Զ��*� <�N�`�r��]��� �������&�8�J� \�n�G����}���� ���� �4F/j |�����/�� 0/Tf??�������w?�?�?�52@��?�?OO+M
?CB2>OgOyO�O�O�O �O�O�O�O	_��*^ U1u$�i�j�,��i�i �"��ߧ	?��_�_o�_ft$�09g�_�Y(�1egQC!>Yрo�=w�l��#�e>L��`�a��R9<#�	
��"p�o,bi��/+f`R��!P%T!�eDre �e@��dX� p?�����v쪉C"/6;B�!�e���0�B�%�f�x�++p>�iq�do
oˏ�SItk$ �$5F>��b	
ď�A�T���8�x��E`+��̄��.�����Da$�{����(4$ܬ��d�v�;��.ؕ>���H�Da5�=���8M�Y �L]�=�`�Db�!-�S�	 J�c�N���r�����ǯ�ٯ������$C�CSCH_GRP�17 2����@�&� �\4>��79  �"m�8rt�r p����\Z��=x����@Ϳ߿@����`R�b�y�cP�?333Le�Md�Y�qD/  �Cq G�P ?fffLa>5q�TPՑ� ���8b��p�x]Lo g�t�P�3�E�f�8% _���Mߧߤ*��F@� ����M�lr��Dz {������ߩ�g��1�?�9 ܵ������� ����!�+�����i�{� �{��������� ������/�A�S�e�w� ����������.��A�������� ���!�'�b� <N`r��P/� �^/�B//&/8/J/ �/B�q?X�2?D?V?`��%n0z#�yT�
? �>�o�S?O�]��p �n0<u9B�tTq�vIp �U�y�*fO�'�`�4n1�T�AD�Nu�VHe4�H��\'_3X>���e43Z�?�?�?�?�? �?O�_%O7OIO[O�O +o�O�O�O�O�O�O�o _!_�oE_W_i_{_�_ W�_�_��_�_oo KoAo�eowo�o�o�o ��o�o��Y|0?b?���.�2��a�s�H����������2�� �����,�>�P�b� t����Ԅާ�ҁ�t� ��im�m�a�v\ ����@�R��v����t!���"�4�8��Γ�q>�!������z�
�>LS�:�z<���<#�
!q��p
ϩ��J���ݢ���q�u�q)����pA�@�B��"�Ϙ�`t q^ �i
��r���B�*�&ߌ߭߿ߢ����ߨ{��>��fđ�x��H��It$ a�-$��>�g�
A��A���;��_�q�°�+����.��y����$敕��(4$�)�����;���.U�>��H�a���5��q�8'M�Y}�ɭ=:�����j�����	������ ��=�/DVhz����$CCSC�H_GRP18 �2�����&� \���v/��   m�� ��5Ғ� ٪��&8J\��(saݢ�� o��%?333ɵ"ʴ��A�D/  C�pG�P ?fffɱ>����%)!%�� ��"�-��ɿ��)�� �/�/�/�u��P/�/$?<!�c F@ V5b!���c Dz�w4b/�T?&?�*T�4�&� �2/D/V/h/z/@O�/ �?jO|O�/�/!�?
O O.ODORO�OB_T_u_ �O�O�O�O�O__*_@l_o,o�_�_>l��_  ?�oD?V?h?z?�?�? �oo�oO�o�o�o �o�7I�m �������5�`�?����ӏ�8Ȣ_ ��sL����E�A�� ����fe�Z�jb뀹� ��V���u���9�9�*� �-�R�*���
��<���jӘ����ϒ�<����>���ℰ� �$�6�H�Z�l�~�W� ����Ɵ؟���� � 2�D�V�h�Aό���w� ¯ԯ������.�@� �d�v�����ȿ��|� �����*��N�`� 9���̭�ߏq�����2 <������%�	�=�28�a�s��� ������������
4 >$O�oԚ����] �����_�W�9� ���n���3���	��_K��>�S�z�qbfb�Ӈ�>L���ρ�<'#�
��~�p�&pce��%Z���@J�NѦ>"_о@a �R�j/����R�ϝ& �Z�/=��0�Bѧ �/	?*?<??`?r?%� >c!��?��It$ �?$/�>%��
�?GA�O�?2O�?�6?+��=�~E.����E>�$敕�E(4$�ܦE^OpK;��.��E>��H�E>5����E8M�Y�EF=�U>��'_MK	DO]_H_�_lW�O��_�_�_�_�_	ok��$CCSCH_G�RP19 2����:a&� \.��1�  ��g�2" $�" �eeV
�a7( �o�o�o�o:R�o�nZ��\��J�?33�3F�bG�	�!D/�  Ck�G�P /?fffF>/!� J��y�q���\o�j� rFawn�J?-�?�`��2��G������pF@ Ӆ�qGuf"�pDzup��я��a�8���� ܯ� ������%���� c�u���u��������� ϟ���ѯ�)�;�M� _�q�������鯗���(�����;������ ӏ���	��!Ϛ � ���6�H�Z�l�~ϐ� Jߴ���X���<�� � 2�Dߎ�<�k�R�,�>�P�Z���h�t��) Ng������� Wr� �h�6%3��$N! �&C ��)��`���� ��h�Nj;���%�fP��_�BO|/!->���_�-
���� ����������1�C� U���%���������� ���	�?Qc u�Q/���/�� E;�/_q� ���/���?/S,@*�\��? OO(E2}� [OmOO�O�M�?�B2�O�O�O__&_8_ J_\_n_�_��~��^�1 �$yz<c�gygy[2 p�V��?��:oLoyopo�f�$@�go.i2A�g�C�!>���o�=p��t3u>LMp�4qt/�R�9<#�
!�"p�b�D?�f�R���!�%�!#u�r� ;u@��<t��� �?Z$k�X/�c� ��"�/�;B�!$u �����@����ݏ+�p>�q�`t�o�oB�cIt$� [�$�F>�ar
;���Ad��5���Y��k��`+�����.������a$�=��(4$�#�۟��;��.O�>���H[��a5���k�8M�Yw��]=@4p���bd1��ʛ	�� گů���7�)�>�P��b�t������$CC�SCH_GRP1�A 2������&� �\�>p߮9  g2�Яr�t/��p ����Z��x �2�DϠVϷ�m�[��R���<is��?333�e���di;�D/  C�� G�P ?fff�a>�qd��� � /�8ٿ�����]�o�� ��Ǐ�߼��߯%�_J�����:]�F@ `P�\����r]�Dz�� q�\�N� ���NA.O I �,�>�P�b�t� :��ߢ�d�v�����/ ����(�>�L�~�< No����������  $f&�~8���>�P�b�t� ���r}�I/� ����/�/1/C/ �/g/�/�/�/�/�/?����?��?�?�?��Ȝ�0�#F�˷�??N ;c�?�O`��T�d �0�u�BP��qo��p3e 3�$:�O'7Lp$D�1˺@�D6^�ud��H�4�����\�_�X>��� �4�ZOO0OBOTOfO xOQo�O�O�O�O _�o __,_>_P_b_;�_ �_q�_�_�_�_o� (o:o�^opo�o�o�o �ov��o�o $
� HZ3�~�|�?�?k�}�����2��؟���$����7�22�[� m��������ǯٯ� ������I�i��ɔ� �������؂������ٷ�ɿ����h����-Ǚ�����Y�E��>M1t��k`���>L�����{���<#�
�qx�p��� �]���T����D�H���8�Y���@��L2d���t������
}�7��*�B y��ŝ��$�6��Z�l��	�>]��������It$ ��$�)�>���
��
�A���
���,�����9�+����x�.������8�$敕��(�4$ܠ�X�j�;�{�.��>��H���8�5����8M�Y��@�=��8��!G�	>�WB{ f���������$CCSCH�_GRP1B 2����4&� \(�|�/+�  � a0,�Ԭ�	БyP� ~1؝���4���T��V0��D5?333@řAĄ����D/  Ce�GÿP ?fff@�> )х�D5�)}!��V �"d=l�@�['h9D�'? 9?Z?,���/A?�?��� F@ �5�!A%`�� Dzo �4�/�?��?[:ˑ���� � �/�/�/�/�/�O?O �O�O]?o?�oO�O�O �O�O�O�O�_�_�_#_ 5_G_Y_k_}_�_�_�_ �o�o"o�_�l�5o�? �?�?�?�?OO ���o�0BTf x�D���R��6� ��,�>���6Ee�LO0&�8�J�TH�ob� n���H�����ς�� ��eQ"���bb�0�-� ��H���=а��١�Z� ������b�H5�����J�Y�<�v�	��'�>���Y�'��� ������џ���ο� +�=�O�}�υ����� ��ͯ߯������9� K�]�o���Kߥ����� ۿ����?�5���Y� k�}Ϗϡχ����ϰ� ��M�$�V������"��2w<U�g�y�����{��2��������  2DVhz�4x> �����)*�]ma) a)U�joPgz�|94Fsj����P(,������>ʁ�����b�bn��>�LG .!n����<#�
���p���e8>�������� ��%�"��5%@�a6$ ɂ�/��T�ebR�6]j�/�҅ߧ�B��%? �?�?�?�?�?�?�ۆ �>�!Z$�{<OI�t$ UO$��>�["
5O�GA�O/O�OSOeF�+��̞�E.���U�$�敕U(4$�xU�O�K;��.IU�>��HUU�5{��eU8M�YqU�=. �U�^�_�K	�O�_�_�_�W1_#o�8oJo\ono�o�k�$�CCSCH_GR�P1C 2�����a&�� \��j���  a�ހ�"~$ )2� u�e�
�a�(�,>P�RgU~���Ӏc#��?333�r�51D/ � C��G�P ?fff�>�!�� ��qߏ��o|��� ��w��?����׏����D�����W�F�@ J�V��u�"W�Dz�pk�V�H��؊H�(�� �&�8�J� \�n�4�����^�p�ڏ ������"�8�F� x�6�H�i�����į֯ �����`�� ϟ�x�2̸�����8�J� \�n�������"wω� C߭Ͽ���������� +�=���a߳߅ߗߩ� ��ﳕ��ɟ�����јȖ�����@9�g {�9�5/����Z��r N0^���%��J4�!i6 � --9���!�F � ���j��0�%^v������O�/���>�����
��*�<� N�`�r�K�������� ���&8J\ 5/��k/���� �/"4?Xj| ���p?���/ /?B/T/-Ox/�,�� ��eOwO�O�E2��O��O�O_]�?1R2 ,_U_g_y_�_�_�_�_ �_�_�_����nCAc4 �y�z�<ڽ�y�y�2� ͷ�?���o�o�o�ovb4�@'w�o�i�ASw
?S�!>G�n	Me�8Z��3{u>L�p�qx�/ub
I<#�
�!r2p{rWŻ?vNb���!>5B1�u2�S0�u@���tF�^�	O �$��/��ںw�12?$KBs1�u�����0� �T�f�;�>W��t��o���cIt$ Zҟ$#V>��r
���A�d���&�П��3p+���r�.����~�2q$敕��(4$ܚ�R�d��;��.ƥ>��yHҥ2q5���O8M�Y�:m=�p 
�2r�1�A�	8�Q� <�u�`�������ǿٿ������$CCS�CH_GRP1D 2���.��&� �\"N��%I  �2[�&��t����� s�Jjx�+��ϩϻ���P.�����Nb�P��s>�?333:u��;t|~i��D/  C_0�G�P ?fff:q>#�d>��wі/ HP���^�fm:U�b� >�!�3�T�&5o��;�x��:��F@ ��0��;�Z���Dzi��������U��A�O�I ܣߵ������߱� ������W�i�/i� {������������� �/ASew��������� /��/���������� �/�r�/�/*/</ N/`/r/�/>?�/�/L? �/0???&?8?�?0��_OF� O2ODON�� \@h3��B��?�N� |cO _�K�ˀ�\@ *�'RǄB��7��e�� �:T_�7�p�D\AB�/T �^���DXSD6�p�xlo!h>���SD !j�O�O�O�O�O�O�O �o_%_7_I_w__ �_�_�_�_�_��_o �3oEoWoio�oE��o �o���o�o�o9/ �Sew����� ����G�OPO�����2q�O�a�s�����u���2��ү� ����,�>�P�b�t� {�r������ � W[�[�O�dJt�v�@.�@�m�dω�߄�@���"�&��Ǽ�|�>�1�φ���h���>LA�(�h�򲇙O<#�
��p������8���˲���|�����կ�Ѐ/�@ |0��2�߆�N�_L�@�W�߮����B�� ��z������������>��T��u�6�^�It$ O�$��K>�U�
/���A����)���M�_���+�{����.�����ޯ�$敕(4�$�����;��=.C>��HO���5��_8M�	Yk��=(Ї��X����	������ +2DVhz���$CCSCH_�GRP1E 2�����?&� \��d?>��  [��0 ��x�#��%�Ǻ� ��/&/8/J/�a/O.�˲��0]ӻ5?3�33��"����/�D�/  C܀G�P_ ?fff��>�� ���5�)�!����v2 �=㽷��'�9��?�? �?����>?�?O�Q0F@ DEP1�%��Q0Dz� eDP?BOOp�:B�"�� � ? 2?D?V?h?._�?�OX_ j_�?�?��O�O
__ 2_@_r_0oBoco�_�_ �_�_�_�_ooZo�oro,|��oO� 2ODOVOhOzO�O�� q�=������ ���%�7�ɏ[���� ���������Eܟ�O�������HȐoِ� :�u�3�/�����}� Tu�"H�Xrِ�դ�D� ��c��'�'��ѯ� @��ّ���*��X&��Д���߀�����>���Д�� �� $�6�H�Z�l�Eϐ��� ��Ư������� �2� D�V�/�z���e߰�¿ Կ�����.��R� d�vψ϶Ϭ�j����� ������<�N�'�r߀�ܛ�͟_�q�����2@�<��������+2&Oas�� ������4�> =�]�)�*}��m�)�) ���o�g���9����&\���!'��(��M'9��>A�h/��_rTr��u%>L� �!��o�<#�	
��l�pu/"Qu��&H����8�<��%,2M�%@�a�$@� X?����b�ߋ6�jq?+����Bm�%�?�?�O*OONO`O�� >�Q1�$���O�Itk$ �O$>��"	
�O�GA��O�O _x�O�F- +���lU�.���xU,!$�{���U(4$ܔU�L_^[;��.�U>���H�U,!5�=��U8M�Y�U4�=� e,"��o;[	 2_Ko6oooZg�_�o�o��o�o�o�o{�$C�CSCH_GRP�1F 2����(q&� �\���  ��U� 2�$�2 � �umuDrq%8��@��(b��~H�J�y�#8�?3334%��r5$x�1D/  �CY�G�P ?fff4!>1y8�y� q����J�X�`4/ O�\�8O�-�N� �໏5�����΀F@� ��́5�T2΀Dz c��͏����O������ ܝ�����ӏ 叫�	��կ�Q�c� ��c�u���������� ������)�;�M�_� q�����׿�ϗ����̸)ϋ�߯���ӟ ���	�߈"�� ߺ� $�6�H�Z�l�~�8�� ��F���*���� �2� |�*�Y�@��,�>�H���V�b�9<w�� ���/v�����E��0 ��V�$5!�4<1�610 ��9��N�� ��V�<z)��%�v>M��0_j?�>���M�}��������� �����1Cq /y������/ �	�/-?Qc� ??���?���/ 3/)/�?M/_/q/�/�/ {?�/�/�O�/A<�J��O�O _U2k�I_[_Hm__�]oO�R2�_ �_�_�_oo&o8oJo \onou�l��n�A�4� ��<Q�U�U�IB^�D� nOp�(:g^�v�4	P�w
y Q�w�Sv1>����M����bC�u>L;�"�b?<�b�I<#�
	1�2�p��r��2O�v�b��v1�5�1����0)�@v�*���Տ�OH4 Y�F?�Q�2y?�KB�1��t�������˟ݟ�;z�>΁N�yxo0�sIt$ I�-$�V>�O�
)�{�At{�#���G�Y��p�+����.��y����q$敕��(4$��ɯ۫;���.=�>��H�I��q5��Y�8'M�Ye��m="����rRA����	��ȿ�� �׷%��,�>�P�b��tσ��$CCSC�H_GRP1G �2������&� \��N^�I   UB����r��z���� �j����� �2�Dߥ�([�I��b���W���?333�u
Ҳt�i�)�D/  C�0G�P ?fff�q>���d������?�H ��p����m����鵟 �����5�o8���<	JK�F@ >�J���тK�Dz��_�J��<����<Q_Y ��,�>�P�b�(�� ��Rd����	?���� ,:l*<] ������ @T//�l&,�� �~/,�>�P�b�t��� �/�k/}/7?�/�/�/ �/�/�/�??1?�?U? �?y?�?�?�?�?���O`���O�O�O��Ȋ �@�34���oO-^)��c ~Ow_N%��B�R"�@�� �R>���]���!u!�J �_G:�T�A�ʦT$ny�RֻX�D���zl<�o�h>����D�j �O__0_B_T_f_? �_�_�_�_�_��_o o,o>oPo)�to�o_� �o�o�o�o��( �L^p���d� ��� ����6�H� !�l����O�OY�k�}���2��Ưد����	�%�2 �I�[�m� �������ǿٿ��� ���7�W��ق�w�� ����ƒ������ ������ �V���נ�ϙɝ�G�3��>�;Ab���Y"N"ߓo��>L�П�ߏi���<'#�
��f�po��pK%���B����@2�6���&�G���@� ��:BR���ń�Ï�� �k�%����Bg��� �����$��H�Z����>K������ϭ��ïIt$ ��$�>%���
����A����������'�+��=�f.���r&��$敕�(4$�܎FX;��.��>��H�&�5����8M�Y�.�=���&�ϑ5	,E0iT�������� +��$CCSCH_G�RP1H 2����"!&� \��?�  ҒO@� �Ԛ���%g%>�l!� �/�/�/�/"�/�.B���D@��2E?33�3.Շ"/�rɦ�D/�  CS�G�P /?fff.�>�s� 2Es9k1�� �D/�2RM Z�.�I7VI2�O'OHO��ϵ?/O�O���0F@ �E�1/5N��0Dz]0�D�?�O�OIJ8������ ܗ?�? �?�?�?�_O_�_�_ KO]O��]_o_�_�_�_ �_�_�o�o�oo#o5o GoYoko}o�o�o��o�|�#�O��O �O�O�O�O_	���� ����0�B�T�f�x� 2�����@�ҏ$���� �,�v�$US�:_�&�8�BX�P�\��� 6'쟪���p������u ?2���rP�����6� ��+��Ş鏚H����� ��P�6*#������&8��G�*d���	��>���G��w����� ����ѯ㯼���+� =�k��s��������� Ϳ������'�9�K� ]��9�ϥ�~����� ����-�#���G�Y�k� }ߏ�u���ߞ���;�@�D�������2eL CUgy�i��2�����  2DVhoDfN��� ���)�*��K}O9O9C� X>wh�jI"/4/a/X/}&�� �'/)�'�p�>���/z�p�r�r\��%>L50�1\��{�<#�
���p�/�"�u,��&���p���5�2��#5@pq$4���? z�B�Sr@�FKz�?��s��B��5OnO�O@�O�O�O�O��t0>�1�H4s/i/*_#It$� C_$�>�I2
#_uWA $u__�_A_�SV� +����U.�����U�!$�=��U(4$�e�_��[;��.7e>���HCe�!5���Se8M�Y_e�=@0{e�"L�o�[	�_ �o�o�o�go&8�J\n}{�$CC�SCH_GRP1�I 2�����q&� �\��X���  O�̐�2l4Bt0 �u�u��q�8��,��>��bU�C�����<Q3��?333�%���$�#AD/  C���G�P ?fff�!>�1������ �}��j�ϝ��/Ƈ ә�O����ş��2����E�F@ `8�D����2E�Dzڀ Y�D�6��ƚ6	 ��&�8�J�\� "�����L�^�ȟڟ� گ����&�4�f�$� 6�Wώ�����Ŀֿ� ���N���ߍ�f� �����x�&�8�J�\� n������"e�w�1�� �߿������߯��+� ��O��s������������������Ȅ�����.I�wi�' #?�x�qHռ�<@L� ��5�8D�1WF�0% I���40��z@�s5L�����_��?t��>��� �����*<N `9/������/ �&8J#?n �Y?������? /"/�?F/X/j/|/�/ �/^O�/�/�/�/?�? 0?B?_f?�<����S_e_w_�U2��_�_�_$�_m�Ob2oCo Uogoyo�o�o�o�o�o �o��~1QQD|�|� qL��̉̉�B�ϻ��O�癟����vPD��P���y�QA�-c�1>5�\��MS�H��Ci�>L�����?cr��I<#�
�1`Bp�i��EթO�<r���1,E0A�� �A@��@����4�L��O�4��?���e�B�?[B aA��������B�T�K�>E�ń�����~sIt$ ��$�f>�Ƃ
���A�}t򯚯���Ц!�+����`�.����l� �$敕|�(�4$܈�@�R�;�{�.��>��H��� �5��е8M�Yܵ(}=���� ��A	�/�	&�?�*�c� Nǜ��ϣϵ�����������$CCSCH�_GRP1J 2�����&� \^|��Y  �B I��鄔��y�a�8z f���ߗߩ߻���ߔ��<r�>�΃,�?333(���)�ly���D/  CM@GÿP ?fff(�> �mt,�m�e�?�H>� ��L�T}(�C�P�,�� !�B�E�o��)����J��F@ ����)�H���DzW���������C��Q�_�Y � ���������� ��E�W��?Wi{ ������� /ASew�� y/�/
/��,�/� �/������������? |��/�/�??*?<?N? `?r?,O�?�?:O�?O �?OO&OpOM_40_ _2_<�/JP VC��0��O�^��js�O �_�%9⹐�"JP�b ��0�Ԗ%��u���JBo �G���TJQ0�d�n����2hAT$�^��lx>���ATzq_ �_�_�_�_�_�_�o o%o7oeo�moo�o �o�o�o���o�o֏! 3EWy3���x� ����'��۟A� S�e�w���o������� �5�_>_Я���
��2_�=�O�a�s���c���2����ҿ��� ��,�>�P�b�i�`� �ή�Δ�����E-I� I�=�R/8'b�d��.�[�R�w�͔������P���ת�j�>�A���t��"�"V���>�L/��V���u�<#�
��ݒp�߅��%8&��ֹ���j��� ���⾐�@j!� �B��t�<�M":���E*�m���Bޑ�� h�����~�������n��>��B�m�c�$��I�t$ =$��>�C�
oA��o�;M��+��̞�.������$�敕�(4$�x��;��.1�>��H=��5{��M8M�YY��=�u��F���	�����/� /2/D/V/h/w+�$�CCSCH_GR�P1K 2�����!&�� \��RO��  I��@��f� �n��%�%���!��?�?&?8?�O?=>����@K�E?333���"�����D/ � CʐG�P ?fff��>���ĩE �9�1�w��/dB�M�� ���7�I���O�O�O���y�,O�O _��?@F�@ 2U>A�5��?@Dz�0ST>O0__�J0��� �O O2O DOVOozO�_FoXo�O �O���_�_�_
o o.o `o0Q�o�o�o�o �o�o�oH���`����Or� _2_ D_V_h_z_����_�q� +�������ˏݏ� �%���I���m���� ��ퟛUʯ�_�������X�~Ǡӓ(��' c�!����r�k�B��2 6�F�Ǡ�咲2���Q� �������	�.�� ǡ�*���m�F6��������ǹό�>�������� ��$� 6�H�Z�3�~������� ⿄����� �2�D� �h�z�S�ϰ����� �ϰ�
����@�R�d� vߤߚ�X��������� ���*�<�`�쉯 ��M_q�2�L�������2 =Oas��� ����D�N .+K� v9v:k��}�9�9��� �w���I�/�/�/�/�&J�z 7{/�)�;7
'��>/�V?��M�8B���c5>L�0�1x��]"��<#�
z�Z�pc?2?���66"����&�*�5B;�5@�q�4.�FO�� ���r��yF�z_O���B[�5O�O__ �O<_N_��0>?A�4��/�/�_x#It$ Z�_$>��2
�_�WAw$�_�_o�_�V�0+���Ze.����fe1$敕ve(4$܂e:oLk�;��.�e>��yH�e15���eO8M�Y�e"-=�0 �e2��)k	 o9 $]Hw�o���� ��$[