��  I��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT�&2�*  � �����$$CLA�SS  ���������� V�ERSION��  �5~�IRTUAL���'  1 �� T���C?R-35iA��� � aiS1�2/4000 8�0H
H1 D�SP1-S1��	P01.00W,  	� v��
�  ��}# :�������� {�F��2r9  �9����� HH��  ������ ����  C ���Z 
t
t������ ���s 1�2���?�u��|�u3��	8����&���<
= ^ ����� J����hI����;� 2 ������H�a����~#�	� � � !� ��� :�?8���'by�c/�/�/�/?��?;?;(X?xj?|?��1�3C( � �b����II2.����>�����wm"��܎?�?"4�<N*`6i2|2��~� ����׶����{���4�	���� @l� 
����n�m ��'!!%�F��� �34��=���!�	����;	':+�}J V 
��R �UV$jO����;��z'��-  � ���(%c	�	`� �#o
��%z�'� �
B_�_�_�_0�_$?�_��3�_o�+o=o��4����<��.����L.�m5�����;7������;G 	EFo�o���c\�?Sb8gBw3|b@ORK ��&����p�tG�p���}S�8HB\P��@�.��+; I'7A7�a#y����2B+�0�����+;= �x":+��� ����� �X"��o�� w��Z2X���w��)�()B�"�� d�#c A���#:rY:q�K�]�o����_ �� oɏۏ����#�@5�G��&�B�oR�bW4/5!A4�k4|�4�ov����ϓ�H�X�!2�D���K9�9~�5
�� �������l� ����0��%'��S@A�S��u� ����� 5V$�b�(S ���z#V@���� c�XR7 (�t Z�ֲ#rY�!����'�9���]���fd���������0ѿ����6d�N�biSR1C��x5|}����˚p�`�Mn����tG���������"�� D@��r�X��$� b*�<����#  z�  �V$�rA� ����Y���PB������`�(Ư%�ZP2Σ_� A��$�rZT�C߻������� L��p�9�K�]�o��������;" �R	@�r6|�h�z�j�̜`R=V����������� �����Ͻ���U`� ���x�V$����C�|�Cz#� ���O���;�( |ߎߠ�i{���� ����/A�Sew�����xTa��Ng%�	�,��� �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
??.?@?P<�P?t?�? �?�?�?�?�?�?OO (O0C��FO��� �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_o^?&o8oJo \ono�o�o�o�o�o�o 6OhOZO#~O�OXj |������� ��0�B�T�f�x��� ����
o������� ,�>�P�b�t������o ����*<N�(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�ȏ������ƿؿ� ��� �2�D�V�ҟğ n�����������
� �.�@�R�d�v߈ߚ� �߾���������*� ��N�`�r����� �������^ϐς�K� �ϸπ����������� ����"4FXj |�����2�� 0BTfx� ������R�d� v�>/P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?��?�? �?�? OO$O6OHOZO lO~O���O/"/4/ �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRo�?vo�o�o �o�o�o�o�o* �O�O�Os�O�O�� �����&�8�J� \�n���������ȏڏ ���Zo�4�F�X�j� |�������ğ֟�D � �z��f�x��� ������ү����� ,�>�P�b�t������� �������(�:� L�^�pςϔϦ�"�� ��8�J�\�$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ֿ�����������
� �.�@�R������ϛ� ���������* <N`r���� ���&��8 \n������ ��/l�5/(/���� ���/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?@OO ,O>OPObOtO�O�O�O �O�OJ/</�O`/r/�/ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�?�o�o�o �o 2DVhz �O_�O�_0_�
� �.�@�R�d�v����� ����Џ����*� <�N��o`��������� ̟ޟ���&�8�� ]�P������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� �h�0�B�T�f�xϊ� �Ϯ���������r�d� ߈�����t߆ߘߪ� ����������(�:� L�^�p������� &��� ��$�6�H�Z� l�~�������0�"��� F�X� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/���/x/�� �/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4O�XOjO |O�O�O�O�O�O�O�O __�/�/6_�/�/�/ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�oNO(: L^p����� &_X_J_�n_�_H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� �����o��ԟ���
� �.�@�R�d�v���� �����,�>���*� <�N�`�r��������� ̿޿���&�8�J� \ϸ��ϒϤ϶����� �����"�4�F�¯�� ^�د����������� ��0�B�T�f�x�� ������������� v�>�P�b�t������� ��������N߀�r�; �ߨ�p����� �� $6HZ l~����"�� �/ /2/D/V/h/z/ �/�/�/�/�/BT f.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O��O�O �O�O�O__&_8_J_ \_n_�/�/�_ ??$? �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0B�Ofx� �������� v_�_�_c��_�_���� ��Ώ�����(�:� L�^�p���������ʟ ܟ�J �$�6�H�Z� l�~�������Ưد4� ���j�|���V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �����������*� <�N�`�r߄ߖ��� ��(�:�L��&�8�J� \�n��������� �����"�4�F�X�j� �ώ������������� 0B�����ߋ �������� ,>Pbt��� ����//r�(/ L/^/p/�/�/�/�/�/ �/�/ ?\%??�� �~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O0/�O
_ _._@_R_d_v_�_�_ �_�_:?,?�_P?b?t? <oNo`oro�o�o�o�o �o�o�o&8J \n���O��� ���"�4�F�X�j� �_�_�_��o o��� ��0�B�T�f�x��� ������ҟ����� ,�>��P�t������� ��ί����(��� M�@���̏ޏ����ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��X� �2�D�V�h�z� �ߞ߰�������b�T� ��x�����d�v��� �����������*� <�N�`�r��������� �����&8J \n���� ��� 6�H�"4FXj |������� //0/B/T/f/��x/ �/�/�/�/�/�/?? ,?>?P?�u?h?�� �?�?�?OO(O:O LO^OpO�O�O�O�O�O �O�O __$_�/H_Z_ l_~_�_�_�_�_�_�_ �_o�?|?&o�?�?�? �o�o�o�o�o�o�o
 .@Rdv�� ����>_��*� <�N�`�r��������� oHo:o�^opo8�J� \�n���������ȟڟ ����"�4�F�X�j� |������į֯��� ��0�B�T�f�x�ԏ ����
��.����� ,�>�P�b�tφϘϪ� ����������(�:� Lߨ�p߂ߔߦ߸��� ���� ��$�6ﲿ�� N�ȿڿ쿴������� ��� �2�D�V�h�z� ��������������
 f�.@Rdv�� ����>�p�b�+ ���`r���� ���//&/8/J/ \/n/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?��?�?2D VO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�/�_�_ �_�_�_�_oo(o:o Lo^o�?�?vo�?OO �o�o $6HZ l~������ �� �2��_V�h�z� ������ԏ���
� fo�o�oS��o�o���� ����П�����*� <�N�`�r��������� ̯ޯ:���&�8�J� \�n���������ȿ$� ��Z�l�~�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �������������� ,�>�P�b�t����� ���*�<���(�:� L�^�p����������� ���� $6HZ ��~������ � 2�����{ ��������
/ /./@/R/d/v/�/�/ �/�/�/�/�/?b? <?N?`?r?�?�?�?�? �?�?�?LOO�� �nO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_ ?�_�_ oo0oBoTofoxo�o �o�o*OO�o@OROdO ,>Pbt��� ������(�:� L�^�p����_����ʏ ܏� ��$�6�H�Z� �o�o�o���o؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.���@�d�v����� ����п�����t� =�0Ϫ���Ο�ϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� ��H��"�4�F�X�j� |��������R�D� ��h�zό�T�f�x��� ������������ ,>Pbt��� ����(: L^p������ &�8� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?�h? �?�?�?�?�?�?�?
O O.O@O�eOXO�� ��O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oop?8oJo \ono�o�o�o�o�o�o �o�ozOlO�O�O�O |������� ��0�B�T�f�x��� ������ҏ.o���� ,�>�P�b�t������� 8*�N`(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�ڏ����ƿؿ� ��� �2�D�V�h�ğ �π���������
� �.�@�R�d�v߈ߚ� �߾���������*� <`�r����� ��������&��ϔ� >������Ϥ������� ����"4FXj |������� V�0BTfx� ����.�`�R�/ v���P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�? �?�? OO$O6OHOZO lO~O�O��O�O"/4/ F/_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodo�?�o�o �o�o�o�o�o* <N�O�Of�O�O_ �����&�8�J� \�n���������ȏڏ ����"�~oF�X�j� |�������ğ֟��� V�zC���x��� ������ү����� ,�>�P�b�t������� ��ο*����(�:� L�^�pςϔϦϸ�� ����J�\�n�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ��述���������
� �.�@�R�d�v����� ����,���* <N`r���� ���&8J ��n������ ��/"/~�����k/ �����/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?RO ,O>OPObOtO�O�O�O �O�O�O</_�Or/�/ �/^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�oO�o�o �o 2DVhz ��__�0_B_T_ �.�@�R�d�v����� ����Џ����*� <�N�`�r��o������ ̟ޟ���&�8�J� ������ �ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��z�0�T�f�xϊ� �Ϯ����������d� -� ߚ������ߘߪ� ����������(�:� L�^�p������� ��8� ��$�6�H�Z� l�~���������B�4� ��X�j�|�DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�� ���/ (�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFO�XO |O�O�O�O�O�O�O�O __0_�/U_H_�/�/ �/�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o`O(: L^p����� ��j_\_��_�_�_ l�~�������Ə؏� ��� �2�D�V�h�z� ���������
� �.�@�R�d�v����� �(���>�P��*� <�N�`�r��������� ̿޿���&�8�J� \�n�ʟ�Ϥ϶����� �����"�4�F�Xߴ� }�p����������� ��0�B�T�f�x�� ������������� ,���P�b�t������� ���������߄� .�ߺ��ߔ��� �� $6HZ l~������ F�/ /2/D/V/h/z/ �/�/�/�/PB? fx@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O��O �O�O�O__&_8_J_�\_n_�_�%�$SB_R2 1 5�P� T0 � ' C?7 �_�_ �_o o2oDoVohozo@�o�o�o�o�o�Q�o �_!3EWi{ ��������o � A�S�e�w����� ����я�����+� �O�2�s��������� ͟ߟ���'�9�K� ]�@���d�����ɯۯ ����#�5�G�Y�k� }���r�����׿��� ��1�C�U�g�yϋ��ϯ��Ϥ�~�_���� �!�3�E�W�i�{ߍ� �߱������������ (�:�L�^�p���� �������� ����� H�Z�l�~��������� ������ 2D(� :�z������ �
.@Rdv Z������/ /*/</N/`/r/�/�/ �/��/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�/�?O"O4OFO XOjO|O�O�O�O�O�O �O�O_�?0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>o"_boto�o �o�o�o�o�o�o (:L^pTo�� ���� ��$�6� H�Z�l�~������Ə ؏���� �2�D�V� h�z����������� ��
��.�@�R�d�v� ��������Я���؟ �*�<�N�`�r����� ����̿޿���&� 
�4�\�nπϒϤ϶� ���������"�4�F� X�<�|ߎߠ߲����� ������0�B�T�f� x��n߮��������� ��,�>�P�b�t��� ������������ (:L^p��� ������$6 HZl~���� ���/ /D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?6/v? �?�?�?�?�?�?�?O O*O<ONO`OrOV?h? �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�O �O�_�_�_o"o4oFo Xojo|o�o�o�o�o�o �_�o0BTf x������� ��o,�>�P�b�t��� ������Ώ����� (�:��^�p������� ��ʟܟ� ��$�6� H�Z�l�P�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ��ϴ���� �*�<�N�`�r߄ߖ� �ߺ����������&� 8�J�\�n����� ���������"��� X�j�|����������� ����0BT8� J�������� ,>Pbt� j�����// (/:/L/^/p/�/�/�/ �/��/�/ ??$?6? H?Z?l?~?�?�?�?�? �?�?�/O O2ODOVO hOzO�O�O�O�O�O�O �O
__ O@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo2_ro�o�o �o�o�o�o�o& 8J\n�do�� �����"�4�F� X�j�|��������֏ �����0�B�T�f� x���������ҟ��ȏ ��,�>�P�b�t��� ������ί���� ��:�L�^�p������� ��ʿܿ� ��$�6� �D�l�~ϐϢϴ��� ������� �2�D�V� h�Lόߞ߰������� ��
��.�@�R�d�v� ���~߾�������� �*�<�N�`�r����� ����������& 8J\n���� ������"4F Xj|����� ��//0/T/f/ x/�/�/�/�/�/�/�/ ??,?>?P?b?F/�? �?�?�?�?�?�?OO (O:OLO^OpO�Of?x? �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�O �O�_�_o o2oDoVo hozo�o�o�o�o�o�o �_�o.@Rdv �������� ��o<�N�`�r����� ����̏ޏ����&� 8�J�.�n��������� ȟڟ����"�4�F� X�j�|�`�����į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ�����Ŀ�� (�:�L�^�p߂ߔߦ� �������� ����6� H�Z�l�~������ ������� �2��(� h�z������������� ��
.@RdH� Z������� *<N`r�� z����//&/ 8/J/\/n/�/�/�/�/ �/��/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?�/O0OBOTOfO xO�O�O�O�O�O�O�O __,_OP_b_t_�_ �_�_�_�_�_�_oo (o:oLo^oB_�o�o�o �o�o�o�o $6 HZl~�to�� ���� �2�D�V� h�z��������� ��
��.�@�R�d�v� ��������П�Ə؏ �*�<�N�`�r����� ����̯ޯ����� 
�J�\�n��������� ȿڿ����"�4�F� *�T�|ώϠϲ����� ������0�B�T�f� x�\Ϝ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� �����2DV hz������ �
//./@/$d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?V/�? �?�?�?�?�?OO&O 8OJO\OnO�O�Ov?�? �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�O �O�_oo0oBoTofo xo�o�o�o�o�o�o�o �_,>Pbt� �������� (�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�