��   u��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����UI_CON�FIG_T  �� A$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�62�ODE�
3�CFOCA �4VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�;�  &USTOM~0 t $} RT_SPID�r,DC4D*PAG� �?^DEVIC�EPISCREuE�F��IGN�@$/FLAG�@C��1  h 	$P�WD_ACCES� E �8��C��!�%)$LABE�� $Tz jа@�3�B�	CUS�RVI 1  < `�B*�B��A7PRI�m� t1�RPTRIP�"m��$$CLA�@ O���sQ��R��RhP\ SI�qW�  �5�QIRTs1q_�P'�2 L3hL3!�pR	� ,��$?����R�P�S�S��Q@o�P� � o��
 ���)/SOFTP�.@/GEN�1?c�urrent=m�enupage,?1133,18o�o��o�o��Mo_o,13�88vo/A �'�o�n9�o�����ocmc480`|�%�7�I� �zQ a�s���������͏\� ���'�9�K�ڏo� ��������ɟX���� �#�5�G�Y��}��� ����ůׯf������1�C�U��� TPTX��y��|��o� s �o����$/soft�part/gen�link?hel�p=/md/tpia.dgd����"��4��r&ɿۻpwd 꿁ϓϥϷ������ ���#�5���Y�k�}� �ߡ߳�B�T�������1�C����zQ2'f	oC ($�ߕ����������i  zQ�Q�op��������SBg*��Q(a���*�����  1��P����@�R�n���)��#`  �V������SB� 1�XR �\ }%`wREG VED��� wholemod.htm4	�singlEd�oub\tr�iptbrows�@�!��� �/AS|��/Adev.s�Jl�o�1�	t���w�G/Y/ k/5/�/�/�/�/�/ ?� �P?*?<?N? `?r?�?�?�?�?�6�@ ?�?�?�? O2ODOE 	�/�/wO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_��_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-??z�� �����
��O @�R�!�3�����QOcO I�ݏ��*�%�7� I�r�m��������ǟ ٟ�����_/�)�W� i�{�������ïկ� ����/�A�S�e�w� ����iֿ����� 0�B�T�f�x�s��Ϯ� }Ϗ����ϭ�����>� 9�K�]߆߁ߓߥ��� ��������#�5�^� Y�k�9��������� ������1�C�U�g� y��������������� ſ2DVhz�� ������
�� @R	����� ����/*/%/7/ I/r/m//�/�/�/�/ ���/�/?!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSO!�O �O�O�O�O�O�O__ 0_+T_f_5_G_�_�_��Z�$UI_TO�PMENU 1��P�QR� 
d�QfA)�*default�qOZM*lev�el0 *\K	 #o� So�_Qo�cbtpio[23�]�(tpst[1�heo�ouo3oEo�-�
h58e01.�gif�(	me�nu5&ypHq13&zGr%zEt4M{4�a�������� �eB�C�U�g�y������,�prim=�Hqpage,1422,1��ݏ�� �%�0�I�[�m�������2���class,5������4)�4���130�f��x�������5���53ʏ���� �2�5���8ٯm������ ��4�ٿ����!�3�^I�P�Q�_k�m]�`�a[ϕ�ϝfty�m<�o�amf[0�o��}	��c[164�g.�59�h�a���k�Ax2uK}��azmWw %{�ߩsK�]�6�H�Z� l�~�ɿ��������� ��� �2�D�V�h�z�	���2���������� 	��ʟ?Qcu� (T�������Ѥ1$�N`r������ainedic����//��config�=single&>��wintpĀ / `/r/�/�/E�W��/{���gl[47��ow�H?���!8��� 6�i.?h?>82ڀ??�?��?z\rLz\r4s&x�? OVx`�6O� �O�O�O�O�O�O��O _#_5_G_Y_k_�O�_@�_�_�_�_�_,$;4$�doub?%o��1}3ؠ&duali38#�,4�_Pobo�_9o,n'o9ato�o �o�o}_,>Pb t������ �����o4�F�X�j�|� �����ď֏���=J�/,�wω¯���YOw���s�͔����ϡ�u��l�V�ȟ.��?RO�<��߬ߚ�6��u7 ��� �����/�A� ��e�w���������N� �����+�=�O�."$13�ϛϭϿ� ��ܿ����+�=�O� ��s߅ߗߩ߻����� "���'�9�K�]�����6d��������,$۬74��/�A��S�e�C����?�	�TPTX[209�,���2�(��������1I8��
����0P2���1_�1�Y�tv�������0�
�1�
ïqC:�4$treevie�wA#.f3�m381,26=o��� l����//+/� O/a/s/�/�/�/�_B�5$oq�?)?;? F/_?q?�?�?�?�?H? �?�?OO%O7O�/�/�1�/r2V��O�O��O �6XO�edit2azO�O_._@_ �?���OSL_�_�_ �_~��_�_G�o}o �CoUogoyo�o�o�o �o/o�o�o	-? Qduӥ���� ����?2�D�V�h� z������ԏ��� 
����@�R�d�v��� ��)���П����� ��<�N�`�r�����%� ��̯ޯ���&��� J�\�n�������3�ȿ ڿ����"��_�_X� o|��o��ϱ����� �����ߋ�)�S�e� x߉ߛ߭߿��ߓ� �,�>�P�b�t￿�� �����������(� :�L�^�p�������� ������ ��$6H Zl~���� ��� 2DVh z������ 
/�./@/R/d/v/�/ 7�IϾ/m��/I���? ?)?;?M?`?q?�?�/ �?�?�?�?�?OO%O 7O��nO�O�O�O�O�O �O%/�O_"_4_F_X_ �O|_�_�_�_�_�_e_ �_oo0oBoTofo�_ �o�o�o�o�o�oso ,>Pb�o�� �������(� :�L�^�p�������� ʏ܏/�/$��/H� �?MOk�}�������ş ؟�W����1�C�U� h�y�����_Oԯ��� 
��.�y�@�d�v��� ������M������ *�<�˿`�rτϖϨ� ��I�������&�8� J���n߀ߒߤ߶��� W������"�4�F��� X�|��������e� ����0�B�T����*defaul�ta�2�*level8����������{� tpst�[1]��ytpio[23��u�������	menu7.gkif�
�13�	B�5�
��
�4�u6�
ʯ?Qcu �������/ /�;/M/_/q/�/�/��/6"prim=��page,74,1�/�/�/??+?�6"�&class,130?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO~O`�O�O�O�/�"18�/��O__'_9_DON26�@_u_�_�_�_�_���$UI_USERVIEW 1���R 
���_>��_
o�m(oQocouo�o�o <o�o�o�o�o�o) ;M_qo~�� ����%��I� [�m������F�Ǐُ ������.�@��� {�������ßf���� ��/�ҟS�e�w������F�*zoom>��ZOOM��W� I��$�6�H�Z���~� ������ƿi������ �2�DϦ�maxr�esH�MAXRES߯E�㿬Ͼ��� ���ϗ��*�<�N�`� ߄ߖߨߺ���w��� ����o�%�J�\�n�� ��5����������� "�4�F�X�j��w��� ����������� BTfx��?� �����'= �t����_� �//(/�L/^/p/ �/�/?�/�/�/7/�/ ?$?6?H?Z?�/~?�? �?�?�?i?�?�?O O 2O�/?OUOcO�?�O�O �O�O�O�O
__._@_ R_d__�_�_�_�_�_ sQ