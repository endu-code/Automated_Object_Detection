��   u��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����UI_CON�FIG_T  �� A$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�62�ODE�
3�CFOCA �4VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�;�  &USTOM~0 t $} RT_SPID�r,DC4D*PAG� �?^DEVIC�EPISCREuE�F��IGN�@$/FLAG�@C��1  h 	$P�WD_ACCES� E �8��C��!�%)$LABE�� $Tz jа@�3�B�	CUS�RVI 1  < `�B*�B��A7PRI�m� t1�RPTRIP�"m��$$CLA�@ O���sQ��R��RhP\ SI�qW�  �5�QIRTs1q_�P'�2 L3hL3!�pR	� ,��d?����Q�P�R��T�Q�����P?�  �����
 ��)/SO�FTP.@/GEN��1?curren�t=menupa�ge,1133,18o�o�o�o��Mo_o,1388vo�/A �'�o�n9 �o�����ocmc480|�%�7�I� �zQa�s������� ��͏\����'�9� K�ڏo���������ɟ X�����#�5�G�Y� �}�������ůׯf������1�C�U���� TPTX���y�򨑿o� s� �o���$/s�oftpart/�genlink?�help=/mdw/tpia.dgd� ���"�4��r&ɿۻpwd꿁ϓϥϷ� ��������#�5��� Y�k�}ߏߡ߳�B�T߀������1�C�����zQ'f	bN� ($�ߕ���������i zQ�Q� c�Sj�n������A
)��Q(aa
a����  ��P����@��n���q��P#`  �V�p�����SB 1�X�R \ }|%`REG �VED�� w�holemod.�htm4	sing}lEdoub\�tript?brows�@� !����/�AS|�/Ad/ev.sJl�o�1�	t��� w�G/Y/k/5/�/�/p�/�/�/ ?� �P ?*?<?N?`?r?�?�? �?�?�6�@?�?�?�?  O2ODOE	�/�/wO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_��_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? ?z������ �
��O@�R�!�3� ����QOcOI�ݏ� �*�%�7�I�r�m�� ������ǟٟ���� �_/�)�W�i�{����� ��ïկ�����/� A�S�e�w�����iֿ �����0�B�T�f� x�s��Ϯ�}Ϗ����� ������>�9�K�]߆� �ߓߥ���������� �#�5�^�Y�k�9��� ������������� 1�C�U�g�y������� ��������ſ2DV hz������� �
��@R	�� ������� /*/%/7/I/r/m// �/�/�/�/���/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSO!�O�O�O�O�O �O�O__0_+T_f_�5_G_�_�_�Z�$U�I_TOPMEN�U 1�P�Q�R 
d��QfA)*def�aultqOZM�*level0 =*\K	 o� �So�_Qocbtpi�o[23]�(tpst[1�heo�o�uo3oEo�-
h58e01.gif~�(	menu5&ypHq13&zGr%zEt14M{4�a���� �����eB�C��U�g�y�����,�p�rim=Hqpag�e,1422,1 ��ݏ���%�0�I�@[�m������2���class,5��@����)�4���130�f�x�������5���53ʏ���P� �2�5���8ٯ m��������4�ٿ� ���!�3�^I�P�Q �_k�m]��a[ϕ��Ɲfty�m�o�amf�[0�o��	��c[g164�g.�59�h �a���k�Ax2uK} ��azmWw%{�ߩsK� ]�6�H�Z�l�~�ɿ�� ����������� �2�@D�V�h�z�	���2�� ��������	��ʟ? Qcu�(T��@�����Ѥ1$�@N`r�����?ainedic�����//�co�nfig=sin�gle&��wintpĀ /`/r/�/�/�E�W��/{���gl[�47��ow�?���!8���� 6�i.?h?>82 ڀ??�?�?z\rLz\r4s&x�? O Vx`�6O��O�O�O�O �O�O��O_#_5_G_ Y_k_�O�_�_�_�_�_��_,$;4$doub�?%o��13ؠ&d�uali38#�,!4�_Pobo�_9o,n 'o9ato�o�o�o}_ ,>Pbt�� ���������o4� F�X�j�|������ď֏���=J�/,�w�@�¯���YOw���s�������ϡ�u��l�V� ȟ.��?RO<��߬ߚ�6��u7��� ��� ��/�A���e�w��� ������N������P+�=�O�."$13 �ϛϭϿ���ܿ��� �+�=�O���s߅ߗ� �߻�����"���'� 9�K�]�����6d����������,$۬74���/�A�S�e�C�����?�	TPTX�[209�,���2 �(��������1I8��P
����0P2��`�1_�1�Y�tv�������0�
�1��
ïqC:4$tre�eviewA#.f3��m381,26 =o���l���� //+/�O/a/s/�/ �/�/�_B�5$oq �?)?;?F/_?q?�? �?�?�?H?�?�?OO %O7O�/�/�1�/r�2V��O�O�O �6<XO�edit2azO �O_._@_�?���O SL_�_�_�_~��_�_ G�o}o�CoUogo yo�o�o�o�o/o�o�o 	-?Qduӥ ��������? 2�D�V�h�z������ ԏ���
����@� R�d�v�����)���П �������<�N�`� r�����%���̯ޯ� ��&���J�\�n��� ����3�ȿڿ���� "��_�_X�o|��o� �ϱ����������� ��)�S�e�x߉ߛ߭� ���ߓ��,�>�P� b�t￿�������� ����(�:�L�^�p� �������������  ��$6HZl~ �������  2DVhz�� ����
/�./@/ R/d/v/�/7�IϾ/m� �/I���??)?;?M? `?q?�?�/�?�?�?�? �?OO%O7O��nO�O �O�O�O�O�O%/�O_ "_4_F_X_�O|_�_�_ �_�_�_e_�_oo0o BoTofo�_�o�o�o�o �o�oso,>P b�o������ ���(�:�L�^�p� �������ʏ܏/ �/$��/H��?MOk�}� ������ş؟�W��� �1�C�U�h�y����� _Oԯ���
��.�y� @�d�v���������M� �����*�<�˿`� rτϖϨϺ�I����� ��&�8�J���n߀� �ߤ߶���W������ "�4�F���X�|��� ������e�����0��B�T���*de�faulta�2�*level8����������{� tpst[1]���ytpioG[23��u������	men�u7.gif�
&�13�	�5�
�4�
�4�u6�
ʯ ?Qcu���� ���//�;/M/�_/q/�/�/�/6"p�rim=�pag?e,74,1�/�/��/??+?6"�&class,130?�f?x?�?�?�?=?O25��?�?�?O O2O5# D<�?lO~O�O�O�O�/�"18�/�O__'_9_DON26@_u_�_�_��_�_��$UI_�USERVIEW� 1���R 
�� �_>��_
o�m(oQo couo�o�o<o�o�o�o �o�o);M_q o~����� �%��I�[�m���� ��F�Ǐُ����� �.�@���{������� ßf������/�ҟ�S�e�w�����F�*�zoom��ZOOM��W�I��$�6� H�Z���~�������ƿ i����� �2�DϦ�maxresH�?MAXRES߯E� 㿬Ͼ������ϗ�� *�<�N�`�߄ߖߨ� ����w�������o�%� J�\�n���5���� �������"�4�F�X� j��w���������� ����BTfx ��?���� ��'=�t�� ��_��//(/ �L/^/p/�/�/?�/ �/�/7/�/?$?6?H? Z?�/~?�?�?�?�?i? �?�?O O2O�/?OUO cO�?�O�O�O�O�O�O 
__._@_R_d__�_ �_�_�_�_sQ