��   m�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING,��<$1_8k  �FMS*�t *v M_LIF��u,(8*x��M(DSTB0+_0>*_���*#�z&+CL_TIM>�PCCOMi��FBk M� �MAL_�EC�S��P!Q%XO �$PS� �TI����%�"r $D�TY?R. l*1E�ND14�$1�ACST1#4V22\93\9�4\95\96\6_O3VR\6� GA[7�2 h7�2u7�2�7�2�7�2ޜ8FRMZ\6DE��DX\6CURL� HSZ27Fh1DG u1DG�1DG�1DG�1DC�NA!1?( �sPL� + ���STA23TRQ_�M��/@K"�FSUX�JY�JZ�II�JuI�JI�D �$U1�SS  ����6Q����+PV�ERSI� 4W  �5GQ?IRTUAL3_EQ�' 1 TX W ��(P���_�_�_�Vm���څ �!� ���~����������R?����?��J�B�y4���=�t��7�Q��]�����V���u�������� � �^_P�dygwe�YAQ�o�^A����O ����a I ������o�o�_�l0/VSet�$�w�gAPB�w�un�Q�� Su����g`� ���`��	 j�����& ~�����j��b%��d�o#�5�G����=L��R�y�?�z���@�����я� ����+�=�O�a�s���� rU������ޟ:T  2��!� 3�E�W�i�{���������<��ۯ����#� 5�G�Y�k�}���������$$ 1�\��aP��J���`J}8*T[���P��$N��}�p�kD�EJ���:Ha�@��J`BB��@�G(�mA��\�1��\�mB�@k�B����`���C+���Pk��.dP�o�Ϙ�����+�=ϟ���M�x���2ߡ�V�A�z���� @P�� ��֠՞՞� ����{Ђ�K�}�gL��3L�X�������L��c�MZQ�M�ZR<MZS�MWZZ��3��8�H�L�VM]+NMoUq؉td ���t����פ�6Q�Q� ������8NS$T�i���i����/U �� ��� �x
� x��������NQ�U�Q�sQ�WQ�BM��C�T�C����C���������E����������������Ə���%����^��p���C��C�F��C�4�C����C������� ��6g�� �7� 4�7 m�t� �ZN �X�� �W �Ts� �1�5���&N� �s�W �/4� �4� �5�9�m9�������{��M��Q��� ��r��Na�,a�$a� �2��ړ����� ���vc+�{��M�U�M��M��M��M�I���ѡ�š����}� t��� 0q� 1�� 1�L 1ح��ρu��EA���@��s����������������}z��N����M��Ƞ7��9��O��K͋ w�3�W�n	 1	 i	 �� �Ġ��1�g���F Av_��q�����U#��+��&��8��'��>�HdUc

BeAIHJ��`�K��k}+����1"sP���xtesPe�E�Q���`EhsP�td��8�f������}� 2  ��B?S	-��sewasP�!?PO�sP������9��������l>�����ahi�A�s�sPE쩀>����� ������{� �©���H楄��s�sP�bsP�sP�zsP���(����������sPd��ͭM��>AQ���4-8���P�Ǡ_� =/��WSsP��эLiF.�'ce�+�/`,�/�$���� ??���*���I��ڭD�@�^��0g�0p�D���=�.�Ħ^��ħ��0��0��?�����&J���L��.c���/m�@�z��0��06�0G�0Pz�0Y�?�s��0��?�t_?�.�k����?-���?-��?-���?-�x?����@��?����?)�?�~��?���?�q}`!@�?�r")@��)@���z�w�9@��z����鬾�b?���>���I.���\ž�v�u��l��ſ���]�2����!�{.��z�ۮ�z�;y@��y@�9@��@?����@��BA�=���@K��@5��@D�@N=%���>y�">�w��ޠ�@Gh��@�@?�E�@ߪ�@ԍ@ʍ@�5Bh��b�hΪ�@���"�V��>�����,���m���;B���f���/?����?�׫�M�?�:E�i�_��hճ�h�9��h�W�hѻ�)Pm��B���B��9Q�ݫ��?�K��Jvh��Ju�MP}MP8�?����i���C͆?+���u�9P!5P
�5P5P 5P9P��� ,($not �a program|?���_�_�_�_�_PLACE�_%o�_Io0hZERXmoTo fo�o�o�o�o�o�o4dFRAM�o,7oP�7I�($A�q_?POSPIC���xA��_q�� ��#�`�G���k�}�𺏡�ޏ��PLCL�ų��� D1�ѐ?��  �>���?C��q�T�m�x� c�������������� ��>�P�