��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�0J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA!R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B!SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C?CFS_UT~p0 "�1�3�#�ؗ`qX"�}R0  4F OIMCM�`O#S�` ��upi �_�p��B}�a���M/� h�pIMPEE_F�N��N���@O��r�D_�~�n��Dy�F��K��_8�r0  T� '��'�DI�n0"���p�P�$Ix���� �CF�t7 X� GRP0�z�M=qNFLI�<7��0UIRE��$�g"� SWITCH^5�AX_N�PSs"�CF_LIM�� � �0EED��!��qP�t�`P�J_dVЦMODE�h�.Z`�PӺ�ELBOF� �������p� ���3���� F@B/��0�>�G�� �� WARN	M�`/��qP��n�wNST� COR-�0bFLTRh�T�RAT�PT1�� $ACC1a��N ��>r$ORI�o"6V�RT�P_S� WCHG�0I��rQT2��1�I��T��I1��� x �i#�Q��HDR�BJ; CQ�2L�3�L�4L�5L�6L�7�L� N�9s!gACO`S <F +�=��O��#92��LLEC�y�"MULTI��b�"N��1�!���0T��� �STY �"�R`�=l�)2`�p���*�`T  |�  �&$��۱m��P�Ḻ�UTO���E��EXT����ÁB���"2� (䈴![0������<�b+��� "D"���ŽQ���<煰kcl�9�# ���1��ÂM�ԽP���" '�3�$ L� E���P<��`=A�$JOBn�T����l�TRIG3�% dK�������<����\��+�Y�6�CO_yM��& t�p3FLܐBNG AgTBA� ���M��
 �!��p� �q��0�aP[`��O�'[����0tna*���"J���_R���CDJ���IdJk�D�%C��`�Z���0��P_��P��@ ( @F RaO.��&�t�IT�c�NOM�
���P�S���`T)w@����Z�P�d���RA��0��2b"����
$�T����MD3�TD��`U31���p(5!YHGb�T1�*E�7�c�KAb�WAb�cA�4#YNT���PD'BGD�� *(��PUt@X��W����AX��a��eTAI^cBUF��0!�+ � 7n�P�IW�*5 P�7M��8M�9
0�6F�7S�IMQS@>KEE�3PATn�^�a"� 2`#�"�L64F;IX!, ���!dĶ�D�2Bus=CCI��:FPCH�P:BAD�aHCEhAOGhA]H"W�_�0>�0_h@�f �Ak���F�q\'M`#��"�DE3�- l �p3G��@FSOES]FgHBSU�IBS9WC���. ` ��M�ARG쀳��FAyCLp�SLEWx�Qe�ӿ��MC�/�\pSM_JBM����QYC	g��e�q�Q�0 �n��CHN-�MP�G$G� Jg�_� <#��1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�fJR���rSEG�FR�PIO� S�TRT��N��cP!V5���!41�r�Ӏ
r>İ�b�B�O�2` +�[��� ,qE`&�,q`y�Ԣ}t8��yaSIZ%����t�vT�s� �z�y,qRSINF}Oбc����k��`��`�`Lp�ĸ T`7�CRCf�ԣCC/�9��`a�ua8h�ub'�MIN��uaPDs�#�G�D�YC��C�����e�q0��� ��EV�q�F�_
�eF��N3�s�ahƔ�Xa+p,5!�#=1�!VSCA?� �A��s1�"!3 ��`F/k��_�U��g�@�]��C�� a�s���}R�4� �ߠ��N����5a�R�HwANC��$LG��lP�f1$+@NDP�t�AR5@N^��a�q���c��ME�18����}0��RAө�AZ� 𨵰�%O��FCATK��s`"�S�P.FADIJ�OJ�ʠ �ʠ���<���Ր���GI�p�BMP��d�p�Dba��AESآ@	�K�W_��BA�S�� �G�5  �M�I�T�CSXh[@@�!62�	$X�K��T9�{sC���N�`�a~P_HEIsGHs1;�WID�06�aVT ACϰ��1A�Pl�<���EXqPg���|��CU�0_MMENU��7�TIT,AE�%�)�a2��a��8 YP� a�ED�E ��PDT��REM�.��AUTH_K�EY  ������ ��b�O	�0�}1E�RRLH� �9 \�� �q-�OR�DB�_�ID�@l �PUN_�O��Y�$SYSP0��4g�-�I�E��EV�#q'�PXW�O�� �: $SqK7!f2p�DBTd�wTRL��; �'�AC�`��ĠIND&9DJ.D��_��f1���f���PL�AF�RWAj���SD�A���!+r|��UMgMY9d�F�10d��&���J�<��}1PR�� 
3�POS���J�= �M$V$�q�PL~�!>���SܠK�?�����CJ�@����ENE�@T��A���S_��RECOR��B�H 5 O�@=$LA�>$~�r2�`R��`�q�b`�_Du�&�0RO�@�aT[�Q� �b������! }У��PAUS���dETgURN��MR�U�  CRp�EWyM�b�AGNAL:�s2$LA�!�?$PX�@$P��y A �Ax�C0 #ܠDO�`X�k��W�v�q�GO_AWAY��MO�ae����]�CSS_CCwSCB C �'N��CERI��гJ`u�QA0�}�\�@�GAG� R�0��`��{`��{`O�F�q�5��#M5A��X��&ш�LL�D� �$���sU�D)E%!`|���OVR10W��,�OR|�'�$E�SC_$`�eDSB#IOQ��l ��B.�VIB&� �c,������f�=pSSW����f!VL��PL|���ARMLO
���`����d7%SC� �bALspH�MPCh �Ch �#h �#
h 5�UU���C�'��C�'�#�$'�d�#C \4�$�pH��Ou��!Y��!�SB���` k$4�C�P3Wұ46�$VOLT37$$`�*�^1���$`O1*�$o��0R�QY��2b4�0DH_THE����0S�<�4�7ALPH�4�`����7�@ �0�qb7
�rR�5�88� ×@���"��Fn�	MӁVHBPFUAF�LQ"D�s�`�THR��i2dB�����G
(��PVP�����������1�J2�B�E�C�E�CPSu�Y@��F b3���H�(V�H:U�G��
X0��FkQw�[�N�a�'B���C INH=BcFILT��� $��W�2�T1�[ @��$���H YАAF�sDO��Y�R p� fg�Q�+�c5h`�Q�iSh�QPL��x�Wqi�QTMOU�# c�i�Q\��X�gmb��Hvi�h�bAi�fI�aCHIG��ca	xO��hܰ��W�"vAN-uX!��	#AV�H!Pa8$P�ד#p�RE_:�A�a��B�qN0�X�MCN�0��f1[1�qVE�p��Z2;&f�I�QO�u�r�x�wGldDN{G|d��aF>!�9��a9M:�U�FWA�:�Ml���X�Lu��$!����!l�ZO����0%�O�lF�s�13�DI�W�@��Q����_��!CURVAL԰0rCR41ͰZ�C <�r�H�v���<�`��<�(�f�CH�QR3��S���t���Xp�VS!_�`�ד�F��ژ����d?NS�TCY_ E 	L����1�t�1��U���24�2B�NI O�7������DEVIn|� F��$5�wRBTxSPIB�P���BYX����yT��HNDG��G H tn����L��Q�C���5�:�Lo0 H���閻�FBP�{tFE@{�5�t��T��I��DO���uPMCS��v>�f>�t�"HO�TSW�`s�ІE;LE��J T���e �2��25�� O� ��HA7�E��344�0>ܘ�A�K �� MD�L� 2J~PE ��	A��s��tːÈ�s�JÆG!��rD"��0������\�TO��W��	��/��SLAV��L  �0IN�Pڐ���`%ن_C�Fd�M� $n��ENU��OG��`b�ϑ]զP�0`�<��]�IDMA�Sa��\�WR�#��"]�sVE�$a�SKI�S!Ts��sk$��2u���J�������	��Q����_SVh�EXC�LUMqJ2M!ONLD��D�Y��|�PE �ղI_V�APPsLYZP��HID-@�Y�r�_M�2��VRFY�0��r�1�c�IOC_f�� 1�������O��u�LS����R$DUMMKY3�!���S� L_TP/Bv�"����AӞ�ّ N ����RT_u��� �G&r[�O �D��P_BA�`3�3x�!F ��	_5���H��N���� >�� P $�Kw�ARGI��� q��2O ��SGN�Z�Q �~P/�/PICGNs�l�$�^ �sQANNUN�@�T<�U/�ߴ�LAzp]	Z�d~��EFwPI�@ �R @�F?I�T�	$TOTA@%��d���!�mM�NIY�S+����E�A[�
DAYS\�ADx�@���	� �EFF_AXI?�TI��0z�COJA �AD�J_RTRQ��UBp��<P�1D �"r5̀Ll�T�0?  ]P�"p��mtpd��V 0w�G����Z����SK�SU� ���CTRL_C�A�� W�TR�ANS�6PIDLE_PW���!��A��V��V_�l�V �DIAGS�~��X� /$2�w_SE�#TAC����t!�!0z*@��R�R��vPA���p ; SW�!�!�  ��dol�U��oOH�f�PP� ��IR�r���BRK'#��"A_Ak���x 2x�9ϐ Zs2��%l�W�0t�*�x%RQDW�%MSx�t5AX�'�"��LIFECAL���10��N�1{"�5 Z�3{"dp5�ZU`}�/MOTN°Y$@�FLA�cZOVC�@p�5HE	��SU�PPOQ�ݑAq� L0j (C�1_X6�IEYRJZRJWRJ�0TH�!UC��6�XZ_A�R�p��Y2�HCO4Q��Sf6AN��w$��ICTE�Y� `��CACHE��C9�M�PLA�N��UFFIQ@��Ф0<�1	��6�
�N�MSW�EZ }8�KEYIM�p��TM~�SwQq��wQ#����OCVI�E� �[ A�B�GL��/�}�?� Q	�?��D\p�ذST��!�R� �T�� �T� �T	��PEM�AIf�ҁ��_/FAUL�]�Rц��1�U�� �T�RE�^< �$Rc�uS�% IT��BUFW}�Wr��N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTQT����sP��M��OtT�LwAX � ��X~`9#�c_G�3
N�YN_1�_�QD��1 �2M�U��T�F��H�@ g�`� p0p��Gb-sC_R�A�IK���r�t�RpoQ�u7h�qDSPq�2�rP��A�IM�c6�\����s2�U�@�A�sM*`IP���s�!DҐ6�TH�@n�)��OT�!6�HSDI3�ABSC���@ �Vy��� �_D^�CONVI�GÐ��@3�~`F�!�pd0��psqSCZ"����sMERk��qFB���k��pET���a6eRFU:@DUr`����x�CD,���@p�;cHR�A!��b`p�ՔՔ+PSԕ�C��C��p��ғSp�cH *�LX�:cd�Rqa� | ����W��U��U�@�U�	�U�OQU�7R��8R�9R��0T�^�1�k�1x�1��1��1���1��1��1ƪ2RԪ2^�k�2x�2��U2��2��2��2��U2ƪ3Ԫ3^�3k�Bx�3���o���3���3��3ƪ4Ԣ�AEsXTk!0�d <�  7h�p�6�pO��p�����NaFDRZ$eT^`V�Gr�����.�2REM� Fj��B�OVM��A�T7ROV�DT�`-�MX<�IN��0,�NW!INDKЗ
w�<׀�p$DG~q3�6��P�5�!D�6�R�IV���2�BGEA-R�IO�%K�¾DN�p��J�82�PB@>�CZ_MCM�@�1���@U��1�f ,<②a? ���P�I�!?I�E���Q����`m���g�� _0Pfqg RI�9ej�k!UP2_ gh � �cTD�p ���! a����bwBAC�ri T�Ph�b�`�) OG���%���p��IFI��!�pm�>��	�PT��"��MR2��j ��Ɛ+"�� ��\��������$�B`�x%��_ԡ�ޭ_����� M������D�GCLF�%DGDMY%LDa��5�6P�ߺ4@��Uk���? T�FS#p�Tl P���e�qP�p$EX_����1M2��2� 3�5���G ���m ���Ѝ�SW�eOe6D�EBUG���%G�R���pU�#BKUv_�O1'� �@PO�I5�5�MS��OOfswS�M��E�b���0�0_?E n �p� �TERM�}o� �ORI+���p�$Z �S�M_���b�q�T�A�r����UP�Rs� -��1�2n$�' o�$SEG,*> EL�TO��$USE.�pNFIAU"4��e1���#$p$UFR���0ؐO!�0����3OT�'�TAƀU��#NST�PATx��P�"PTHJ��©�E�P r�PV"AR�T�``%B`�abU!R�EL:�aSHFTp��V!�!�(_SH+@M$���� ��@N89r����OVRq��r�SHI%0��UN� �aAYLO����q�Il����!�@��@ERV]��1�?:�¦'��2��%��5�%�RyCq��EASYM�q��EV!WJi'��}�E ���!I�2��U@D� �q�%Ba��
5Po��0,�p6OR�MY� `GR��t2b5n�� � ��UPa�Uu �Ԭ")���TOCbO!S�1POP ��`�pC�������O,ѥ`REPR3��a�O�P�b�"ePR��%WU.X1��e$P�WR��IMIU�2R9_	S�$VIS��#�(AUD���Dv" �v��$H���P_�ADDR��H�G �"�Q�Q�QБR~pDp.1�w H� SZ�a���e�ex�e��S�E��r��HS��M�Nvx `���%Ŕ��OL���p<P��-��ACR�OlP_!QND_C���ג�1�T �ROUIPT��B_�VpQ�A1Q�v��c_��i�� �i��hx��i���i��6v�ACk�IOU���D�gfsu^d�y3 $|�P_D��V�B`bPRM_�b�]�ATTP_אH�az (��OBJ�Er��P��$��L�E�#�s`{ �s ��u�AB_x��T~�S�@�DBwGLV��KRL�Y�HITCOU�B�GY LO a�TEM��e�>�+P'�,P�SS|�P�JQUE�RY_FLA�b��HW��\!a|`�u@�PU�b�PIO ��"�]�ӂ/dԁ=dԁ~�� �IOLN���}����CXa$�SLZ�$INP7UT_g�$IP#�1P��'���SLvpa~��!�\�W�C-�CyX���pF_ASv��$L ��w �DF1G�U�B0m!���0HY��ڑ���$���UOPs� `������[�ʔ[�і"�[PP�SIP�<�і�I�2��IP_MEsMB��i`� X��cIP�P�b{�_N�`����R�����bSP��p$FO�CUSBG�a~�U=J�Ƃ �  � �o7JOG�'�DI�S[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A���APHIb�Qt�]�D� J7J\����� _KEYt�� �KՀLMO�Na���$XR���ɀ��WATCHa_��3���EL��b}Sy~���s� ���!V�g� �CTR�3򲓥��LG�D�� �R��I�
LG_SIZ���J�q XIƖ�I�FDT�IH� _�jV�GȴI�F�%S O���q �Ɩ���v������K�S����w�kR�N����E�@�\���'�*�U�s�5��@L>�4�DAUZ�EA�pՀ�Dp�f��GH�B,�OGB�OO��� C���PIT���� ���REC��SCRNě���D_p�b�aMARGf�`��:���TH�L���S�s��W�Ը��Iԭ�JGMO�MgNCH�c��FN���R�Kx�PRGv�UqF��p0��FWD��HL��STP��V`��+���Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*� a28����Gh�0CPO��������M8��Ģ��EX��TUIv�I��(�4� @�t�x�J0J�~�P���J0��N�a�#ANqA��O"�0VAIA���dCLEAR�6DCS_HI"�/cj�O�O�SI�r�S��IGN_��vpq�uᛀT�d� DEV-�LLA �°SBUW`��x0mT<$U�EM��PŁ�����A�R���x0�σ�a�@OS1�2�3�`�`� �ࠜh�AN%�-���-�IDX�DP��2MRO��Գ!�S�T��Rq�Y{b! _�$E&C+0��p.&A&T���`� L��ȟ%Pݘ��T\Q�UE�`�Ua~��_ � �@�(��`�b���# �M�B_PN@ R`r��<R�w�TRIN��P���BASS�a	6IkRQ6aMC(��� ��CLD�P�� ETRQLI`��!D�O9=4FLʡh2�Aq3zD�q7���LDq5[4q5ORG �)�2�8P�R��4�/c�4=b-4�t� ��rp[4*�L4q5S�@T�O0Qt�0*D2FRCLMC@D�?�?RIAtr,1ID`�D� d1���RQQprpDS3TB
`� �FᆻHAXD2���G�LE�XCES?R�q�BM�hPa�͠�BD4��E�q`�`�F_�A�J�C[�O�H� K���� \���bTf$�� ��LI�q�SRE�QUIRE�#MOx�\�a�XDEBU���E� L� M䵔 ��p���P�c�AA",1N��
Q�q�/�&����-cDC��B�IN�a?�RSM�Gh� �N#B��N�iPST�9� � 4��L�OC�RI���EX�fANG��A,1�ODAQ䵗�@1$��9�ZMF���� �f��"��%u#ЖV�SUP�%ؐ�FX�@IGGo�� �rq�"��1��#B��$���p%#by��rx��x�vbPDATAK��pE;���Z ��M܋�*� t�`MD
�qI��)�v� �t�A��wH�`��tDIA<E��sANSW��t(h���uD��)�bԣ�(@$`� PCU�_�V6�ʠ�d�PLODr�$`�R���B����B�p�����,1R�R2�E�  ���V�A/A d$OCALI�@��G~��2��!V��<$R�SW0^D"�kC�ABC�hD_J2�SE�Q�@�q_J3:M�
G�1SP�,��@PG�n�3m�u�3p
�@��JkC���2'A�O)IMk@{BCS�KP^:ܔ9�wܔJy�{BQܜ������`_AZ.B��?�E�L��YAOCMP0�c|A)��RT�j�ƚ�1�ﰈ��@1�茨����Z��SMG0��pԕ� ER!���*aINҠACk�p����b�n _�������D��/R��DIU��CD�H�@
�#a�q$�V�Fc�$x��$���`@���b���̂�E�H �$�BELP����!ACCEL���kA°�IRC_R�p�@��T!�$PS�@B2L`���W3��ط9� ٶPAT!H��.�γ.�3���p�A_��_�e�-B�`�C���_MG��$DD��ٰ��$FW�@�p����γ�����DE��PPAB�N�ROTSPE�Eu��O0��D�EF>Q��`$U�SE_��JPQPCD��JY����-A 6qYN�@A�L�̐�nL�MOU�NG���|�OL�y�INC U��a�¢ĻB��ӑ�AENCS���q�B��X���D�IN�I��0���pzC�VE�����23_U ��b�/LOWL���:�O0��0�Di�B�PҠȠ ��PRC����MOS� gTMOpp�@-GPERCH  M�OVӤ �����! 3�yD!e�]�6�<�� ʓA����LIʓdW�ɗ��:p3�.�I�TRKӥ�AY����?Q ^���m�b��`p�CQ�� MOM�B?R�0u��D���y�0Â擰DUҐZ�S_BCKLSH_C�� ��o�n��TӀ���x
c��CLALJ���A��/PKCHKtO0�Su�RTY� B�q��M�1�q_
#Nc�_UMCP�	C�΂�SCL���LMTj�_L�0X����E�� �� ����m�h���6��P	C����H� �P�Ş�CN@�"XT����C�N_��N^C�kCS	F����V6����ϡpj���nCAT�SHs�����ָ1����֙���������PAL���_P���_P0�� e���O1u�$xJaG� P{#�OG�>��TORQU(�p� a�~����Ry������"_W��^�����4t��
5z�
5I;I ;Iz�F�`�!��_8�1���VC��0�D�B�21��>	P�?�B�5JRK��<�2�6i�DBL_�SM�Q&BMD`_D9Lt�&BGRV4
D0t�
Dz��1H_���31�8JCOSEKr�EHLN�0hK�5oDt�jI���jI<1�J�LZ1�5Zc@y��1MYqA�HQB�THWMYTHET=09�NK23z�/Rln�r@CB4VCBn�CqPASfaYR<4gQt�gQ4VSBt��R?U'GTS���Cq��a���P#���Z�C$DUu ��R䂥э2�V�ӑ��Q�r�f$NE��+pIs@�|� �$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b�FP�c�j�FR�VrhVghTd��lV�jV�kV�kUV�kV�kV�kV�iHrh�f�r�m!�x�kUH�kH�kH�kH�kUH�iOclOrhO���nO�jO�kO�kO��kO�kO�kO�FF�.bTQ���E��egSPBALANCE���RLE�PH_'US�P衅F��F��FPFULC�3��3��E��1�l�UTOy_p �%T1T2t���2NW�����ǡ@��5�`�擳�T��OU���� INSE9G��R�REV��R����DIFH��1�l��F�1�;�OB��;C��2� �b�4?LCHWAR��i��ABW!��$ME�CH]Q�@k�q��AXk�P��IgU�i��� 
���!����ROB��CR��ͥ_T� �C��_s"�T � x ?$WEIGHh�9�#$cc�� Ih�.�sIF ќ�LAGK��8SK��K�BIL�?�OD��U��STŰ�P�; ����������
�Ы�Lў�  2�`�"�D�EBU.�L&�n���PMMY9��N8A#δ9�$D&����$��� Q ��DO_�A��� <	���~��L�IBX�P�N��+�_7��L�t�OH  �� %��T���Ѽ�T�����TICK,/�C�T1��%����B��N��c�Ã�R �L�S���S�����PR�OMPh�E� $IR� X�~ ���!�MAI�0��j���_9����t�l�R�0COD��F9U`�+�ID_" =������G_SUFF<0 3�O����DO��ِ��R� �Ǔن�S����!{���ꗰ�	�H)�_FIv��9��ORDX�3 ����36��4X�����GR9�S�n�ZDTD�\ t��ŧ4 *�L�_NA4���K��DEF_I[�K���g� ��_���i��Ɠ�š���IS`i �萚�D���e����4��0i�Dg����D�� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{ԓ�{� ��{����}��v�� ���g������^�� ��K�Փ����!w�N�P'���^���,`�W\�[R�7�T�EFĨ �O?ULOMB_u��0�VISPIT�Y�A�!OY�A_�FRId��(�SI���R������)3���W�W��0��0_,�EAS %��!�& "����4p�G;� h ���7ƵCOEFF_Om���m�/��G!%�S.�߲CA�5����u�GR` � � $R�4�� �X]�TME�$`R�s�Z�/,)�ER�qT;�:䗰�  ]��LL��S�_S�V�($~�����@���� "SwETU��MEA���Z�x0�u������ g� � �� ȰID�"���!*��&P���*�F�'�� ��)3��#���"��5;`*��RECt���!7�SK_���� P	�1_USER��,��4��8�D�0��VEL,2�0����2�5S�I�|���MTN�CFG}1�O  ���Oy�NORE��3��2�0SI���� ��\��UX-�ܑPDE��A $KEY�_����$JOG<EנSVIA�WC�� 1DSWy���
���CMULT�GI��@@C��2� 4� �#t�+�z�XYAZ��|�����z� �@o_ERR��� ��S L�-���@��s0�BB$BUF-@X�17ࡐMOR�� H	�CU�A3�z��1Q�
��3����$��FV��2�SbG�� � �$SI�@ G�0V�O B`נOBJE<&�!FADJU�#E�ELAY' ���SD�WOU�мE1PY���=0QT i�0�W�DIR$ba�8pےʠDYNբHeT�@��R�^�X�����OPWORK�}1�,�SYSsBU@p 1SOP�aHR�!�jU�k�PR��2�ePA�0�!�cu�V 1OP��UJ��a�'�D�QIMAGb�A	��`i�IMAC�rIN,�bsRGOVRD=a�b�0�aP�`sʠ� �^u�z�LP�B�@��!P�MC_E,�Q��N"@�M�rǱ��1Ų7�=qSL&�~0���$OVSL\G*E�D��*E2y�Ȑ�_=p �w��>p�s���s	�����y��t�#}1� �@�@;���O/�RI#A��
N��X�s�f�Rՠ���PL}1�,RyTv�m�ATUSRBTRC_T(qR��B �����$ �Ʊ��,�~0� D��`-CSALl`�SA���]1gqXE���%���bC��J�
���UP(4����PX��؆�q��y3�w� �PG�5�� $SU�B������t�JMPWAITO��s���LOyCFt�!D=�CCVF	ь�y���R`��0��CC_CTR��Q�	�IGNR_{PLt�DBTBm�P��z�BW)����0�U@���IG�a��I�y�TNLN��Z�R]aK� N��`B�0�P�E�s���r��f�SP]D}1� L	�A�`0gఠ�S��UN�{�传]�R!�`BDLY��2���7�PH�_PK�E��2RETRIEt��2�b5�����FI�B� �x���8� 2��0�DBGLV�LO�GSIZ$C�KT�ؑUy#u�D7�_�_YT1@�EM�@C\1�aA����R��D�FC�HECKK�R�P��0����@&�(bLYEc�" PA9�T����P�C߰PN�����ARh�0���Ӯ��PO�BORMATTnaF�f1h���2�S��UXy`	���LB��4�  ^rEITCH��W7��9PL)�AL_ �� $��XPB�q� C,2D�!��+2��J3D��� T�pPDCKyp��oC>� _ALPH����BEWQo���� ���I�wp � �~b@PAYLOA�Öm�_1t�2t���J3AR��؀դ֏�^laTIA4��5��6,2MOMCP������������0BϐAD���������PUBk`R��;���;��Ғ��z4�` I$PI\Ds�oӓ1yՕ�w�T2�w�Z��I��I��I���p����n���y�e`�9S)bT�S/PEED� G��(� Е��/���Е�`/��e�>��M��ЕSAMP�6V��/���Е#MO�@ 2@�A�� QP���C��n������� ����LRf`kb�ІE9h�EIN09��7 S.В9
yPy�/GAMM%S���D$GET)bP�ciD]��2
�IB�:q�I�G$HI(0;�A��LREXPA8)LWVM�8z)��g���C�5�CHKKp]�0�I_��h`eT��n� q��eT,����� �$�� �1�iPI� RCH�_D�313\��30L�E�1�1\�o(Y�7 ¾t�MSWFL �M.��SCRc�7�@�&���%n�f�SV���PB``�'�!�B�sS_SAV&0ct5B3NO]�C\�C2^� 0�mߗ�uٍa��u� ��u:e;��1���8��D�P��������� )��b9��e�GE��3��V�tQ��Ml��o � �YL��QNQSRlbfq XG�P�RR#dCQpH� �S:AW70�B�B�[�CgR:AMxP�KCAL�H���W�r�(1n�rg�M�!o�� �F�P@}t$WP�u�P  r��P5�R<�RC� R��%�6�`��� �Ôqsr X��OD�qZp�Ug�ڐ>D� ��OM#w�J?\?n?��?�?��9�b"�7�PuL]�_��� |� �X0��bf��qf��q`��ڏgzf��Eڐ� Q��Ce�"�ܰ�кFdPB��PM�Q}U�� � 8L��QCOU!5�QT�HI�HOQBpHY�SY�ES��qUE��`�"�O���  b�P�@\�UN��ʄCf�O�� �P��Vu��!����O�GRAƁcB2�O��tVuITe �q:pINFO�����{�q�cB�e�OI�r� =(�@SLEQS��q���p�vgqS����� 4L�ENAB|DRZ�PTIONt������Q���)�GCF:��G�$J�q^r�� R���U�8g�����_ED����'� �F��PK��5E'NU߇و�AUT$1܅COPAY�����n�00M�N���PRUTj8R �Nx�OU���$G[rf�@bRG�ADJ���*�X_:@բ$�����P��W��P��} ��)󂐶}�EX�YCDR[$~�NS.��F@�r�LGO�#�NY�Q_FREQR�W`� �#�h�TsLAe#�����ӄ �CRE�� s�IF��sNmA��%a�_Ge#STATUI`e#MAIL�����q �t�������ELE�M�� �/0<�FEASI?�B��n��ڢ�vA�]� � I �p��Y!q]�t#A��ABM���E�p<�VΡY�BASR�Z���S�UZ��0$�q���RMS_TR ;�qb ���SY�	�ǡ���$���>C�Q`	~� 2� _ �TM������̲�@ ��A��)ǅ�i$DOUd�s]$Nj���PR+@z3���rGRID�q�M�BARS �TY�@�|�OTO�p��� Hp_}�!����d��O�P/�� � �p�`POR�s��}�.��SRV��)����DI&0T����� �#�	�#�4!�5!�6J!�7!�8�e�F��2��Ep$VAL�Ut��%��ֱ��/��� ;�1�q��1���(_�AN�#��ⓡRɀ(���TOTcAL��S��PW��Il��REGEN�1�cX��ks(��a����`TR��R��_!S� ��1ଃV������⹂Z��`��E�Sp�3Vr���V_H���DA�S����S_Yh,1�R4�S� AR�P�2� ^�IG_CSE	s����å_Zp��C_�Ƃ�ENH�ANC�a� T� ;�������I#NT�.��@FPsİ/_OVRsP�`p� `��Lv��o��7�}�8�Z�@�SLG�AA�~�25�	��D��S�BĤDE�U������TE�P��ޏ� !Y��
�Jx��$2�IL_MC�0x r#_��`TQ�`�P�q���'�BV�C��P_� 0�M�	V�1�
V1�2�2��3�3�4�4 �
�!���� � m�Av�2IN~VIBPP���1�2�2�U3�3�4�4��A@-�C2���p�� MC_Fp+0��0L	11d���Mb50Id�%"E� S`��R/�@KEEP�_HNADD!!H`$^�j)C�Q���$��"	��#O�a_$A��!�0�#i��#REM�"�$��½%�!�(�U}�e�$HPWD�  `#SBM�SK|)G�qU2�:�P	�COLLAB� �!K5�B�� ��g��pITI1{9p�#>D� ,�@FL|AP��$SYN ��<M�`C6���U_P_DLYAA�Er�DELA�0ᐢY��`AD�Q��Q�SKIP=E� �4��XpOfPNTv�A�0P_Xp�rG�p�R U@,G��:I+�:IB1:I G�9JT�9Ja�9Jn�9Jt{�9J9<��RA=s� X���4�%1��QB� NFLIC��s�@J�U�H�LwN�O_H�0�"?��RIuTg��@_PA�p=G�Q� ��^��U��W��LV�d�NGRLT�0_q��O��  " ��OS��T_J�vA V	�APPR_�WEIGH�sJ43CH?pvTOR��vT��LOO��]�+�tVJ�е�ғA�Q�U�S��XOB'�'�@aJ2TP���7�X�T� <a43DP=`Ԡ\"<a�q�\!��RDC��L�+ �рR��R�`� ��RV��jr�b�R�GE��*��cN�FL�G�a�Z���SPC��s�UM_<`^2�TH2NH��P.a �1� m`EFv11��� lQ `�!#� <�p3AT�  g�S�&�Vr�p�tMq�Lr���HOMEVwr u2'r�-@?Qcu��w3'r�������w4'r�'�9�K�]�o����w5'r뤏��ȏPڏ����w6'r�!�@3�E�W�i�{��w7'r힟��ԟ����w8'r��-�?�Q�c��u��uS$0�q�p �� sF��`S0p� `P�����`/���&-�IO[M�I֠����1R�pWE��# ��0Za*���� �5��$DS=B GNAL���0�Cp��m`S232N3�� �~`��� �/ ICEQP��PE�p��5PIT����O�PBx0��FLOW�@TRvP��!U����CU�M��UXT��A��w�ERFAC��� U��ȳC�H��� tQ  _���>�Q$����O)M��A�`T�P#�UPD7 A�ct�T��UEX@�ȟ�U �EFA: X"�1RS9PT�����T ���PPA�0o񩩕`EXP�IOS���)Ԃ��_���%��C�WR�A��ѩD�ag֕`~ԦFRIENDsa�C2UF7P����TO;OL��MYH C2�LENGTH_V�TE��I��Ӆ�$SE����UFI�NV_���RsGI�{QITI5Bb��Xv��-�G2-�G17�w�SG�X��_��UQQD=#���AS��d~C�`��qᾭ� �$$C/�S�`�����S0�0|����VERSI� ����0�5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����S0����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT&�����  ��DINp�O�A�Dq�EXE�HiPV_��ATQ�z
��LARMRECOV ��RgLMDG �*�5�OLM_�IF *��`d �O�_�_�_�_j�_'o�9oKo]onm, 
 ��odb��o�o�o�o�^��$� z, A�   2D{�PPINFO u[ �Vw��������`������ �*��&�`�J���n�����DQ����
� �.�@�R�d�v����������a
PPLIC�AT��?�P���`Han�dlingToo�l 
� 
V8.30P/40Cp�ɔ_LI
88�3��ɕ$ME�
F0G�4�-

398�ɘ��%�z�
7D�C3�ɜ
�Non�eɘVr���ɞ@/6d� Vq?_ACTIVU�r�C죴�MODP����C�I��HGAP�ON���OU�P�1*��  i�m����Қ_�����1*�  �@��������Q����Կ�@�
������ ���5��Hʵl�K�HTTHKY_��/�M�S� ����������%�7� ��[�m�ߝߣߵ��� �������!�3��W� i�{���������� ����/���S�e�w� �������������� +�Oas�� �����' �K]o���� ����/#/}/G/ Y/k/�/�/�/�/�/�/ �/�/??y?C?U?g? �?�?�?�?�?�?�?�? 	OOuO?OQOcO�O�O �O�O�O�O�O�O__ q_;_M___}_�_�_�_`�_�_�_kŭ�TOp���
�DO_CLE�AN9��pcNM  !{衮o�o�o��o�o��DSPDgRYRwo��HI��m@�or���� �����&�8�J���MAXݐWdak�H�h�XWd�d���PLUGGW�Xgd���PRC)pB�`"�kaS�Oǂ2^DtSEGF0�K�  �+��o�or�������8���%�LAPOb� x�� �2�D�V�h�z��������¯ԯ�+�T�OTAL����+�U�SENUO�\� �e�A�k­�RGDI_SPMMC.����C6�z�@@Dr\�O�Mpo�:�X�_STRING 1	(��
�M!�S��
��_ITE;M1Ƕ  n�� ����+�=�O�a�s� �ϗϩϻ����������'�9�I/O SIGNAL���Tryout� ModeȵI�npy�Simul�ateḏOu�t��OVER�RLp = 100�˲In cyc�l�̱Prog� Abor��̱~u�Statusʳ�	Heartbe�atƷMH F�aul	��Aler�L�:�L�^�p�����������  ScûSaտ��-�?�Q� c�u������������� ��);M_q��WOR.�û�� ����+= Oas��������//'.PO ����M �6/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�?�?H"DEVP.�0d/ �?O*O<ONO`OrO�O �O�O�O�O�O�O__�&_8_J_\_n_PALT	��Q�o_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o�_GRIm�û9q �_as���� �����'�9�K��]�o�������'�R 	�݁Q����)�;� M�_�q���������˟ ݟ���%�7�I�ˏPREG�^����[� ����ͯ߯���'� 9�K�]�o����������ɿۿ�O��$AR�G_� D ?	����0���  	$�O�	[D�]D���O�e�#�SBN_C�ONFIG 
�0˃���}�CI�I_SAVE  �O�����#�TC�ELLSETUP� 0�%  O�ME_IOO�O�%?MOV_H���ώ��REP��J��U�TOBACK�����FRA;:\o� Q�o����'`��o���{� �� f� o�����*�!�3�`�����f������ ����o�{��&�8�J� \�n������������ ������"4FXj |������\끁  ��_i��_\ATBCKC�TL.TMP 6�.VD GIF PHD_q���N�t#��f�IN�I�P�Օ�c�MESSAG�����|8��ODE_D�����z��O�0�c�P�AUSM!!�0� (73�U/g+(Od/�/x/�/�/ �/�/�/�/???P?�>?t?1�0$: TSK�  @-��T�f�UgPDT��d�0�
&XWZD_ENqB����6STA��0��5"�XIS��U�NT 20Ž�� � 	 ���z��e�ng�-�?���S�o�U@��H����zF�OTo�}Cw�g�^�	���.�O�O�O�O�/_2FMET߀2�CMPTAA��@��$A-�@����@���@����]5���5�(d5��P�5�r�5F*�5�338]SCR�DCFG 1�6/�Ь�Ź�_�_oo(o:oLo��o�Q���_�o�o�o �o�o�o]o�o>P bt���o9�iуGR<@M/�s/N5A�/�	i��v�_ED�1�Y� 
 �%-5�EDT-�'�G?ETDATAU�o��9��?�j�H�o��f�\��A��  ���2�&�!�E���:IB���~�ŏ׏m����3��&۔� �D��ߟJ�����9�ǟ�4���ϯ�(�����]�o�����5 N������(�w��)�;�ѿ_��6ϊ�g� ��(�CϮ���ϝ�+��7��V�3�z�(��@z�����i����8��&���~�]���F����5����9~������]����Y�k�����CR�!ߖ��� W�q���#�5���Y��p~$�NO_DEL���rGE_UNUS�E��tIGALL_OW 1���(*SYST�EM*S	$S?ERV_GR�Vܖ : REG�$8�\� NUM�
���PMUB U�LAYNP\?PMPAL��CYC10#6x $\ULSU0�8:!�Lr��BOXORI�C�UR_��PM�CNV�1�0L�T4DLI�0��	����BN/ `/r/�/�/�/�/�/����pLAL_OUT� �;���qWD_ABOR=f�q�;0ITR_RTN��7�o	;0NONS�0�6 
HCCF�S_UTIL 9#<�5CC_@6Aw 2#; h ?��?�?O#O6]CE_�OPTIOc8�qF@RIA_I�c f5Y@�2�0FF�Q�=2q&}�Ao_LIM�2.�� ��P�]B�T�KX�P
�P�2O��Q��B�r�qF�PQ5T1)TR�H��_:JF_PARAMGP 1�<g^&S�_�_�_�_~�VC�  C�dE�`�o!o`�`U�`�`�Cd��T@ii:a:e>eBa�Gg�C�`� D� kD	�`�w?��2{HE ONFI� �E?�aG_P�1#; ���o�1CUgy�aKoPAUS�1�yC ,����� ����	�C�-�g� Q�w���������я���rO�A�O�H��LLECT_�B�IPV6�EN. QF�n3�NDE>� �G��71234?567890��sB�TR����%
 H�/%)������� W���0�B���f�x��� 㯮���ү+����� s�>�P�b��������� �ο��K��(�:�Г�^�|��B!F� ��I|�IO #��<U%e6�'�9�lK���TR�P2$���(9X�t�Y޼`%��̓ڥH��_MOR֮3&�=��@XB��a��A�$� �H�6�l�~���~S��'�=�r_A?�a�a`D��@K��R�dP��y)F�ha�-�_�'�9�%
�k��G�� ��%Z�%���`�@c.�PDB�+���cpmidbg��	�`:�����p��N  ��@��.����]ܭ@�s<�^��@bsg�$� s�fl�q��u�d1:��:J��D�EF *ۈ��)��c�buf.�txt����_�L64FIX ,������l/[Y/�/ }/�/�/�/�/
?�/.? @??d?v?U?�?�?�?��?�?�?,/>#_E -���<2ODOVO�hOzO�O6&IM��.zo�YU>���d�l
�IMC��2/��b��dU�C��20�M�QT:Uw�Cz  �B�i�A���A����Au�gB�3�*CG�B�<�=w�i�B.���B���B���5B�$�D��%B���ezVC��q�C�v�D����D-lE\D�n�j��ؤB9"��22o�DT|����� ����C�C����2
�xObi�D4cdv`�D��`/�`v`s]E��D D�` E�4�F*� E�c��FC��u[F����E��fE���fFކ3FY�F�P3�Z���@�33 ;���>L���Aw�n�,a@��@e�5Y����a���`A��w�=�`<#�*
��?�o�zJRSMOFS�T (�,bIT�1��D @3��
д��'�a��;��b�w?���<�{M�NTEST�)1O�CR@�4��>VC5`A�w�Ia+a��aORI`CTPB�fU�C�`4���rN��:d�*�qI?��5��qT_�P�ROG ��
�%�$/ˏ�t��NUSER  �U�������KEY_TBL � ����#a��	
��� !"#�$%&'()*+�,-./��:;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������������������������������������������������������������������������L�CK�
����ST�AT/��s_AUT_O_DO �	��c�INDT_EN�BP���Rpqn�`�T92����STOr`��v�XC�� 26��) 8
SONY? XC-56�"b�����@��F( �А�HRC50w���>�P�7b�t�Aff����ֿ� Ŀ����C�U� 0�yϋ�fϯ��Ϝ���������-ߜ�TRLޡ�LETEͦ ���T_SCREE�N ��k�cs���U�MM�ENU 17�� <ܹ���w��� ������K�"�4� ��X�j�������� ����5���k�B�T� z������������� ��.g>P�t ������ Q(:�^p�� ��/��;//$/ J/�/Z/l/�/�/�/�/ �/�/�/7?? ?m?D? V?�?z?�?�?�?�?�? !O�?
OWO.O@OfO�O�vO�O�O(y��REG� 8�y����`��M�ߎ�_MANU�AL�k�DBCOΊ�RIGY�9�DB�G_ERRL��	9�ۉq��_�_�_� ^QNUMLIT�pϡ�pd
�
^Q�PXWORK 1:���_5oGoYoko|}oӍDBTB_Nѧ ;������ADB_AW�AYfS�qGCP� 
�=�p�f_AL�pR��bbRY�[�
��WX_�P 1<{y�n�,�%oc�P�6�h_M��ISO��k�@L��sONTIM6X��
���vy�
��2sMOTNE�ND�1tRECO�RD 1B�� y���sG�O�]� K��{�b��������V� Ǐ�]����6�H�Z� ��������#�؟� �����2���V�şz� �������ԯC���g� �.�@�R���v�寚� 	���п���c�χ� #ϫ�`�rτϖ�Ϻ� )ϳ�M���&�8ߧ� \�G�Uߒ�߶�����@I������4�� �p 7�n���ߤ����� �����"���F�1��� |��������[����� i���BTf����bTOLEREN�C�dB�'r�`L���^PCSS_CC?SCB 3C>y�`	IP�t}�~� <�_`r�K�@����/�{�� 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�OX_�~�LL� D���&qET�c�a 7C[C��PZP\^r_ A� p� ��sp��QGPt[	� A�p�Q�_�[?� �_�[oU�p1�P�pSB�V�c �(a�PWoio{h+�o��X�o�oY��[	r�hLW���N:p�����}6ګ��c��aD@�VB��|�G����+��K� �otGhXGr��So����eB   =��Ͷa�>�tYB�� �pC(�p�q�aA"�H�S�Q -��q���ud�v���|��AfP ` 0����D^P��p@�a
�QXTHQ�$���a aW>� �a9P��b�e:�L�^�h�Hc�́PQ�RFQ� PU�z�֟�o\^�� -�?��c�u����zKCz�ů�b2᤼Щ�RD�����l)*����S̡0��]��0�.��@���EQ� �p��F�X�ѿUҁп��VSȺNSTCOY 1E��]�ڿ��K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߒ���DEVICE 1F5� MZ�۶a ��	� ��?�6�c����	{䰟���_HN?DGD G5�VP����R�LS 2H �ݠ��/�A�S�e�w������ ZPARAMG I�FgHe��RBT 2K���8р<��WPpC�*C��,`¢P�Z�z���%{�C�� 2�jMTLU,`"nPB, s��M� `}�gT�g��
B��!�bcy�[2D chz����/���/gT#I%D��C�` b!�R���A��A,�ͿBd��A��P���_C4kP�!2�C���$Ɓ�]�ffA��À��B�� ��| ���/�/�T ( ��54a5�}%/7/ d?/M?_?q?�?�?�? �?�?O�?OO%O7O IO�OmOO�O�O�O�O �O�O�OJ_!_3_�_�_ 3�_�_�_�_�_o�_ (ooLo^oЁ=?k_Io S_�o�o�o�o�o�o �o#5G�k} �������H� �1�~�U�g�y�ƏAo �Տ���2�D�/�h� S���go����ԟ���� ϟ���R�)�;��� _�q����������ݯ �<��%�7�I�[�m� ��������}�&�� J�5�n�YϒϤϏ��� ��ѿ������F�� /�Aߎ�e�w��ߛ߭� ��������B��+�x� O�a��������� ��,���%�b�M���q� ������������� �L#5�Yk} ��� ��6 1CUg��� �����	//h/ ���/w/�/�/�/�/�/ 
?�/.?@?I/[/1/ _?q?�?�?�?�?�?�? �?OO%OrOIO[O�O O�O�O�O�O�O&_�O _\_3_E_W_�_?�_ �_�_�_�_"ooFo1o joE?s_�_�om_�o�o �o�o�o0f= Oa������ ����b�9�K��� o���Ώ��[o��(� �L�7�I���m�������$DCSS_S�LAVE L����ё���_4D  �љ��CFG MMѕ��������FRA:\�ĐL-�%04d.wCSV��  }��� ���A i�CH
q�z������|���.��  �����Ρ�ޯ̩ˡҐ-��*�����_CRC_O_UT N�������_FSI ?}њ �� ��k�}�������ſ׿  �����H�C�U�g� �ϋϝϯ���������  ��-�?�h�c�u߇� �߽߫��������� @�;�M�_����� ����������%�7� `�[�m���������� ������83EW �{������ /XSew �������/ 0/+/=/O/x/s/�/�/ �/�/�/�/???'? P?K?]?o?�?�?�?�? �?�?�?�?(O#O5OGO pOkO}O�O�O�O�O�O  _�O__H_C_U_g_ �_�_�_�_�_�_�_�_  oo-o?ohocouo�o �o�o�o�o�o�o @;M_���� ������%�7� `�[�m��������Ǐ ������8�3�E�W� ��{�����ȟß՟� ���/�X�S�e�w� ������������� 0�+�=�O�x�s����� ����Ϳ߿���'� P�K�]�oϘϓϥϷ� ��������(�#�5�G� p�k�}ߏ߸߳�����  �����H�C�U�g� �������������  ��-�?�h�c�u��� ������������ @;M_���� ����%7 `[m���� ���/8/3/E/W/ �/{/�/�/�/�/�/�/ ???/?X?S?e?w? �?�?�?�?�?�?�?O 0O+O=OOOxOsO�O�O��O�O�C�$DCS�_C_FSO ?�����A P �O �O_?_:_L_^_�_�_ �_�_�_�_�_�_oo $o6o_oZolo~o�o�o �o�o�o�o�o72 DVz���� ���
��.�W�R� d�v����������� ��/�*�<�N�w�r� ��������̟ޟ�� �&�O�J�\�n����� ����߯گ���'�"� 4�F�o�j�|������� Ŀֿ������G�B�|T��OC_RPI�N_jϳ����ς��O�����1�Z�U��NSL��@&�h߱������� ��"��/�A�j�e�w� ������������ �B�=�O�a������� ����������' 9b]o���� ����:5G Y�}����� �///1/Z/U/g/ y/�/�/�/�/�/�/�/ 	?2?-???Q?z?u?�� ߤ߆?�?�?�?OO @O;OMO_O�O�O�O�O �O�O�O�O__%_7_ `_[_m__�_�_�_�_ �_�_�_o8o3oEoWo �o{o�o�o�o�o�o�o /XSew �������� 0�+�=�O�x�s����� ����͏ߏ���'��P�K�]�o����� �P�RE_CHK �P۪�A ��,8�2���� 	 8�9�K���+�q���a������� ݯ�ͯ�%��I�[� 9����o���ǿ��׿ ���)�3�E��i�{� YϟϱϏ�������� ���-�S�1�c߉�g� y߿��߯����!�+� =���a�s�Q���� �����������K� ]�;�����q������� ������#5�Ak {����� �CU3y� i������/ -/G/c/u/S/�/�/ �/�/�/�/??�/;? M?+?q?�?a?�?�?�? �?�?�?�?%O?/Q/[O mOO�O�O�O�O�O�O �O_�O3_E_#_U_{_ Y_�_�_�_�_�_�_�_ o/ooSoeoGO�o�o =o�o�o�o�o�o =-s�c�� �����'��K� ]�woi���5���ɏ�� ������5�G�%�k� }�[�������ן�ǟ ����C�U�o�A��� ��{���ӯ����	�� -�?��c�u�S����� ��Ͽ῿�����'� M�+�=σϕ�w����� m������%�7��[� m�K�}ߣ߁߳��߷� ���!���E�W�5�{� ��ϱ���e������� 	�/��?�e�C�U��� ������������ =O-s���� ]����'9 ]oM����� ��/�5/G/%/k/ }/[/�/�/��/�/�/ �/?1??U?g?E?�? �?{?�?�?�?�?	O�? O?OOOOuOSOeO�O �O�/�O�O�O_)__ M___=_�_�_s_�_�_ �_�_o�_�_7oIo'o moo]o�o�o�O�o�o �o!�o1W5g �k}����� �/�A��e�w�U��� ����я��o���� 	�O�a�?�����u��� ͟�����'�9�� ]�o�M���������ۯ ��ǯ�#�ůG�Y�7� }���m���ſ����� ٿ�1��A�g�E�w� ��{ύ�������	�� ��?�Q�/�u߇�e߫� �ߛ��������)�� �_�q�O������ �������7�I��� Y��]����������� ����!3WiG ��}���� %�A�1w�g ������/+/ 	/O/a/?/�/�/u/�/ �/�/�/?�/9?K? �/o?�?_?�?�?�?�? �?�?O#OOGOYO7O iO�OmO�O�O�O�O�O _�O1_C_%?g_y__ �_�_�_�_�_�_�_o �_+oQo/oAo�o�owo �o�o�o�o�o); U__q���� ����%��I�[� 9����o���Ǐ��� ��ۏ!�3�M?�i�� Y�������՟�ş� ���A�S�1�w���g� ���������ӯ�+��=��$DCS_S_GN QK�c���7m� 0�9-MAY-19� 14:33  � O�14-J�ANt�08:38�}����� N.DѤ����������h�x,rWf*�σ�^M��  �O�VERSION� [�V3�.5.13�EF�LOGIC 1R�K��  	���P�?�P��N�!�PROG_E_NB  ��6����o�ULSE  �TŇ�!�_AC�CLIM�����Ö��WRSTgJNT��c��K�EMOx̘��� ���INIT S.��G�Z���OPT_S�L ?	,��
 	R575��VY�74^�6_�7_�+50��1��2_�@�����<�TO  �Hݷ���V�DE�X��dc����P�ATH A[�A�\�g�y��HC�P_CLNTID� ?��6� �@ȸ����IAG_�GRP 2XK�� , `���� �9�$�]�H������1234?567890����S�� |�������8!�� ��H؀��;�dC�S��� 6�����. �Rv�f�� H��//�</N/ �"/p/�/t/�/�/V/ h/�/?&??J?\?�/ l?B?�?�?�?�?�?v? O�?4OFO$OjO|OO E��Oy��O�O_�O 2_��_T_y_d_�_,
�B^ 4�_�_~_ `Oo�O&oLo^oI��T jo�o.o�o�o�o�o  �O'�_K6H�l �������#� �G�2�k�V���B]� ��Ǐُ�������(���L�B\Drx�@���PC�����4  79֐�$��>���:������ߟʟܟ���CT_�CONFIG �Y��Ӛ��egU���STBF/_TTS��
��b�����Û�u�O�MA�U��|��MSW_�CF6�Z��  ~�OCVIEW��3[ɭ������ -�?�Q�c�u�G�	��� ��¿Կ������.� @�R�d�v�ϚϬϾ� ������ߕ�*�<�N� `�r߄�ߨߺ����� ����&�8�J�\�n� ���!���������� ���4�F�X�j�|�����RC£\�e��! *�B^������C�2g{�SBL_FAULT ]��|ި�GPMSKk���*�TDIAG �^:�աI���UD1: 67�89012345�G�BSP�-? Qcu����� ��//)/;/M/� �
@q��/>$�TRECP��

��/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOi/�{/xO�/UMP_OPTIONk���A�TR¢l��	�EP�MEj��OY_TE�MP  È�g3B�J�P�AP�DUNI��m�Q���YN_BRK �_ɩ�EMGDI_STA"U�aQSU�NC_S1`ɫ ��FO�_�_�^
�^d pOoo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{�E �����y�Q�� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d��z����� ��˟����%�7� I�[�m��������ǯ ٯ����!�3�E�W� i���������ÿݟ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�{�iߗ� �߻�տ������'� 9�K�]�o����� ���������#�5�G� Y�s߅ߏ�����i��� ����1CUg y������� 	-?Qk�}�� �������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?u?�?�?�?� �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_m?w_ �_�_�_�?�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9Ke_W����_ �_����#�5�G� Y�k�}�������ŏ׏ �����1�C�]o y��������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;���g�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�_� i�{ߍߟ߹������� ����/�A�S�e�w� ������������ �+�=�W�E�s����� �ߧ�������' 9K]o���� ����#5O� a�k}�E���� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-?GYc?u?�? �?��?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ Q?[_m__�_�?�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/I_Sew ��_������ �+�=�O�a�s����� ����͏ߏ���'� A3�]�o������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����9�K�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� ��C�M�_�q߃ߝ��� ����������%�7� I�[�m������� �������!�;�E�W� i�{��ߟ��������� ��/ASew ������� 3�!Oas��� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?+=G? Y?k?!?��?�?�?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O 	_#?5??_Q_c_u_�? �_�_�_�_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o-_7 I[m�_���� ����!�3�E�W� i�{�������ÏՏ� ���%/�A�S�e� q�������џ���� �+�=�O�a�s����� ����ͯ߯���� 9�K�]�w��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� �����'�1�C�U�g� ���ߝ߯��������� 	��-�?�Q�c�u�� ����������m�� )�;�M�_�y߃����� ��������%7 I[m���� ����!3EW q�{������ �////A/S/e/w/ �/�/�/�/�/�/�/ �/+?=?O?i_?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O��O�O�O? �$E�NETMODE �1aj5��  00�54_F[PRROR�_PROG %�#Z%6�_�YdUTA�BLE  #[�t?�_�_�_gdRSE�V_NUM 2R?  �-Q)`�dQ_AUTO_ENB  PU+SaTw_NO>a b#[�EQ(b  *�*�`��`��`��`4`�+�`�o�o�oZdHI�S%c1+PSk_AL�M 1c#[ �24�l0+�o;@M_q���o_b.``  #[aFR��zPTCP_VE/R !#Z!�_��$EXTLOG_7REQ�f�Qi,��SIZ5�'�STK�R�oe�)�TOoL  1Dz�b��A '�_BW�D�p��Hf��D�_D�I�� dj5�SdDT1KRņSTE�Pя�P��OP_�DOt�QFACTORY_TUN�g�d<�DR_GRP� 1e#YNad 	����FP��x�̹ ���� �$�f�?�� ��� ǖ��ٟ�ԟ���1� �U�@�y�d�v������ӯ����LW
 JG��>�,��tۯ��j�U���y�B� � B୰���$ � A@��s�@UU�UӾ�������E��� E�`F@ �F�5U/�,��L����M��J�k�Lzp�JP��Fg�f��?�  s��9��Y9}�9���8j
�6̿�6�;���A���O ���� � I� ������[F�EATURE �fj5��JQ�Handling�Tool � "�
PEng�lish Dictionary��def.4Dw St�ard��  
! h�Analog I�/OI�  !
�IX�gle Sh�iftI�d�X�u�to Softw�are Update  rt s����matic B�ackup�3\�st��gro�und Edit���fd
�Camera`�F�d�e��CnrRn�dIm���3�C�ommon ca�lib UI�� /Ethe�n��"�Monitor�oLOAD8�tr�?Reliaby�O��ENS�Data ?Acquis>���m.fdp�iag�nos��]�i�Do�cument V�ieweJ��87�0p�ual C�heck Saf7ety*� cy� ��hanced U�s��Fr����C� �xt. DIOm :�fi�� m8����end��Err�I�L��S������s�  t Pa�r�[�� ���J94�4FCTN /Menu��ve�M�� J9l�TP I�nT�fac{�  �744��G��p �Mask Excz��g�� R85��T��Proxy �Sv��  15 �J�igh-Sp�e��Ski
� R�738Г��mm�unic��ons��S R7��ur8r�T�d�022��a����connect� 2� J5��I�ncr��stru�,Қ�2 RK�AREL Cmd�. L��ua��R�860hRun-�Ti��EnvL�o�a��KU�el +:��s��S/Wѹ��7�License����rodu� o�gBook(Sy�stem)�AD� pMACR�Os,��/Off�s��2�NDs�MH��� ����MM�RC�?��ORDE�� echStopr��t? � 84fcMi$�|� 13d�x��]е�׏���M�odz�witchBI�VP��?��.� sv��2Opt�m�8�2��filз�I ��2g 4� !+ulti-�T�����;�P?CM funY��Po|���4$�b&R�egi� r �P�ri��FK+7���g� Num Sel�W  F�#�� �Adju���60q.��%|� fe�ў�&tatu�!$6����%��  9 J�6RDM R�obot)�sco{ve2� 561��RemU�n@� �8 (S�F3Ser�vo�ҩ�)SNPX b��I�\dcs�0}�L�ibr1��H�� �5� f�0��5�8��So� tr�s�sag4%G 91E�p ��&0����p/I��  (i~g TMILIB(M<Ӌ�Firm�����gd7���s�Accd����0�XATXN�Heln��*LR"1x��Spac�A�rquz�imul�aH��� Q���To�u�Pa��I��T���c��&��ev.� f.svU�SB po��"�iuP�a��  r"1�Unexcept���`0i$/����H5-9� VC&�r��[6���P{��RcJP�RIN�V�; d �T@�TSP CS�UI�� r�[XC���#Web Pl6�%d -c�1�R�@4d�����I�R�66?0FV�L�!FVG�ridK1play C�lh@����5R�iR�R.@���R-�35iA���Ascii���"���� 51f�cUpl�� � (T����S���@rityAv�oidM �`��C�E��rk�CoYl%�@�GuF� 5P��j}P����
 B�L�t� 120C C�� o�І!J��P��yH��� o=q�b @oDCS b ./��c��O��q��`�; ����qckpaboE4�DH@�OTШ�?main N��19.�H��an.��A:> aB!FRLM����!i ���MI D�ev�  (�1� #h8j��spiJP�� � �@��Ae1/�r����!hP� M-2 � i��߂^0i�p�6�PC��  i�A/'�Passw�o�qT�ROS �4����qeda�SN��Cli����Gr6x Ar�� 47�!t���5s�DER��.�Tsup>Rt�I��7 (M�a�T2D�V�
�3D Tr�i-���&��_8t;�
�A�@Def?�����Ba: deRe p 4t0�Пe�+�V�st64MB DRAM��h86΢FRO�֫0�Arc� vi�sI�ԙ�n��7| �), �b�Hea�l�wJ�\h��Ce�ll`��p� �sAh[��� Kqw�c�G - �v���p	V,Cv�tyy�s�"�/�6�ut��v�m���xs ���T�D_0��J�m�` 2���a[�>R tsi��MAILYk�/�F2�h��ࠛ 90C H��F02]�q�P5'���T1C��5��F��FC��U�F9�OGigEH�S�t�0/A� if�!2���boF�dri=c ^�OLF�S�����" H5k�OP3T ��49f8���cro6��@ꊠl�ApA�Syn�.(RSS) 1�L�\1y�rH�L� (`2x5�5�d�pCVx9\����est�$SРl��> \pϐSSF��e$�tex�D o@���A�	� BP����a�(R00�Qirt��:���2)�D��1��e�VKb@l B�ui, n��WAP!Lf��0��Va�kTF�XCGM��D��L����[CRG&a�YBU��YKfL��p�f��k�\sm�ZT�Af�@�О�Bf2��и��V#�s���� r���CB���
f(���WE��!��
����T�p��DT��&4 Y�V�`��EaH����
�61Z���
�R=2�
�E (Np��F�V�PK�B��D�#��Gf1`?G����H�р?I�e �����LD�L��N��7\s@���`�z��M��dela<,���2�M�� "L[P��`?��_�%������S��-F�T�SO�W�J57η�VGF�|�VP2֥ 5\b�`0&@�cV:���T;T� ܨ<�ce,?VP�D��$
T;F���DI)�<I�a\so<��a-�6Jc6As6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P�
� ����`��Im'g PH�[l���I/A  VP�S��U�Ow��!%S�S>kastdpn)ǲt��� SWIMES5T�BFe�00��-Q�� �_�PB�_�Ru#ed�_�T�!�_�Sx ��_bH573ob2c2��-oNbJ5N�HIojb)�Cdo�cxE� �o�_�lp��o�TdP�o �c�B�or�2.rٱ`(Jsp�EfrSEop�f1�}�r3 RGoNeELS��sL�� ��s�����B	��S�\ $�F�ryz�ft	l�o~�g�o�����@����?�����P  �n�&�"�l ��T�@�<�^��Y��e�u8<Z���alib��Γ���ɟ3���埿�\v� ��e\c�6�Z�f8�T�v�R VW���98S��UJ91�����i�ů[c91+o�w8<���847�:� �A4�j��Q��t6�m���vrc.����HR���ot�0ݿ��'  ��8ޯ�3460�>eS0L��97���U�ЄϦ�60.� g�н�+��'��ܠ�Ϻ�8co��DM�߱U"�����ߕpì߲T! ��na;�� ���u%�����I��loR�d��1a59gϱŭ���95�ϔ�R����1 ��?��o�#��1A�/�d��vt{�UWeǟ����ￇ73[���7��ρ�C W��6I2K�=fR���8��@������d����2��ڔ����@�@"< "http������t7 �� v R7��78����p4�� ��TTPT�p#	��ePCV4/dv߀�j�Q�Fa7�b�$N�0�/2�rIO�p)/;/M/6.sv3��64i�oS�l? to�rah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��O�B4c.K?�g'�)�294g?�� (B�Ofd�\iOA5sb�?U_�?vi�/i��/�/BWn��`�o%�Fo��4l�$of��oXF sI)xo�cmp\7f��mp���duC��0lh����o(A�_Bt� �o]6P��m�I?�w��@���naO��4*O0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե1�1?o��DMs�B	C��7J�\���(�952�XFa AP�ڟ�<�v�`/şaqs8����/Of��I1�9�VRK�0��ph�քH5+�=�sIN/¤SkiW�/�IF��_�%�F�fs�I�O�l����"<𜿚$�`�����\jԿz5bO�vro�uς�3(�ΤH (DϮ��?sG��|��F �Ou�������D)O��*�3P$�FӅ�k���ϻ���럴� �PLx��ʿ��pbox��f�ebo���Sh �>�R.�0wT{����fx6��P��D��03��#_I\m;YE	e�OԆM�hxW�=E�te,���dct\���O$kR�����2�Xm*���ro3��D�l�j9��V<'�  FC����|@�ք f?6KA�RE0�_�~ (Kh��.cf���WcpoO�_K�up���a���H/j#- E�qd/�84���$qu�o��/ o2o?Vo"<�7C�)�s�NJԆx�|?�3l\sy�?0�40�?Τwio�u�]?�w58�?,F�0$OJ�
?Ԇ"io�!��V��u&A��PR��ߩ5, s��v1\�  H5352B�Q21p0�R78P51�0.R0  ne�l J614�Ҡ/WAT�UP��d8P545�*�H8R6��9�VCAM�q97PC�RImP\1tPUIF��C8Q28  in�gsQy0��4P P63rP @P PSCH��?DOCVڀD ��PCSU���08Q0�=PqpVEIO�Cr��� P54Pu;pd�PR69aP����PSET�pt\h�PQ`Qt�8P7`Q�!�MASK��(P�PRXY���R7�B#POCO  \pppb36���PR �Q��b1Pd60Q$c/J539.eHsb��?vLCH-`(��OPLGq\�bPQ0]`��P(`H�CR��4`S�au;nd�PMCSIP`e)0aPle5=Ps�p(`DSW� �  qPb0`0�aPa��(`PRQ`Tq0�RE`(Poa601P<cgPCM�PHcR0@q\j23b�V�`E`8�S`UPvisP`�E` c�`UPcPRS�	a�bJ69E`sF�RDmPsRMCN�:eH931PHcSNsBARa�rHLB�U�SM�qc�Pg52΁fHTCIP0cTMCIL�e"P�`eJ ��PA�PdSTPTXv6p967PTEL�p@��P�`�`
Q8P8$Q�48>a"PPX�8P915�P`[�95qqbwUEC-`F
PGUFRmPfahQCmP;90ZQVCO�`@�PVIP%�537nsQSUIzVSX�P��SWEBIP�SHT�TIPthrQ62�aP�!tPG���cIGt؁�`c�PGS�e�IRC%��cH76D�P�e Q�Q|�Ror��R51P s:P�P&,t53=P8u8=Py�C�Q6]`�b�PI��q52]`sJ56`E`s���PDsCL�q�Pt5�\rd�q7�5UP cR8���u5P sR55]`,s�  P8s��P�`CP�PP��SJ77P0\o��6��cRPP�cR�6�ap�`�QtaT�7�9P`�64�Pd87]`�d90P0c���=P,���5�9ta�T91P� ��1P(S��n�Qpai�P06=PW- C�PF�T	�0��!aLP PTS�pL��CAB%�I БI�Q` ;�H�UPPai-ntPMS�Pa��D��IP|�STY%�t\patPTO�b�P��PLSR76�`�5ؐQ��WaNN�Pai�c�qNNE`�OR�S�`�cR681Pi;nt'�FCB�P(��6x�-W`M�r��!�(`OBQ`plug��`L�aot �`O#PI-���PSPZ��PPG�Q7�`73nΒPRQadRL��(Sp�PSⳲn�@�E`��� �PTS-�� 8W��P�`apw�`���P`cFVR�PlcVs3D%�l�PBVI��SAPL�Pcycn+PAPV1�pa_��CCGIP - U���L�Prog+PC�CR�`�ԁB�P 4�PԁK=�"L�P��$p��(h�<�P��h��̱�@g�Bـ
TqX�%���CTC�p�tp��2��P927�"0ҝPs2�Qb��T�C-�rmt;�	`#�1ΒTC9`HcCT�E�Perj�EIPp.p/�E�P�c��I��use��Fـvr2v�F%���TG�P� �CP��%�d -h�H�-�Tra�PCTI��p��TL� TRS���p�@נ��IP�PuTh�M%�lexsQ{TMQ`ver, �p�SC:���F��Pv�\e�PF�IPSV"`+�H�$cj�ـtr�a�CTW-���CPVG�F-��SVP2mPv'\fx���pc�b���e��bVP4�fx_qm��-��SVPD-���SVPF�P_moҟ`V� cV��t\z��LmPove4��\-�sVPR�\|�tPV�Qe5.W`V 6�*u"��P}�o`���`N��CVK��N�IIP��CV����IPN9�Gene���D�@�D�R�D����  ��yf谔�pos.��/inal��n��D"eR���`��d�P��somB���on,��иR�D�R��\��TXpf��D$b��omp��G "N��P��m����! ��=C-f8����=FXU�����g F��(��Dt� II��r�D��u��� "����Cx_�ui X������fa2��h	Crl2��D,r9ui�Ԣ�� it2c�0c�o��e"�����ާ(.)� ��{�� ��� �IQnQ �I�[ ��_= wwo��,bD� ���|GG�� �����4� �e� v�ʷ� ��&�� 2��Z uz������� �w�TW&q~q �5�׷&�o?� ;0��  �{2� �y� ����W&���� ?�3� A���e�/> �{\�3&T��� �77߸ ��ֽ� ���� �{���&��8 ��l1��S�)� ���d *{J� F's �~��� 6:0�� ��,��s�- Q�v� ���� �,�T� �ZBLx6����6 ��6���N�Par ��s>�tE��j�6dsq��F  �������ЁDhel�����ti-S�� �Ob��Dbcf�O�����+t OFT��P<A� _�V�ZI��D��V�\�qWS��= dt�le�Ean�(bz=d��titv�Zҥz�Ez XWO �H6�6���5 H^�6H691�E4܀�TofkstF� Y6�82�4�`�f80M4�E91�g�`30oBkmon_�E��e�ݱ�� qlm��0� J�fh��B�_ / ZDTfL0�fw(P7�EcklKV0� �6|��D85��ّ�m\b����xo�kn�ktq��g2.g����yLbkLVtms��IF�bk��x����Id I/f���GR� �han�L��Vy��%��%ecre�����io��w ac�- A�qn�h���cuACl�_�^ir��)�g�2�	.�@�& G��R630���p v�p`�&H�f��un���R57v�OJavpG�`Y��owc��-ASF��O��7���SM�����v
af��raf�La�vl�\F c�w a���?VXpoV �{30��NT "L�FFM��=����yh	�a�G-�w�� �m�2.�,�t��̹�g6ԯ��sd_�#MC'V����D����fslm�isc�.  Hg5522��21&d�c.pR78�����0�708�J614Vip ATUu�@�OL�545ҴI�NTL�6�t8 (�VCA���sseCRI���ȑ��UI���rt\�rL�28g��NRmE��.f,�63!���,�SCH�d Ek�DOCV���p���C,�<�L�0Q�isp��EIO��xE,У54����9��2w\sl,�SETĸ��lр�lt2�J�7�ՌMAS�K��̀PRX�Y҇��7���OC-O��J6l�3�l�� (SVl�A�H�pL�@Օ��539R�sv���#1��L�CH���OPLG.f�outl�0��D��HCR
svgb��S@�h��CSaԌ!�{�50��D�l�5�!�lQ��DSW��S0����̀��OP����M7��PR���L�Ҟ��(Sgd���P�CM���R0 \Es��5P՝���0��X��n�q� AJ�1��tN�q�2��PRSa����69�� (AuFRD�Խ���RMCN���93�A�ɐCSNBuA�F9� HLB���� M��4���h�2vA�95z�HTCa�ވ�TMIL6�j9y5,��857.,�PA1�ito��T�PTXҴ JK�T�EL��piL�� 4XpL�80�I)��.и!��P;�J95��s� "N���H�UE�C��7\cs�F�R��<Q��C��57\{VCOa�,����IP1jH��SU�I�	CSX1�A�WEBa��HT�Ta�8�R62��md`��GP%�IG %�tutKIPGS�j�| RC1_meN�H76��7P��ws_+�?x�R51�\iw�N��ԦH�53!��wL�8!�h�R66��H����Ԡ���@;J5�6��1���N0��9�j2��L���R5`%�AJ|�5q�r�`,�8 5���{165!��@�"5l��H84!�29��Ⱦ0��PJ���n �B[�J77!Ԩ�RA6�5h3n���y36P��3R6��-`;о Ը�@��exeKJs87��#J90!��stu+�~@!䬵��k90�kop �B����@!�p�@|B�A�g*�n@!��Q��06!�@[�F�FaP��6��́,�TS� �NC[�CAB$i4Ͱl1I��R7��@�q�y�CMS1�r�og+QM�� �� T�Y$x�CTOa�n�v\+��1�(�,�6��con�~0��1]5��JNN�%e:�8�P��9ORS%xк��8A�815[�FCBaUnZQ�P!��p�{��CMOB��"�G��OL��x�OP]I�$\lr[�SŠ��T	D7�U��CPRMQR9RL���S�V��~`���K�ETS �$1��0���3�Ԯ��FVR1�LZQVc3D$ ���BVa��SAPL1�CLN�[�PV��	rCCG�aԙ��CL�3C{CRA�n "W!�B�H�CSKQn�\0�p��)�0CTPn�ЌQe��p!$bCt�aT0U�pGCTC�yЋRC1��1 (�s��trl�,�r��
TX��T�Caerrm�r�M�C"�s��#CTE���nrr�REa�XqPj�^��rmc�$^�a"�P�QF!$�\��$p "�rG1䖈tTG$c8��QHܑ$SCTI�! �s��CTLqdAC�K�Rp)��rLa�R82��M��YPk�.���OF��.���e�{��CN���^�1�"M �^�a�С�Q`US��T!$��M�QW�$m��VGF�$R MHv��P2�� H5� �ΐq��ΐ�$(MH[�VP�uoY����$�)��D��hg��V{PF��"MHG̑�`e!�+�V/vpcm��N��ՙ�N��$�VcPRqd)��CV�x�V� "�X�,�1�(${TIa�t\mh��K��etpK�A%bY�VP%ɠ�!PN����GeneB�ri�p����8��e�xtt���Y�m �"�(��HB�� �)��x������x�Ȣ�res.�yA�ɠn�����*���p�@M�_�NĀ6L���Ș�yAvL�Xr�Ȉ2��s"R;�Ƚ\ra���	P�� h86��Gau+ʸ�Ͽ�SeL��m�9�69�P�Ȩr`�Ȩ2�ɹ1��n2��h� �0L�XR}�RIB{�e� L�x���c�Ș���N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1��/�k�@���A���ruk�ʘ L�so1p��H�}�ts{���ĺ��s��9��j965��Sc��h��O5 J9�{�
�P�L�J	een��ts I[
x�com��9Fh�L�4 J�v�fo��DIF+��6�Q����rati�|��p��1�0�
R8l߾�M�����P��!8� �j�mK�X� HZ����N��oڠ��3�q��vi̋��80�~�l aSl�yQ��tpk�xb�j�.�@�R�d�������,/n(�8�8 �0���
:�O8�<�LQ}�CO���PT��O (��.�Xp|��~H���?�v f�wv��8�22�p�m���722��j�7�^�@ƙ���cf��=Yvr���vcu���O�O�O�O_�#_5_7�3Y_��wv�4{_�_w�ʈ�u�st_�_�cus �_�Z��oo,o>oPo8�io��nge��(p�Ly747�jWel�ʨHM47ZKEq� {���[m�MFH�?�(wsK�8J��n���o��fhl�;��wmf���? �:�}(4	<g J�{��II)̏މw��X�774kﭏ/7�ntˏ݊e+���se�/�aw��8�ɐR��EX \�!+: �p,��~�00��nh�,:�Mo+�xO��1 "YK�O��\a��#0 ��.8���{h�L?�j+N�mon�:��t�/&�st�?-�w�:� ��)�;��(=h�;
�d Pۻ�{:  ��� �J0���re����S�TD�!treLANG���81�\tqd�������rch.��ռ���htwv�WxWָ� R79���"Lo�51 (��I�W�h�Ո�4�aSww� �vy ��623c�h a?�cti�֘!�X��iؠ�t ��n@,�։����j��"AJP@�3p�Svr{�H�6��!��o- SeT� E3ּ) G�J934��L=oW�4 (S����p��� <���91 ��8!4�j9�所+��ٲy�
��	�btN�ite{�R ��I@� ������P�������p	 ����Z�vol���X ��9�<�I�p���l�d*���F�864{��?��K�	�k�����֘1�wmsk���M�q�Xa�e ����p��0�RBT�1ks.OPTN�qf�Uz$ RTCamT ��y��U��y��U��UlU6L�T�1 Tx����SFq�U�e�6T��USP W�b DT�qT2h�T�!/&+��TX�U\j6&�Up U�UsfdO&��&ȁT���66�2DPN�b0i��%�Q�%62V��$����%�� �#(�(6T=o6e St�%���#5y�$�)5(T�o�%tT0�%5�W6Tp���%�#�#orc���#I���#���%ccat�6ؑ?�4\W6�965"p6}"�#\j536���4�"�?GkruO O,Im?Np�C �?t�0<O�;�e �%���?
;{gcJ7 "AV�?�;avsf�O__�&_8WtpD_V_0GT��F|_:UcK6�_�_r��O�3e\s�O2^y\`O:�migxGvgW'! m�%��!�%T�$E A{6�po6�f�#37N�)5R5_�2E���$0���$Ada�Vd���V�?;Tz78�_�e7DDTF9���#8�`�%��4y�?ted Z@�A}�@�}�04N�}�}���}�dc& }���	�u 6�v��v1�u1\b�u$2}���}� R83�u�"}�<�"}�valg���Nrh�&�8�J�Y��o�ue��� j70��v=1��MIG�uerfa��{q���E�qN�ء��EYE�ce A���񁏯p V�e�A!���2Յ�Q�%��u1�e�i�@��H� e����J0� '��bx��T��E In��B�  W�|��53q7g����(MI��t�Ԇr��ݟ�a!m���nеv!g�U -�v J߆8⹖F���P�y�ac���2���Rɏ jo��2��� djd�8r}� Gog\k�0��g��wmf�Fro�/� Eq'�4"}�3� J8��oni�[��ᅩ}Ĵ�� !o� ��ʛ��m@�RΉe��{n�Д�V�o������  �����裆"PO�S\����ͯ me�nϖ�⑥OMo�4q3��� �(Coc� An[�t���"e��a\�vp��.��c7flx$�le��8ٰhr�tr�NT� �CF+�x E/�t0	qi�M�ӓxc��p��f�lx����Z�cxb��
0 h��h8��3mo��=� H����)� (�vSER,����g�0߆0\r��vX�= ��I � -� �ti��H��V]C�828�5���L"�RC��n G�/���w�P�y�\v�vm "o�lϚ�x`а�=e�ߠ-�R-�3?������vM [�A�X/2�)�S�rxel�v#�0��h8߷^=� RAX�A�����9�H�E/R�צ����h߶"RXdk��F�˦85���2L/�xB885t_�q�Ro�0iA��5\rO�9�K��v�����8���.�n� "�v��88��8 s�i ?�9 ��/p�$�y O�MS"�x��&�9R H74&�`�745�	p��8p��ycr0C�c�)hP0� j�-�a%?�o��6D950R7tr�l��ctlO�AcPC���j�ui"��L���  ����^%棆!�A��qH��z�&-^7����w ��616C��q�794h���� qM�ƔI��99����(��$FE�AT_ADD ?_	���Q%P?  	�H._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n ���������TDEMO �fY    WM_���� ����//%/R/ I/[/�//�/�/�/�/ �/�/�/?!?N?E?W? �?{?�?�?�?�?�?�? �?OOJOAOSO�OwO �O�O�O�O�O�O�O_ _F_=_O_|_s_�_�_ �_�_�_�_�_ooBo 9oKoxooo�o�o�o�o �o�o�o>5G tk}����� ���:�1�C�p�g� y�������܏ӏ��� 	�6�-�?�l�c�u��� ����؟ϟ����2� )�;�h�_�q������� ԯ˯ݯ���.�%�7� d�[�m�������пǿ ٿ���*�!�3�`�W� iϖύϟ��������� ��&��/�\�S�eߒ� �ߛ��߿�������"� �+�X�O�a���� �����������'� T�K�]����������� ������#PG Y�}����� �LCU� y������/ 	//H/?/Q/~/u/�/ �/�/�/�/�/??? D?;?M?z?q?�?�?�? �?�?�?
OOO@O7O IOvOmOO�O�O�O�O �O_�O_<_3_E_r_ i_{_�_�_�_�_�_o �_o8o/oAonoeowo �o�o�o�o�o�o�o 4+=jas�� ������0�'� 9�f�]�o��������� ɏ�����,�#�5�b� Y�k���������ş� ���(��1�^�U�g� �������������� $��-�Z�Q�c����� ��������� �� )�V�M�_όσϕϯ� ����������%�R� I�[߈�ߑ߫ߵ��� ������!�N�E�W� ��{���������� ���J�A�S���w� ������������ F=O|s�� ����B 9Kxo���� ��/�/>/5/G/ t/k/}/�/�/�/�/�/ ?�/?:?1?C?p?g? y?�?�?�?�?�? O�? 	O6O-O?OlOcOuO�O �O�O�O�O�O�O_2_ )_;_h___q_�_�_�_ �_�_�_�_o.o%o7o do[omo�o�o�o�o�o �o�o�o*!3`W i������� �&��/�\�S�e�� ������������"� �+�X�O�a�{����� �����ߟ���'� T�K�]�w��������� �ۯ���#�P�G� Y�s�}��������׿ ����L�C�U�o� yϦϝϯ�������� 	��H�?�Q�k�uߢ� �߫���������� D�;�M�g�q���� ������
���@�7� I�c�m����������� ����<3E_ i������ �8/A[e� �������/ 4/+/=/W/a/�/�/�/ �/�/�/�/�/?0?'? 9?S?]?�?�?�?�?�? �?�?�?�?,O#O5OOO YO�O}O�O�O�O�O�O �O�O(__1_K_U_�_ y_�_�_�_�_�_�_�_ $oo-oGoQo~ouo�o �o�o�o�o�o�o  )CMzq��� ������%�?� I�v�m����������ُ���;�  2�Q�c�u����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�9� K�]�o����������� ������#5GY k}������ �1CUgy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o�o�o�o +=Oas��� ������'�9� K�]�o���������ɏ ۏ����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������ +=Oas��� ����'9  :>U gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����� ����/�A�S�e� w���������я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{�����@��/=C6Yk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/AS ew������ �+=Oas �������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�� ������!�3� E�W�i�{�������Ï�Տ�����/�A���$FEAT_DEMOIN  E���q��>�Y�I�NDEXf�u���Y�ILECOMP g������t�T���SETUP2 h������  N� ܑ��_AP2B�CK 1i�� � �)B���%�C�>���1�n�E� ���)���M�˯���� ���<�N�ݯr���� ��7�̿[��ϑ�&� ��J�ٿWπ�Ϥ�3� ����i��ύ�"�4��� X���|ߎ�߲�A��� e�����0��T�f� �ߊ�����O���s� ����>���b���o� ��'���K������� ��:L��p���� 5�Y�}�$� H�l~�1� �g�� /2/�V/ �z/	/�/�/?/�/c/ �/
?�/.?�/R?d?�/ �??�?�?M?�?q?O��?O<O���P�� 2�*.VRCO�O�0*�O�O�30�O�O�5w@PC�O_>�0FR6:�O=^�Oa_�KT���_�_�&U�_�\h�R_�_�6G*.FzOo�1	(S�oEl�_io�[STM �b�o�^+P�o�m��0iPend�ant Pane	l�o�[H�o �gp�oYor�ZGIF|���e�Oa��ZJPG �*��e����z��JJS�����0�@���X�%
JavaScriptُ�CSʏ1��f�ۏ� %Casca�ding Sty�le Sheet�s]��0
ARGN?AME.DT���<�`\��^���Д����АDISP* ן���`$�d��V�e���CLLB.Z�I��=�/`:\��\������Coll�abo鯕�	PA�NEL1[�C�%@�`,�l��o�o�2a��ǿV���r����$�3 �K�V�9���ϝ�$�4i���V���zό�!����TPEINS.gXML(�@�:\<�����Custom� Toolbar�}��PASSWO�RD���>FRS�:\��� %P�assword ?Config��? J���C��"O��3��� ��i����"�4���X� ��|�����A���e� ����0��Tf�� ���O�s ��>�b�[� '�K���/� :/L/�p/��/#/5/ �/Y/�/}/�/$?�/H? �/l?~??�?1?�?�? g?�?�? O�?�?VO�? zO	OsO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_;_M_�_q_o�_ �_<o�_`o�_�o�o%o �oIo�o�oo�o8 �o�on�o�!�� W�{�"��F�� j�|����/�ďS�e� ��������T��x� �����=�ҟa���� ��,���P�ߟ񟆯� ��9����o����(� :�ɯ^�����#��� G�ܿk�}�ϡ�6�ſ /�l�����ϴ���U� ��y�� ߯�D���h� ��	ߞ�-���Q߻�������,��$FIL�E_DGBCK �1i������ ( ��)
SUMMA�RY.DG,����MD:`�����Diag Sum�mary���
C?ONSLOG��y������$���Con�sole log�%���	TPACC�N��%g������TP Accou�ntinF���F�R6:IPKDM�P.ZIP����
���)����Exception-�����MEMCHECKК����8�Me�mory Dat�a��LN�)�RIPE����0�%� Packet LE����$Sn�ST�AT*#� �%LStat�us�i	FTP��/�/�:�m�ment TBD�=/� >)E?THERNE�/�o�/�/��Eth�ernU<�fig�uraL��'!DCSVRF1//)/B?��0 veri?fy allE?��M(5DIF�F:? ?2?�?F\8d�iff�?}7o0CHGD1�?�?�?LO� �?sO~3&��
I2BO)O;O�O qbO�O�OGD3�O8�O�OT_ �O{_�
VUPDATE�S.�P�_��FR�S:\�_�]��U�pdates L�ist�_��PSRBWLD.CMo����Ro�_9�PS�_ROBOWEL<^/�/:GIG��o�>_�o�GigE� ��nostic�W�N�>�)>�aHADOW�o�o��ob�Shad�ow Changye��8+"rNOTI?=O���Notifi�c�"��O�A�PMIO�o���h��f/��o�^U�*�UI3�E�W��{�UI������B��� f��_�������O�� �������>�P�ߟt� �����9�ί]�򯁯 �(���L�ۯp���� ��5�ʿܿk� Ϗ�$� 6�ſZ��~��wϴ� C���g���ߝ�2��� V�h��ό�߰���Q� ��u�
���@���d� �߈��)��M����� �����<�N���r�� ��%�����[���� &��J��n�� 3��i��"� X�|��A �e�/�0/�T/ f/��//�/=/�/�/��$�$FILE_��PPR�P���� �����(MDONLY �1i5�  
 �z/Q?�/u?�/�? �?t/�?^?�?O�?)O �?MO_O�?�OO�O�O HO�OlO_�O_7_�O [_�O_�_ _�_D_�_ �_z_o�_3oEo�_io �_�oo�o�oRo�ovo �oA�oew �*��`����&�O��*VISB�CK,81;3*.�VDV����FR�:\o�ION\DOATA\��/���Vision VD filȅ ��&�<�J�4�n��� ���3�ȟW������ "���F�՟�|���� ��m�֯e������0� ��T��x������=� ҿa�s�ϗ�,�>��� b���ϗϼ�K��� o��ߥ�:���^�����ϔ��*MR2_G�RP 1j;�C4  B�}Ї	 71������E��� E�  F@ F�5U�������L���M���Jk�L�zp�JP��F�g�f�?�  �S����9�Y9�}�9��8�j
�6��6��;��A�  l���BH��B���B���$��������������@UUU#�����Y�D�}�h� ���������������
C��_CFG {k;T M����]�NO �:
F0� �� \�RM_CHK�TYP  0��}�000��OM�_MIN	x����50X� S�SBdl5:0��bx�Y����%TP_DEF_�OW0x�9�I�RCOM��$�GENOVRD_�DO*62�TH�R* d%d�_�ENB� �R�AVC��mK�� ��՚�/3�/�q�/�/�� �M!kOUW s��}���ؾ��8��g�;?�/7?Y?[?  C��0����(7�?6�<B�?B����2p��*9�N SMTT#�t[)��X�4�$HoOSTCd1ux����?�� M5Cx��;zOx�  27.0�@=1�O  e�O�O 	__-_;Z�O^_p_�_�_�LN_HS	ano?nymous�_�_�_oo1o yO��FhFk�O�_�o�O�o�o �o�oJ_'9K] �o�_����� 4o�XojoG�~�o^� ������ŏ���� �1�T���y����� ������,�>�@�-� t�Q�c�u��������� ϯ���(�^��M� _�q�����ܟ� �ݿ ��H�%�7�I�[Ϣ� ϑϣϵ����l�2� �!�3�E�Wߞ���¿ Կ����
������� /�v�S�e�w���� ���������+�r� �ߖ�s�����߻��� �������'9K] ��������� 4�F�X�j�l>��} ������/ /1/T��y/�/�/�/�/.D\AENT {1v
; P!J/.?  ��/3? "?W??{?>?�?b?�? �?�?�?�?O�?AOO eO(O�OLO^O�O�O�O �O_�O+_�O _a_$_ �_H_�_l_�_�_�_o �_'o�_Koooo2o{o Vo�o�o�o�o�o�o 5�oY.�R��v��zQUIC�C0���3��t1 4��"����t2��`��r�ӏ!ROUT�ERԏ��#�!�PCJOG$����!192.16?8.0.10��s?CAMPRTt�P��!d�1m�����R�T폟�����$NA�ME !�*!�ROBO���S_�CFG 1u�)� �Au�to-start{edFTP&��=?/֯s��� �0�B��f�x����� ����S������,� ��������ϼ�ޯ�� �������ʿ'�9�K� ]�oߒ�ߥ߷����� ����(:~�k� �Ϗ���������� ��1�C�f���y��� ���������,�>� R�?��cu��`� ����(�$ M_q������  /H%/7/I/[/ m/4�/�/�/�/�/� ~/?!?3?E?W?i?� ���?�/�?/�?O O/O�/�?eOwO�O�O �?�ORO�O�O__+_ r?�?�?�?�O|_�?�_ �_�_�_o�O'o9oKo ]ooo�_o�o�o�o�o �o�oF_X_j_~ok �_������o� ��1�TU��y����������U�)�_ER�R w3�я�P�DUSIZ  jg�^�p���>�?WRD ?r�Cq��  guestb�Q�c�u��������"�SCDMNGRP 2xr�w���Cq�g�\�b�K� 	�P01.00 8~(q   �5p��5pz�5pB � �{ ����H���L���L��L�����O�8�����l�����a�4� x��Ȥ�x��V8���\���)�5`�;��������d�.�@�R�ɛ_�GROUېy������	ӑ���Q?UPD  ?u��Y��İTYg�����TTP_AU�TH 1z�� �<!iPend�an��-�l����!KAREL:q*-�6�H�KC]��m��U�VISI?ON SET���� ��g�G�U������R� 0��H�Bߏ�f�x�����߮���CTRL C{����g�
S��FFF9E3���AtFRS:D�EFAULT;��FANUC W�eb Server;�)����9�K��܀����������߄W�R_CONFIGw |ߛ ;���IDL_CPU�_PCZ�g�B��Dpy� BH_�MI�Nj�)�}�GNR_�IO��g���a�N�PT_SIM_D�_�����STAL�_SCRN�� ����TPMODNT�OL������RTY`��y���� �ENO����Ѳ]�OLNK 1}��M���������eMA�STE��ɾeSL?AVE ~��c>�O_CFGٱ�BUO�O@CY�CLEn>T�_A�SG 1ߗ+�
 ����// +/=/O/a/s/�/�/�/��/��NUM�z�
@IPCH��^RTRY_CN Z���@��������� @kI��+E�z?E�a�P_M�EMBERS 2Y�ߙ� $���2����ݰ7�?�9a�S�DT_ISOLC�  ����$J_23_DSM+��3JOBPROC�N��JOG��1��+�d8G�?��+�O�/?
�LQ�O__/_�O S_e_w_�_`�O H�m@��E#?&BPOS�REQO��KANJ�I_���a[�MON ����b�yN_goyo�o�o�o�$Y�`3�<� ��e�_ִ��_L���"?`�EYLOGGIN�LE��������$LANGUAGgE ��<T�Y {q�LGa2�	��b���g�xP�� � ��g�'Զ�b���>�M�C:\RSCH\�00\<�XpN_D?ISP �+G�pJ��O�O߃LOC�p�Dz���AsO�GBOOK �������󑧱����X�����Ϗ���`�a�*��	p� ����!�m��!���=p�_BUFF 1�p��2F幟����՟D� Col�laborativǖ���F�=�O�a� s�������֯ͯ߯����B�9�K���DC�S �z� =���'�f��?ɿۿ����H@{�IO 1��� ~?9ü�� 9�I�[�mρϑϣϵ� ���������!�3�E� Y�i�{ߍߡ߱����ߴ���E��TMNd �_B�T�f�x���� ����������,�>� P�b�t�������L��SEVD0��TYPN1�$6���QRS"0&��<2�FL 1�"�J0���������GTP:pO>F�NGNAM1D��mr�tUPS�GI�"5�aO5�_LO{ADN@G %��%TI�pZUZ�AUN#�(MAXUALRM�'���(���_PR"4F0�d��1�B_PNP�� V 2�C	�MDR0771�ߕ�BL"806=3%�@ �_#?�hߒ|/�C��z��6��/���/Po@P �2��+ �ɖ	�T 	t  ��/�%W?B?{?� k?�?g?�?�?�?O�? *OONO`OCO�OoO�O �O�O�O�O_�O&_8_ _\_G_�_�_u_�_�_ �_�_�_o�_4ooXo joMo�oyo�o�o�o�o �o�o0B%fQ �u������ ��>�)�b�M����� {��������Տ�� :�%�^�p�S��������D_LDXDI�SApB�MEM�O_APjE ?=C
 �,� (�:�L�^�p�������� 1�C � ���4�������4���X���C_MST�R ���w�SC/D 1���L�ƿ H��տ���2��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v� aߚ߅ߗ��߻����� ��<�'�L�r�]�� ������������� 8�#�\�G���k����� ����������"F 1jUg���� ���B-f�Q�u���h�MKCFG �����/�#LTARM_*��7"0��0N/V$� METP�Uᐒ3����ND>� ADCOLp%� �{.CMNT�/ �%� ����.E#�>!�/4�%POSC�F�'�.PRPMl�/9ST� 1���� 4@��<#�
1�5�?�7{?�? �?�?�?�?�?)OOO _OAOSO�OwO�O�O�O�O_�A�!SING_CHK  �/�$MODAQ,#�����.;UDEV �	��	MC:>o\HSIZEᝢ���;UTASK �%��%$1234?56789 �_�U�9WTRIG 1�
��l3%%��9o��"o0coFo5#�VYP�QNe���:SEM_IN�F 1�3'� `)AT?&FV0E0po�m�)�aE0V1&�A3&B1&D2�&S0&C1S0}=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o' ��K������� я:�L�3�p�#�5��� Y�k�}������$�[� H���~�9�����Ư د��������ӟ�V� 	�z�������c�Կ�� ��
��.���d�� )�;��Ͼ�q����� ��˿<���`�G߄ߖ� IϺ�m�ϑϣ���� 8�J��n�!ߒ�M��������h_NITO�R� G ?�[  � 	EXEC�1�/�25�35�4�5�55��P7�75�8
5�9�0�Қ�4� ��@��L��X��d� ��p��|�������2��2��2��2���2��2��2��2���223��3��3@�;QR_GRP_SV 1��k� (�A�z�4��~�K��������K:z�j]�Q_D��^��PL_NAME �!3%,�!�Default �Personal�ity (fro�m FD) �R�R2� 1�L?6(L?�,0	l d���� ����//(/:/ L/^/p/�/�/�/�/�/�/�/ZX2u?0?B? T?f?x?�?�?�?�?\R<?�?�?O O2ODO�VOhOzO�O�O�OZZK`\R�?�N
�O_\TP�O:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHo_)_~o�o �o�o�o�o�o�o  2DVhz�[omo ����
��.�@� R�d�v���������Џ�� Ef  Fb� F7���   ��!��d��@�R�6�t��� ���l���ʝ����� ݘ���� "�@�F�d���� "�|��ݐA�  ϩ�U[�$n�B��E ��� � @D�  &�?�� �?�@��A@�;f��FH�� ;�	l,�	 '|��j�s�d�/>��� ��� �K(��Kd$2�K ��J7w��KYJ˷�ϜJ�	�ܿ�� @�I���_f�@w�z��f򿿾γ�N�������	Xl�����_��S�ĽÔ�}�I ����5�?��  ����A�?oi#�;����� ���l� �Ϫ�-���ܛ�G�G�Ѳ��@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=�����в@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj��a�Be�Ci��#��Bи�ee^��^^ȹBР ��P����̠�����ADz՟�n�3��C��i�@�R�R�Y���� { �@� ����  ���?�ff0������n� ɠ #ѱy9G
(���I�	(�@uP~����t��t���>����;�C�d;��.<���<�g�<F+<L�������,��d�,�̠?fff�?��?&&��@���@x��@��N�@���@T�H�ِ�!-�ȹ �|��
`���� ���//</'/`/`r/]/�/��eF�� �/�/�/�/m?��/tJ?�(E��G�#�� FY�T?�?P? �?�?�?�?�?O�?/O O?OeOk��O�IQO G�?�O1?�OmO_0_�B_T_������A _�_	_�_�_�_ o���A��An0 bФ/o �C�_Uo�_�Op���؃o�o�o�o���W������oC�E�� q�H�d�����a@q��e�F�Bµ�WB]�NB2��(A��@�u�\?�D��������b�0�|�u�R����
x~��ؽ��B�u*C��$�)�`�$ ����GC#����rAU�����1�eG�D�I��mH�� I:��I�6[F�﫹C�I���J�:\IT��H
~QF�y���p�*J��/ I8Y�I��KFjʻCe �o��s�����Џ��� ߏ�*��N�9�r�]� �����������۟� ��8�#�\�G�����}� ����گů���"�� �X�C�|�g�����Ŀ �������	�B�-� f�Qϊ�uχ��ϫ��� �����,��P�b�M� ��qߪߕ��߹����� ��(��L�7�p�[��@�������s($�ϳ�3:����$���3���d�,��4��@�R�wa�ǲ��l�~�wa����e����wa4 �{������(L�:ueP�P~�A �O������	����G2 W}h����� �/���O�O7/m/[(d=�s/U/�/�/�/ �/�/?�/1??U?C?�y?�=  2 E�f9gFb��77�b9fB)aa)`C9A`	�&`w`@-o�?w`e�@O)O�?MO�Ow`�?@�?�O�O�O�O9c?�0T�A7ht4w`w`�!w`xn
  �O9_K_]_o_�_�_�_ �_�_�_�_�_o#ozz�Q ��h��G����$MR_CA�BLE 2�hO �a�T� @@�0�Ae��a�a��a��`��0�`C��`�aO8�tB�^n�d��`�aE�4�E�#��o�f�#��0�|�0�DO��By`���Š��bED4E�c,��o�g8  ���Cu�07�d4
v�ے�0 �b���XE�Z&�lȠ`y`
qC�p�bHE݈
v#g�5DͣҮ�qz�lҠ`�p�0�q�p�b0�
v׸%c���b=%	E;h��u/o�c -��4tH�\�?�9�K� ]�o�ԏϏ��
�ɏۏ�@���?��eo �a���������b����� �����`�	 ���������`�� ���퐺@�����ŀ�U�ݐ����������������*,� ,�-�\c�OM �ii���3� � �]0%% 23�45678901�i�{� f��������ԋ��1����
���`�not �sent3������;�TEST�FECSALGRG  e�qiG�1d.�Zš
:�� �D�CbS�Q�c�u��� 9�UD1:\ma�intenanc?es.xml��ֿ�q� =���DEFAULT�-�i4\bGRP 2�M�  =��a����   �%Force��sor chec�k  ���b�z��p����h5-[ �ϻ��������dID�%!1�st clean�ing of c�ont. v�i?lation��}�Rߗ+��[�ߔߦ������mech��cal`����B��0��h5k߀@�R�d�v�����(�rolle_Ƶ�����/���(�:�����Basic �quarterl!y�������,����`������M��M��:C@"GpP�a�b`i4��������#C���M"���{Pbt����Suppq�gre�ase����?/&/8/J/\/��C�+ ge��. ba�tn�y`/��/h5	 /�/�/�/? ?_���en'�v��/�/��/��?�?�?�?�?F�G=?O�qp"CrB1O��0�/`OrO��O�O�O�t$��Lf���C-m��A�O:��OO$_6_H_Z_l_��t*cabl�Om����S<m��Q�_:�
 _�_�_oo0oo)(��/�_�_���_�o�o��o�o�o�O@h�au1�l�2r !xm�<qC:��op�������ReplaW�fUȼ2�:�._4�F�X�j�|�m�$%���o������� #���
��.�@���d� ��ŏ׏����П��� �U�*�y�����r��� ������	�q��?�߯ c�8�J�\�n���ϯ�� ���ڿ)����"�4� Fϕ�jϹ�˿����� �������[�0�ϑ� fߵϊߜ߮�����!� ��E�W�,�{�P�b�t� ����߼�����A� �(�:�L�^������ �������� $ s�H������q�� ���9]o� Vhz���U� #�G/./@/R/d/ ��/�/��//�/�/ ??*?y/N?�/�/�? �/�?�?�?�?�???O c?u?JO�?nO�O�O�O8�O+J�r	 H�O�O __6M2_@OBE:_p_ >_P_�_�_�_�_�_ o �_�_oHoo(oZo�o ^opo�o�o�o�o�o ��o :z �bA?�  @�q  _���Fw��� �H* �** @q>v�p2T�f�x��:�������ҏ�� eO^C7�Տ#�5�G�	� k�}���ُ���c�� ���W��C�U�g��� ß)�����ӯ���	� �-�w�����9����� ��m�Ͽ��=�O�E�	A�$MR_H�IST 2�>u�N�� 
 \�$Forc�e sensor� check  �12345678�90q�3�������N}SB�� -319.8� hours R�UN 9.�Y�!�1st clea�ning of �cont. ve�ntilatio�n0ÄϖϨ�-�� $��mech���cali�%Ό4���o�DN�t&��95��1����rolleh�+�=��O���Bas�ic quarterlyߒߤ߶� 
O4�F��(���� ��b�t���������� �M�_����:������p���:�SKCFM�AP  >u�Q��r5��������ONREL  .�3���?EXCFEN��:q
��QFNCX�JJOGOVLI�M8dNá ��KE�Y8��_PAN7����������SFSP�DTYPxC��S�IG�:��T1M�OT�G��_C�E_GRP 1�>u\�D�� ���/Ⱥ��/ �/U//y/0/n/�/ f/�/�/�/	?�/??? �/c??\?�?P?�?�? �?�?�?O)OOMO,����QZ_EDIT�5 )TCOM_�CFG 1����[�O�O�O 
�ASOI �y3�
__+[_O_���>O�_bHT_AR�C_UքT_MN_MODE5��	UAP_C�PL�_gNOCH�ECK ?�� �� o.o@o Rodovo�o�o�o�o�o��o�o*!NO_WAIT_L4l~GiNT�A���|EUwT_ERRs2���3��ƱJ������>_)��|MO�s��}x:Ov���?8�?������ l��rPARAuM�r������j���5�5�G� =  r�b�t�s�X��� ���������֟�0����b�t������SUM_RSPA�CE�����Aѯۤ�$ODRDSP�S�7cOFFSET�_CARt@�_�D�IS��PEN_FILE:�7�AF��PTION_I�O��q�M_PR�G %��%$*�����M�WORK ��yf �!�춍�����r����	 �������gT��RG_DSBL  ���C�{u��RIE�NTTO7 ��Cٴ A �UT�_SIM_Dy����V�LCT ��}{B �٭�ď_PEX�P=��R[AT�W dc�>�UP ���`���e�w�]ߛߩ���$�2r�L�6(L?���	l d������ &�8�J�\�n���� �����������"�4�F�X���2�߈����� ��������*�<w�Tfx��������J`�ˣG���Tz�Pg���� ��/"/4/F/X/j/ |/�/�/�/���/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?�/�/ ,O>OPObOtO�O�O�O �O�O�O�O__(_:_��O��y_�]2����_�^�_�_�W^]@^]��/ooSog� Hgrohozo�o�o�o�o��oF`�#|`�AG�  9y����OK��1�k�����<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	 '|�Q�s�r�q/>��u �sF`�H<zH~��H3k7GL�z�HpG�9�9l7�k_B�T�F`C4T��k�H���t��-��Ae���k������s���  ��ሏ����EeBVT����dZ��g���ڏ ����q-�Fk�y�{FbZU���n@6�_  ���z��Fo��Be	'� �� ��I� ��  �:p܋=����ڟ웆�@���B�,���B��g�AgN���� � '|���g��B�*��p�BӀC׏�����@  #�B�u�&�ee�^^މB:p2����>�m�6p�Z���Dz ?o}�܏������׿�������Ǒ��� f� � � �M���*�?�ff�_8�Jφܿ 3pϑ�ñ8@�Чϵʖq.·�(����P���'��s�tL��>��/�;�Cd;���.<߈<��g�<F+<AL ��^oiΚrd@�|�r6p?fff?��?&�п�@���@x��@�N��@���@T� ��Z���ћtމ�u�� �w	�x��ti�>�)�b� M��q��������� ����:�%�^��������W���S�E�  �G�aF�� Fk���������1 U@yd���� ��q��	��{�A ��h�����a��ird��A{/w�/J/5/n/vA��A0���":t�/ C^/�/xZ/ ލ?���/��/1??���W���t�g��pE� ~1��?04�0
1�1@�IӀ��BµW�B]�NB2�(�A��@�u\�?����������b�0�|�uR�����
�>��ؽ��Bu�*C��$�)`��? ���G�C#���r�AU����1��eG���I�m�H�� I:��I�6[F����C4OI���J�:\IT��H
~QF�y��Ol@�*J�/� I8Y�I��?KFjʻC��-? �O�O__>_)_b_M_ �_�_�_�_�_�_�_o �_(oo%o^oIo�omo �o�o�o�o�o �o$ H3lW�{� ������2�� V�h�S���w�����ԏ �������.��R�=� v�a�������П���� ߟ��<�'�`�K�]� ��������ޯɯ��&�8�#�\��3(J��g�3:a������J�3��c4�������������1��㚅ڿ��1����e���14 �{ 2�2�r�`ϖτϺϨ�J�%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ��� �������3��W�B� {�f�4���������d�A����!��1�3� E�{�i��������������  2 Efn�7Fb�7��6�B�!�!� C9� �� �0@�/`r������#x��+=�3?, V�8�v��0�0�:�0�.
 D� ����//%/7/�I/[/m//�/�:� ���ֻ�G����$PARAM_M�ENU ?2���  �DEFPUL�SE�+	WAI�TTMOUT�+�RCV? S�HELL_WRK�.$CUR_ST�YL� 4<OP9TJJ?PTB_?Y2�C/?R_DECSN 0�Ű<�?�?�?�? �?OO?O:OLO^O�O��O�O�O�O�!SSR�EL_ID  �.�����EUSE_PROG %�*q%�O0_�CCCR0��B���#CW_HOSoT !�*!HT�_=ZT��O_�Sh_zQ��S�_<[_TIM�E
2�FXU� GD�EBUG�@�+�CG�INP_FLMS�Ko5iTRDo5gP+GAb` %l�tk�CHCo4hTYPE
�,� �O�O�o# 0Bkfx�� �������C� >�P�b���������ӏ Ώ�����(�:�c��^�p�����7eWOR�D ?	�+
 �	RSc`��P�NS��C4�JO�v1��TE�P��COL�է�2��gLVP 3�����Oj�TRACECTL� 1�2��!{ �� ��Қ�q�DT Q�2�Ǡ��D �� :��f��Ԡ�Ԡ���}�ׯ���;�4��4��4� ��;�u:�q:���;�U8�	8�
8�8�U8�8�8�8�T�@:�8�8����� ���ٱ޴���ؿ�$�6��� 
�l�~�@�R�dϞϰ� ��������
��V�h� zߌߞ߰��������� 
�,�>�P�*�<�v���*� +8� (
��)��*�������� ��)�;�M�_�q��� ������������ %,�>�P�b�t����� �������С�* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6@u bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� V�߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�?��?�1�$PGTR�ACELEN  ��1  ����0��6_U�P ����2A@�1@�1_CFG �ES�3�1
@�<D�0<DZO<C�0uO�$BDEFSPD ��/L�1�0���0H_CONFI�G �E�3 U�0�0d�D��2 �1�APpDsA�A��0��0IN'@T�RL �/MOA8lpEQPE�E��G��A<D�AIL�ID(C�/M	bTG�RP 1ýI �l�1B  ������1A�3�3FC� F8п E�� @eN	��A�AsA�Y�Y�A�@� 	 vO�Fg��_ ´8cokB ;`baBo,o>oxobo�o��1>о�?B�/�o�o~�o =?%<��
C @yd��"�������  Dz@�I�@A0�q� ��� ����ˏ���ڏ��� 7�"�4�m�X���|����Ú)ґ
V7.10beta1HF @�����Aq��Q m �?� �BܠPz�p �C��&�?B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@��8�f������ҡ�R9�ܣ�Rљ���1��i�������t<B!CeQKNOW_M  lE7FbT�SV ĽJ �BoC_�b�t�������@������1�]aSM�S]ŽK ���	NB~�0���Ŀ�K���-�bb ��A�RP����0��Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1�K
 4MU�iǨj� K�]�oߠߓ� �߷�������2��#� h�G�Y��}�����@��
������,�27�9I��1�<t�H���P3^�p�����,�4 ��������,�5(:,�6Wi{��,�7����,�8��!3,�MAD��6 F,�OVL/D  KD�xO�.�PARNUM � �MC/%�SCH� E
9'!G)�3Y%UPD/��E|�/P�_CMP_���0@�0'7E�$E_R_CHK�%5H�&�/�+RS���bQG_MO�+?=5_'?~O�_RES_G6��:�I�o�?�?�?�? O�?O7O*O[ONOO�rO�O�O�{4]��< �?�Oz5���O__|3  #_B_G_|3V b_�_ �_|3� �_�_�_|3�  �_�_o|3Oo>oCo|2V 1�:�k1!��@c?�=2THR_INRc0i!}�zo5d�fMASS�o� Z�gMN�o�cM�ON_QUEUE� �:�"�j0��*O�N� U1Nv�+�DpENDFqd?`yEcXEo`u� BEnp|PAsOPTIOMw�m;DpPROGRAoM %$z%Cp�}o(/BrTASK_�I��~OCFG ��$��K�DAkTA��T���j12/ď֏���� ��+�=�O�a������𩟻�͟��INFO
�͘��3t��!�3� E�W�i�{�������ï կ�����/�A�S��e�w�����Θ� �'��FJ�a K_N�q�T��˶ENBg Hڽw1��2��GN��2�ڻ P(�O�=���]ϸ��@���v� ��u�uɡdƷ_EDIT �T�����>G�WERFL�x�c�)�RGADJ �Ҷ�A�  $�?@j00��a�Dqձӆ5�?�����<u�)%e���Ș��FӨ�2�R��	�H;pl�G�b_�>��pAod�t$��*�/� **�:�j0�$�@�5 Y�T���^��q�߈b ~�L��\�n���� �����������4� F�t�j�|��������� ����bLBT �x����:� �$,�Pb� ��/����/ ~/(/:/h/^/p/�/�/ �/�/�/�/V? ??@? 6?H?�?l?~?�?�?�? .O�?�?OO O�ODO VO�OzO�O_�O�O�O �O�Or__._\_R_d_��_�_�_�_�_�_�f	 g�io�pWo�o{d�o��~o�ozoB�P?REF �Rږp��p
�IORI�TY�w[���MP�DSP�q��pwUT�6����ODUCT�3�����OG��_TG��8�����rTOENT 1�׶� (!AF_INE�p,�7�?!tcp7�_��!udN���!icmv��ޯrkXYK�ض���q�)� ,�����p��&�	��R�9�v� ]�o�����П����� �*��N�`�*�sK���9}�ߢ���Ư �,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE� �R��:�wd��连�2s�9Ks���PORT_NUUM�s�p����_CARTREP�{p�Ω�SKSTAv�w d�LGS)��ݶ��tӁpU�nothing��������{��TEMP ޾y��'e���_a_seiban�o\��olߒ� }߶ߡ���������"� ��X�C�|�g��� ����������	�B� -�f�Q���u������� ������,<b M�q��������(L�VE�RSIyp�w} �disabl�edWSAVE �߾z	260_0H768S?��!ؿ����/ !	5(�r)og+^/yÁe{/�/�/�/�/�*��,/? �p���_��p 1�Ћ�? �����Wh?xz?�W*pURGE��aB�p}vgu,�WF�0#DO�vƲ�vW%��4�(�C�WRUP_DELAY �\���5R_HOT �%Nf�q׿GO�5R_?NORMAL&H�rx6O�OZGSEMIjO��O�O(qQSKIPF3��W3x=_9 8_J_\_]�_�_{_�_ �_�_�_�_�_	o/oAo Soowoeo�o�o�o�o �o�o�o+=a Oq������ ��'��7�]�K���x����)E�$RA{����K/�zĀÁ_�PARAM�A3���K @.�@`\�61�2C<��y�M�C�6$�BÀ�BTIF�4`�RC_VTMOUu�cŻ�ÀDCRF3��I �+Q;�/�CC�SeD��#�1=h��-0�t]�/��ޅ�����1��0��_��k_����Cd;��.<�߈<�g�<?F+<L���Ѱ��d�u�L������� ϯ����)�;�M��_���RDIO_T?YPE  M=U��k�EFPOS1 ;1�\�
 x4/�����+�$/<�� $υ�pϩ�D���h��� ���'������o�
� ��.ߤ�Rߌ������ ��5���Y���i��*� <�v���r������� ��U�@�y����8��� \�����������?��xc����2 1�KԿX�T�x��3 1�����nY�S4 1�'9K�/�|'/�S5 1����/�/�/�/:/S6 1�Q/c/u/�/�-??Q?�/S7 1��/�/
?D?�?�?�?>d?S8 1�{?�?��?�?WOBO{O�?SM?ASK 1L�8�O�D�GXNO���Fx&�^��MOTEZ�hŻ��Q_ǁ�%]�pA݂��PL_RA�NG!Q]�_QOWE/R �ŵ�P1V�SM_DRYPR/G %ź%"O�_��UTART ���^�ZUME_PR�O�_�_4o��_EX�EC_ENB  yJ�e�GSPD`pO`WhՅjbTDBro�jRM�o�hING�VERSION �Ź#o�)I_AIRPURhP� �O(�MMT_ҡ@T�P#_ÀOB�OT_ISOLC��NTV@A'qhuN�AME�l��o�JO�B_ORD_NU�M ?�X#q�H768  �j1Zc@�r
��rV�s���r�?�r?��r�pÀPC_TI�MEu�a�xÀS2�32>R1�� �LTEACH PENDANw��:GX�!O �Maintena�nce Cons�j2����"��?No UseB�׏ ������1�C�y�V��NPO�P@�YQ��cS�CH_Lf`�%^ �	ő~��!UD1:�z��R�@VAIL�q�@�Ӏ�J�QSPA�CE1 2�ż ��YRs�i�@Ct��YRԀ'{��8�?��˯���� "���7�2�c�u����� G���߯ѿ򿵿�(� �u�AC�c�u����� Ͻ�߿���ϵ��(� �=�_�qσϕ�C߹� �����߱��$��9� [�m�ߑߣ�Q����� �߭��� ���	�W�i� {���M�������5� ��.S�e�w��� ��I������� *?as��E �����/&// ;/]o����� �/2/�/?"?�/7?Y/ k/}/�/�/O?�/�/�?��?�?O0OOKA�o�*SYPpM*��8.30261 �yB5/21/2018 A �WP�fG|�H�_TX`�� !$COMM�E�$US�Ap $EN�ABLEDԀ$sINN`QpIOR�B��@RY�E_SIG�N_�`�AP�AIT\�C�BWRK�BD<��_TYP�CRIN�DXS�@W�@%VF{RI{�_GRPԀ$UFRAM�r�SRTOOL\VMY�HOL�A$LE�NGTH_VTE�BTIRST�T ? $SECLP�X�UFINV_PO�S�@$MAR�GI�A$WAI�T�`�ZX2�\�VG-2�GG1�AI�@�S��Q	g�`_WR�BNO_USE_DI�B^uQ_REQ�BC�C�]S$CUR_T�CQP�R"a^f �G�P_STATUS>�A @ �A3`X�BLk�H$zc1�h��P@���@_�F�X �@E_MLoT_CT�CH_�J6�`CO�@OL�E�C�GQQ$W�@w��b#tDEADLO�CKuDELAY_CNT�a3qGt�a�$wf 2 �R1[1$X<�2*[2�{3[3$Zwy �q%Y�y�q%V�@�c�@��b$V�`�RV�UV�3oh>b�@ � q�d�0arMSKJ��LgWaZ�C`NRK�P�S_RATE�0�$���S
`�Q�TAC���PRD���e�SD*��a4�A�0�DG�A� 0�P�flp bquS2ppI�#`\
`�P 
�S\`�  �A�R_�ENBQ ��$RUNNER_SAXI�<`ALPL�Q��RU�THICQ�$FLIP7��DT�FEREN��R�IOF_CHSU�IW��%V)�G1����$P�řA�Q�Pݖ_J�F�PR_P�	�RV_DATA�A�  $�E�TIM���$VA�LU$�	�OP_ �  �A�  2 �S�C*�	� �$ITP_!�SQ]P�NPOU}�o�TOT�L�o�DSP��JO�GLIb��PE_P�Kpc�Of�i��PX�]PTAS�$KE?PT_MIR��¤2"`M�b�APq�aE�@�y�q�g@١c�vq�PG�BRK6��x���L�I��  �?�SJ�q�P�ADE�z�ܠBSOCz�M�OTNv�DUMM�Y16Ӂ$SV��`DE_OP��S�FSPD_OVR4
���@LD�����OR��TP8�LEb��F������OV��CSF��F����bF��d�ƣ&c)�fQc�LC�HDLY��REC�OV���`��W�PM��gŢ�RO�������_F�?� @v�S� �NVER�@�`O�FS�PC,�CSWD�ٱc�ձ���B����T�RG�š�`E_F�DO��MB_CM4}���B��BLQ�¢�	�Q�̄Vza�BUP��g��G
��AM����@`KՊ�e�_M�!�d�AMf�Q��T�$CA����DF����HBKd�v���I�OU��I'R��PA����������p���~��DVC_DB�S�!�x�Q�!�s�d�9�1�A��9�3A��AT�IO�0��͠��U0S����WaAB��R�+c�`tá`DؾA��_�AUXw�SUBCPUP���S�`�����3Եжc���3�FLyA�B�HW_Cwp�"�Ns&�]sAa��_$UNITS�M�>F�ATTRIz�Z�ެ�CYCL�CNE�CA���FLTR�_2_FI��TARTUPJp����Aƴ�LP������_S�CT*cF_F�F_P���b�FS��+�K�CHA/Q��*�d�RSD��Q�����Q���_TH�PRO8r���հEMPJ���rG�T� ��Q�DI�@y�RAOILAC/�bMX�CLOf�xS��ځ����拁���PR#�S�`app�C� {	��FUNC���RIN`QQP� �ԱRA)]R ���AƠ��AWAR�֓��BLZaWrA0kg�ngDAQ�B�rkLD�र&q��M�K���TI����j��$�@R�IA_SW��AF
��Pñ#��%%�p89r1��MOIQ���gDF_~P(�PD"�LM-�FA�PHR�DY�DORG�H�; _QP�s%MULCSE~Pz���*�� �J��Jײ��FAN_ALMLVG���!WRN�%HARDP��UcO�� K�2$SHADOW�]�kp�a02��� ST�Of�+�_^�w�AU�{`R��eP_SBR�z5���:F�� ��3MPINF?�p\�4��3REGV&/1DG�+cVm �C��CFL(��?�D�AiP���Z`�� �8����Z�	 �P(Q�$�A$Z�Q �V�@�[�
� ���EG��o���kAAR���㌵2�axG���AXE��ROB.��RED��W�QD�_�Mh�SYA��AF�:�FS�GWRI�P~F&�STR����E�˰EEH�)��D�a\2BkPB6P��=V��DvЗOTO�1)���ARYL�tR�v�3����FI&�ͣ$LI�NKb!\��Q�_�3S���E��QXY�Z2�Z5�VOFF����R�R�XxPB��ds�G�cFI�03g�������_J��'�ɲ�S�&qR0LTV[6���aT�Bja�"�bC���D�U�F7�TURB� X��e�Q�2XP�ЊgFL�E���x@��`�U9Z8���� +1	)�K��Mw��F�9��劂����OR!Qj��G;W3��� #�Ґd ���uz����1N�tOVE�q_�M�� ё?C�uEC�uKB�v'0 �x-�wH��t��� & `��qڠ�B�ё�u��q�wh�ECh����E)R��K	�EP�$���AT�K�6e9`e�W���AXs� '��v�/�R ��� �!�� ��P��`�@�`�3p�Yp�1�p �� �� �� (��  8�� H�� X�� h�� �x�� ������DEBU�$%3�I��·RAB���ٱ�s9V��� 
d�J� ����@񘧕������ �Q���a���a��3q���Yq+$�`%"<�cLA�B0b�u�'�GR�O���b<��B_ s��"Tҳ*`�0A�u�p�uq�p1}�ANDGp��������U��p1��  �ѷ0�Qθuݸ��P�NT0���SERsVE �Z@ $`�EAV�!�PO ����nP!�P@�$!�Y@  $.>�TRQ�b
=��B2G�K�%"2\��~� _  l���5�D6ERRVb(�I��V0`;���TOQ:�7�L�@
�R��e %G�%�Q�� <�50�F� ,�`�z��>�RA� 2� d!�����S�  M��pxU �����OCuG�  }��COUNT6Q���FZN_CFG�F� 4#��6��T�G4�_�=����(����VC ���M  �"��$6��q ��CFA E� &��X�@@�������A���r�AP��P@HEL�0~�� 5b`�B_BAS��RS)R�6�CSH��R��1�Ǌ�2��3��U4��5��6��7��98��}�ROO���̚P�PNLEA�cAB�)ë ��ACKu�IeNO�T��(B$UR08� =�_PU��!0��OU+�Pd�8j���� V��TPFWD_KAR��� ��RE(ĉ P�P�>7QUE�:RO�p�`r0P1I� x�j�Pp�f��6�QSEM���0��� A��STYfL�SO j�DIX��&�����S!_TM>CMANRQ��P�ENDIt$KEYSWITCH��ذ�kHE�`BE�ATM83PE{@L�E��>]��U��F���SpDO_H�OM# O�@�EF�pPRaB�A#PY��C� O�!���OV�_M|b<0 IOCqM�dFQ��h�;HKYA D�Q�7��UF2��M���p޸cFORC�3WA�R�"�OM|@ G @S�#o0U)SUP�@1�2&3&Q4E���T�O��L�y��8UNLOv��D4K$EDU1  ��SY�HDDN�F� M�BLO�B  p�SN�PX_AS�� �0@�0��81$S{IZ�1$VA{�~��MULTIP-���# A� � $��� /4`��BS��0�C���&F'RIFBO�S����3� NF�ODBUP߰�%@3;9(���܋�Z@ x��SI���TEs�r�cSG%L�1T�Rp&�Н3xB��@�0STMTq2�3Pg@VBW�p�4�SHOW�5@�SmV��_G�� 3p�$PCJ�PИ���F�B�PHSP A�W�EP@VD�0WC�� ���A00 ��PB XG XG XGT$ XG5VI6VI7VIU8VI9VIAVIBVI@�XG�YF�0XGFVH���XbI1oI1|I1��I1�I1�I1�I1��I1�I1�I1�I1��I1�I1Y1Y2�UI2bI2oI2|I2�I2�I�`�X�I2p�X��I2�I2�I2�I2
�I2Y2Y�p�hbIU3oI3|I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3�IU3Y3Y4�i4bIU4oI4|I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4�IU4Y4Y5�i5bIU5oI5|I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5�IU5Y5Y6�i6bIU6oI6|I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6�IU6Y6Y7�i7bIU7oI7|I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7�I�7Y7T��VP� UD�y"ՠ��Q
<A62��t��R��CMD� ��Mb5�Rv�]��Q_hЁR���e����<�Y�SL���  � �%\2��+4�'��xW�BVALU���b��'���FH�ID�_L���HI��I���LE_��㴦��$0C�SAC��! h �VE_BLCK��1>%�D_CPU5ɧ  5ɛ �����C�� ���R " � �PWj��#0��LA��1SBћì���R?UN_FLG�Ś� ���ĳ ���������šH���Хą�T�BC2��# � @ B��e �S�88=�FTDC�����V���3d�Q�TH�F�����R�L�ESERVE9��F���3�2�E��Н��X -$��LEN`9��F��f�RA��LW"G�W_5�b�1�њд2�MO-�T%S60U�Ik�0�ܱF�����[�DEk�21LA3CEi0�CCS#0�� _MA� j��z玤�TCV����z�T �������.Bi�'A�$z�'AJh�#EM5���J��@@i�V�z���2Q �0&@o�h��JK��VK9��{����щ�J0����J�J��JJ��AAL����������4��5�ӕ N1������J.�LD�_�1* v�CF�"% `�GROU���1�A�N4�C�#m REQ�UIR��EBU��#��6�$Tk�2�$���zя #�&{ \�APPR� �C� 0�
$OPE=N�CLOS��St��	i�
��&' �MfЩ���W"N-_MG�7CB@��A���BBRK�@NOLD@�0RTMO_5ӆp1	J��P�����@���������6��1�@ )!�#�(� ������'��+#PATH ''@!6#@!�<#� � 9'��1SCA��l�6IN��UCJ�[1� C0@UM�(Y  ��#�"�����*���*���� PAYLOA�~J2LؠR_A	N^�3L��91�)�1AR_F2LSHg2B4LO4�!F7��#T7�#ACRL_@�%�0�'�$��H���.�$HA�2FL�EX��J!�) P�2�D߽߫��|�0��* :�� ��z�FG]D����z���%�F1]A�E�G4�@F�X�j�|���BE�� �����������(� �X�T*�A���@�XI��[�m�\At�T$g�QX <�=��2TX���emX �������������������+	�J>+ �-�K]o|�٠cAT�F�4�ELFP�Ѫs�J� *� J�EmCTR�!�AT�N�vzHAND_VB.��1��$7, $8`F2Avԍ��SWu	#-?� $$M*0. �]W�lg��PZ����A��� 1����:QAK��]AkAzP��LN�]DkDzePZ G��C�ST_hK�lK�N}DY�� � A����0��<7]A <7W1�'��d�@g`�P�������t"
"J"�. M��2D%"��H����AS�YMj%0�� j&-��-W1�/_�{8�  �$�����/�/�/�/ 3J<�:9�/�89.�D_VI�v��>��V_UNI�ӛ��cD1J����╴�W< ��n5Ŵ�w=4��9���?�?<�uc�4�3{d�%�H���/��j��0�DIzuO��w�k�>0 �`��I��A��#�� �@ģ���@��IPl� 1 � /�ME.Qp��9�ơT}�PT�;pG �+ Gt� ���'���T�0 $D�UMMY1��$�PS_�@RF�@ � G b�'FLA�@ YP(c|��$GLB_TP�ŗ����9 P�q��2 �X� z!ST9�� SBRM M21�_V�T$SV_�ER*0O�p����C)L����AGPO��f��GL~�EW>�3 �4H �$YrZBrW@�x�A1+�A���"	""�U&�4 �8`NZ�"�$GIn�p}$&� -�8 �Y�>�5 LH {��}$F�E��NWEAR(PN�CF��%PTANC�B	!JsOG�@� 6.@$JOINTwa�?pd�MSET>�7�  x�E��HQtpS�{r��up>�8� ��pU.Q?�� L?OCK_FOV06�ޅ�BGLV�sGL�t�TEST_XM�� 3�EMP��8���_�$U&@%�Fw`24� Y��5��h2�d��3��CE- |���� $KAR�Q}M��TPDRA)�����VECn@��kIU��6��HEf�OTOOL�C2V�D;RE IS3ER96��@ACH� �7?Ox �Q�29�Z�H I�  @�$RAIL_BO�XEwa�ROB�O��?��HOW�WAR�1�_�zROLMj��:qw�pjq� �@ O_Fkp�! d�l>�9��� �R O8B:� �@�c�OU�;�Һ�3ơ�r�q�_�$PIP��N &`H�l�@��#@?CORDEDd�p �>f�fpO�� <o D ��OB� �sd���Kӕ����qSYS�ADR��qf��TCHt� o= ,8`ENo�*�1Ak�_{�-$Cq�,Be�VWVA��> �  &��PREV_RT$EDITr&V/SHWRkq�֑ �&R:�v�D��JA��$�a$HEAD��6�� �z#KE|:�E�CPSPD�&�JMP�L~��0R�*P��?��1%&Ij��S�rC�pNE; <�q�wTICK�C���M�13�3HN���@ @� 1Gu�!_�GPp6��0STY'"xLO��:�2l2�?�A t 
m G�3%%$R!{�=��S�`!$��w`��������Pˠp6SQU���E��u�TERC��0��TSUtB ����hw&`gw�Q�)�pO����@IZh��{��^�PR�0kюB1XPU���Eg_DO��, XS�K~�AXI�@���UR�pGS�r� ^0��&��p_) �ET��BPm��o��0Fdo��0A|���R�h���a;�SR�Cl>@P��b_� yUr��Y��yU��yS�� yS���UЇ�U���U�� �U�]��Ul[��Y�bXk�]Cm������ 1@SC�� 7D h�DS~0��fQ�SP���eATހ��A]0,2N�AD�DRES<B} S�HIF{s��_2C�H�p�I��=q�+TVsrI��E"����a�Ce�
��
;�V8W�A��F \��qA��0l|\A@�rC��_B"R{zp�ҩq�T�XSCREE�Gzv��1TINA����t{����A�b?�H T1�ЂB��р��I��A��BE�y RRO������ B��Dv��UE4I �g��!p�S��RSM<]0�GUNEX(@~���j�S_S�ӆ��Á։񇣣�ACY�0�o 2H�pUE;��J�����@GMTJ��Lֱ�A��O	�/BBL_| W8��ЧK ��0s�OM���LE/r��� TO�!�s�RIGH��B�RD
�%qCKGR8л�TEX�@����WIDTH�� �Bh[�|�<��I_��}Hi� L 8K�B��_�!=r���R:�@_��Yґ��O6qJ�Mg0紐U��rh�Rm��LUMh��FpERVw �QP���`�N��&�/GEUR��FP)�M)� LP��(RE%@�a)ק�a�!��f ��5�6�7�8 Ǣ#B�É@���tP�f�W�S@M�U{SR&�O <�����U�Qs�FOC\)��PRI;Qm� �:���TRIP�Om�UN����Pv��0��f%��'���@��0 Q����AG �0T� �a>q�OS�%�RPo���8�R/�A�H�L4$����U¡�SU�g�p�¢5��OFF���T�}�O�� G1R�����S�GUN��6�B�_SUB?���,�SRTN�`TUg2���mCOR| D�RAU�rPE�TZ�#'�VC�C��	3V AC?36MFB1f$c�{PG �W (#�.�ASTEM����L�0PE��T3G��X �\ ��MOV1Ez�<���AN�� ����M���LIM_X��2��2��7�,������ı�
��VF@�`E�� }��04Y�F�IB�7���5S���_Rp� 2��� WİGp+@��}���P��3�Zx ���3���A�rݠCZ�DRID�����Vy08�90� D~e�MY_UBYd�@��6��@��!��X��P_S��3��mL�KBM,�$+07DEY(#EX`������UM_MU� X����ȀUS�� �z��G0`PACI�� �а@��:��:,�:����RE/�3qL�+���:[��TA�RG��P�r��R<�\ d`��A���$�	��AR��SWH2 ��-��@Oz��%qA7p�yREU�Uh�01�,�HK�2]g0�qP� N�� �EAM0GWORx���MRCV3�W^ ���O�0M��C�s	���|�REF_���x(�+T � ���������3_RCH4(a �P�І�hrj�NA�5��0�_ ��2����L@4��n�@@OU~7w�6���Z��a2[ư�RE�p�@;0\��c�a'2K�@SUL���]��C��0�^��� NT��L�3��@(6I�(6q�(3� L��@Q5��Q5I�]7q�}�)Tg`4D`�0.`0ПAP_HUC�5S]A��CMPz�F�6(�5�5�0_�aR��a��1I\!X�9|"GF}S��ad ��qM��0p�UF_x�0�B� �ʼ,RO��Q���'����UR�3GR�`.�3IDp���)�D�;��A��~�IEN��H{D���V@A J���S͓UWm�i=�����TYLO�*�5�$����bot +�cPA�{ �cCACH� vR�UvQ��Y��p�#�CF�I0sFR�XT8���Vn+$HO����P!A3�XBf�(01 ���$�`VPy� �^b_SZ313he6K3he12J�eh chlG�chWA�UMP�j���IMG9uPAyD�iiIMRE�$^�b_SIZ�$P�����0 ��ASYNB{UF��VRTD)u�5tqΓOLE_2�DJ�Qu5R��C��U���vPQuECCUlVEMV �U�r��WVIRC�aIuVTPG���rv1s���5qMPLAqa��v쨣��0�cm� C/KLAS�	�Q�"��d  �ѧ%ӑӠ�@}¾�R���Ue A|�0!�rSr�T�# 0! �r�iI��ml�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f �� >֦3�@Sp�SgLOW>�RO��ACCE���!� 9��VR�#���p:���A1D�����PAV�j��� D����M_B8"���^�JMPG ���g:�#E$SSC@��x&�vPq��hݲ�vQS�`qVN��L;EXc�i T`�s�r���Q�FLD �DEsFI�3�0p2���:��VP2�V�j� �A��V|�4[`MV_PIs���t���A�@��F	I��|�Z��Ȥ����`�A���A��~�GAߥ�1 LOO��1 JC�B���Xc��^`�#P�LANE��R��1F@�c�����pr�M� [`�噴��S����f� ���Af��R�Aw�״t9U��pRKE��d�VANC�A���� k���ϲ�BwR_AA� l���2� ��p�#��m h���O K�$����2��kЍ0OU&A�"eA�
p�pSK�T�M@FVIEM 2l� ��P=���n �<<��dK�UMM�YK1P��`D6�ȟ�CU��#A�U��o $��T�IT�$PR�����OP���V�SHIF�r�p`J�Qsԙ�fOxE[$� _R�`U�# ����s��q������ G�"G�޵'�T�$��SCO{D7�CNT Q i�l�>a�-�a�;� a�H�a�V���1�+�2u1��D���� w � SMO�U�q��a�JQ���%��a_�R[�r�n׍*@LIQ�AA/`��XVR��s�n�T�L���ZABC��t�t�c�
��Z�IP��u���LV�bcLn"���MPkCFx�v:�$��� ���DMY_L�N�������@y�w �Ђ(a�u� MCM��@CbcCART_��DPN� $J71D��=N�Gg0Sg0�BUXW|� ��UXEUL|ByX���	��L�Z��x �	���m�YH�D>b  y 80�֞�0EIGH�3n�?�(� H����$z� ���|�����$B� Kd'��_��L3��RVS�F`���OVC�2'�$|�>PD&��
q���5D��TR�@ �Vc��SsPHX��!{ ,� �*<�$R�B2 2 ���C!��  ���V+L�b*c%Rg!`+g"�`V*~�,8�?�V+ �/V.�/�/?�/�/V(7%3@/R/d/v/�/6? �/�/�?�?�?O4OOION;4]?o?�?�?�? SO�?�?�O_�O0_Q_8_f_N;5zO�O�O�O �Op_�O_o8o�_MonoUo�oN;6�_�_�_ �_�_�oo%o4U j�r�N;7�o�o �o�o�o� BQ�r�@5���������N;8� ����Ǐ=�_�n����R���ş��ڟN;Gw � џ
�
������W� i�{�������ï�.��������A��d W�<�N�|�������Ŀ ֿ�ޯ���0�B� _�R�d�꿤϶����� ��������*�L�^� �rτ�
��������� ���&�8�J�l�~�w `ҟ @�Ѐ�����ߩ��-� ���&�,���9�{� ����a����������� ����A'Y� ������� �a#1�
���N;_MODE  y��S ��[�Y�B���
/�\/*	|/�/R4CW�ORK_AD�	��
�T1R  ����� �/� _I�NTVAL�+$���R_OPTIO�N6 �q@V�_DATA_GR�P 27���D��P�/~?�/�?�9� �?�?�?�?OO;O)O KOMO_O�O�O�O�O�O �O_�O_7_%_[_I_ _m_�_�_�_�_�_�_ �_!ooEo3oioWoyo �o�o�o�o�o�o�o /eS�w� ������+�� O�=�s�a�������͏ ���ߏ��9�'�I��o�]�����$SA�F_DO_PUL�S� �~������C?AN_TIM�����ΑR ��Ƙ�"��5�;#U!P"�1!��� �?E�W�i� {�����.�ïկ���X��'(~�T"2F���dR�I�Y��2�o+@a얿�����)�u��� k0ϴ���_ ��  �T� � �2�D�)�T D��Q�zό� �ϰ���������
�� .�@�R�d�v߈ߚ�/<V凷������߽��R�;��o �W�p��
�?t��Diz$�~ �0 � �T" 1!�������� ����������*�<� N�`�r����������� ����&8J\ n���������"4FX �� ࿁������ �/`4�=/O/a/s/ �/�/�/�/�/�/�!!/ �0޲k�ݵu�0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ ok $o6oHoZolo~o�o�o �o�o1/�o�o 2 DVhz�/5?�� ������&�8� J�\�n���������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u��� ���`Ò�ϯ ����)�;�M�_� q���������˿ݿ�� ����3� ����&2,��	12345678v��h!B!�U�2�Ch���0� �ϵ����������!� 3�9ѻ�\�n߀ߒߤ� �����������"�4� F�X�j�|�h�K߰��� ������
��.�@�R� d�v������������� ��*<N`r ������� &��J\n�� ������/"/ 4/F/X/j/|/;�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �/�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_�?L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o=_�o �o�o�o�o�o 2 DVhz�����h������u�o�.�@�R���Cz � B��   ����2&� � �_�
���  	�_�2�Տ���,�_�p������ďi�{�������ß ՟�����/�A�S� e�w���������N�� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�_�����<v�_��$SC�R_GRP 1
�� �� �t ��� ���	 ��������� �������_�����Ϝ)�a����&�DE� DW8���l��&�G�CR-3�5iA 9012�34567890���M-20��8~��CR35 ��F:�
��������������:֦�Ӧ��G���&������	���]�o����:���H���>�����������&���ݯ:��j����g�X�����B�t�����������A����  1@�`��@� (' ?�=��Ht�P�
��F@ F�`z�y����� � �$H���Gs^p��B� �7��/�0// -/f/Q/�/u/�/�/�/�8���P�� 7%?�����"?W?-2?<���]? H�1�?t�ȭ7�������?-4A, �&E@�<�I@G�B-1 3OZOlO-:HA�H�O�O.|O P�B(�B�O��O_��EL_DE�FAULT  ~����`�SHOTSTR�#]A7RMIPOWERFL  i�z/UYTWFDO$V� /URRVENT 1�����NU L!DU�M_EIP_-8��j!AF_IN�E#P�_-4!FT$�_->�_;o!��`o� �*o�o!RPC_MAIN�o�jh�vo�o�cVIS�oii��o!TMPpPU�Yd�k!
PMON_�PROXYl�Ve Z�2r��]f���!RDM_SR�V��Yg�O�!�R��k��Xh>���!%
�`M��\i����!RLSYNC��-98֏3�!gROS�_-<�4"���!
CE4pMT'COM���Vkn�˟{!	��CONS̟��Wl���!��WOASRC��Vm�vc�!��USBd��XnR���Noӯ��� ����!��E��i�0����WRVICE_�KL ?%�[ �(%SVCPR#G1��-:Ƶ2ܿ�"˰3�	�˰4,�1�"˰5T�Y�˰6|ρ�˰7�ϩ�˰�����	9����ȴf�!�˱ οI�˱��q�˱ϙ� ˱F���˱n���˱�� �˱��9�˱��a�˱ ߉��7߱��_��� �����)���� Q����y��'��� O����w����� ����˰��İd �c������ =(as^�� ����/�/9/ $/]/H/�/l/�/�/�/ �/�/�/�/#??G?2? k?V?}?�?�?�?�?�? �?O�?1OCO.OgORO �OvO�O�O�O�O�O	_��O-_��_DEV ��Y�MC�:5Xd�GTG�RP 2SVK ���bx 	� 
+ ,�PK 5_�_ �T�_�_�_o�_'o9o  o]oDo�ohozo�o�o �o�o�o�o5{�_ g������ ����?�&�c�u� \�������Ϗ���J \)���M�4�q���j� ����˟ݟğ��%� ��[�B��f����� �ٯ�������3�� W�i�P���t���ÿ�� �ο���A�(�e� L�ί��RϿ��ϸ��� ��� ��O�6�s�Z� �ߩߐ��ߴ������ '�~ϐ�]���h�� ������������5� �Y�@�R���v����� ����@�	��?& cu\����� ���;M4q X�������/ �%//I/[/B//f/ �/�/�/�/�/�/�/�/ 3??W?�L?�?D?�? �?�?�?�?O�?/OAO (OeOLO�O�O�O�O�O��O�O�O_iV �N�Ly�6 * �		S=>��+�c"_VU@Tn_Y_B����B�2�J�j~Q´~_g_�_��Q%JOGGI�NG�_�^7T(?Vj�Z�Rf��Y���/e�_%o7e�Tt�]/o�o{m�_�o�m ?Qi�o�o;)Kq%��o�}os ������9�{ `��)���%���ɏ�� �ۏ�S�8�w��k� Y���}���ş���+� �O�ٟC�1�g�U��� y�������'���� 	�?�-�c�Q���ɯ�� ��w���s����;� )�_ϡ���ſOϹϧ� ��������7�y�^� ��'ߑ�ߵߣ����� ���Q�6�u���i�W� ��{������=�� M���A�/�e�S���w� ����������� =+aO������ u���9' ]���M��� ���/5/w\/� %/�/}/�/�/�/�/�/ =/"?4?�/?�/U?�? y?�?�?�??�?9?�? -OO=O?OQO�OuO�O �?�OO�O_�O)__ 9_;_M_�_�O�_�Os_ �_�_o�_%oo5o�_ �_�o�_[o�o�o�o�o �o�o!coH�o{ ������;  �_�S�A�w�e��� ����я���7���+� �O�=�s�a������ П�����'��K� 9�o�������_���[� ɯ���#��G���n� ��7���������ſ�� ��a�Fυ��y�g� �ϋϭϯ�����9�� ]���Q�?�u�cߙ߇� ����%���5���)�� M�;�q�_���߼��� �������%��I�7� m������]������� ����!E��l�� 5������� _D�we� ����%
//� ��=/s/a/�/�/�/ ��/!/�/??%?'? 9?o?]?�?�/�?�/�? �?�?O�?!O#O5OkO �?�O�?[O�O�O�O�O _�O_sO�Oj_�OC_ �_�_�_�_�_�_	oK_ 0oo_�_co�_so�o�o �o�o�o#oGo�o; )_Mo����o ����7�%�[� I�k���������� ُ���3�!�W���~� ��G�i�C����՟� ��/�q�V������w� �������ѯ�I�.� m���a�O���s����� ��߿!��E�Ͽ9�'� ]�Kρ�oϑ����� Ϸ����5�#�Y�G� }߿Ϥ���m���i��� ���1��U��|�� E���������	��� -�o�T������u��� ��������G�,k� ��_M�q��� ����%[ Im���	� ��//!/W/E/{/ ��/�k/�/�/�/�/ 	???S?�/z?�/C? �?�?�?�?�?�?O[? �?RO�?+O�OsO�O�O �O�O�O3O_WO�OK_ �O[_�_o_�_�_�__ �_/_�_#ooGo5oWo }oko�o�_�oo�o�o �oC1Sy�o ��oi����� 	�?��f�x�/�Q�+� ��Ϗ�����Y�>� }��q�_�������˟ ���1��U�ߟI�7� m�[�}����ǯ	�� -���!��E�3�i�W� y�ϯ��ƿ������ ��A�/�eϧ���˿ UϿ�Q��������� =��dߣ�-ߗ߅߻� ���������W�<�{� �o�]������� ��/��S���G�5�k� Y���}����������� ����C1gU� �����{���� 	?-c���S ������/;/ }b/�+/�/�/�/�/ �/�/�/C/i/:?y/? m?[?�??�?�?�??  O??�?3O�?COiOWO �O{O�O�?�OO�O_ �O/__?_e_S_�_�O �_�Oy_�_�_o�_+o o;oao�_�o�_Qo�o �o�o�o�o'ioN `9���� ��A&�e�Y�G� i�k�}�����׏��� =�Ǐ1��U�C�e�g� y����֟���	��� -��Q�?�a���ݟ�� ퟇��ϯ��)�� M���t���=���9��� ݿ˿��%�g�Lϋ� ��mϣϑϳ����� ��?�$�c���W�E�{� iߟߍ߯������;� ��/��S�A�w�e�� �����������+� �O�=�s������c� ����������'K ��r��;���� ���#eJ� }k�����+ Q"/a�U/C/y/g/ �/�/�//�/'/�/? �/+?Q???u?c?�?�/ �?�/�?�?�?OO'O MO;OqO�?�O�?aO�O �O�O�O__#_I_�O p_�O9_�_�_�_�_�_ �_oQ_6oHo�_!o�_ io�o�o�o�o�o)o Mo�oA/QSe�����%{,p��$SERV_MA_IL  +u!���+q�OUTPU]T�$�@��RV 2�v  $� (�q�}���SAVE7�(�TO�P10 2W�� d 6 *_�π(_������ #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽݷ毅YP��'�FZN_CFG �u'$�~����?GRP 2�D�� ,B   A�[�+qD;� B�\��  B4~��RB21��HELL��u��j��k�2�����%RSR�������
�C� .�g�Rߋ�v߈��߬߀����	���-�?�Q�_�  �_�%Q���_���,p�����ޖ�g�2�,pd����HK ;1�� ��E� @�R�d����������� ������*<e�`r���OMM ������FTOV_ENB�_����HOW_REG_�UI�(�IMIO/FWDL� �^�^)WAIT���$V1�^�NT�IM���V�A�_)_UNI�T����LCT�RYB�
�MB�_HDDN 2W� 2�:%0  �pQ/�qL/^/�/�/�/��/�/�/�/�"!ON�_ALIAS ?5e�	f�he�A? S?e?w?�:/?�?�?�? �?�?OO&O8OJO�? nO�O�O�O�OaO�O�O �O_"_�OF_X_j_|_ '_�_�_�_�_�_�_o o0oBoTo�_xo�o�o �o�oko�o�o, �oPbt�1�� �����(�:�L� ^�	���������ʏu� � ��$�Ϗ5�Z�l� ~���;���Ɵ؟��� �� �2�D�V�h���� ����¯ԯ���
�� .�ٯR�d�v�����E� ��п���ϱ�*�<� N�`�r�ϖϨϺ��� w�����&�8���\� n߀ߒߤ�O������� ����4�F�X�j�|� '����������� �0�B���f�x����� ��Y��������� >Pbt��� ���(:L �p����c� � //$/�H/Z/l/ ~/)/�/�/�/�/�/�/�? ?2?D?V?]3�$�SMON_DEF�PRO ����1 �*SYSTE�M*0m6REC�ALL ?}9� ( �}8co�py frs:o�rderfil.�dat virt�:\tmpbac�k\=>147.�87.149.4�0:2896  >�815172]?O�+M}/�2mdb:*.*�?�?�?O�Ol�O7D3x�4:\HO �@ZOu@sO�O_(_;@4�Ea�O�OpE�O_��_�_ }
xyz�rate 61 �J_\_n_�_o#o6E�W�_44 �_�_o �o�o�_Jo\ono�od#6E?o�f02�`@�o�o��9B9�?��?I[qy
��/L0 ?O�Rz������8\�H_�_Vvt����)� }5?_Џ������ ����X�s����(� ;�֟_��������� L�^���$�7�ȯ گm���������ǟP� �}�� �3�E��i� ���Ϟϱ�ïV��y� 
��/�A���e���+� �߭o�_Q�c�u߇��8*�=Oy192^~�� �����mY�k�}��� �3oE�0:9308 ����������8C�3L�outpu�t\tcpser�v3.pcC�: �over =>3�70278p@357235w���� ��ѿI�[�����/O A�\T�o�$�O ���X����;_ L^[�t�/)/�� ������/�/�/:L ���/?%?���/ � ?�?�?6��l ~?O!O���?��? �O�O�/�/M?�/zO_ _0?B?�Of?�O�_�_ �?�?SO�?v_�_o�_ >O�_�_�_o�o�o�O �OW_r_�o':_�o�^_�o�����$�SNPX_ASG 2����q�� P �0 '%R[1]@1.1��y?��s%�!�� E�(�:�{�^������� Տ��ʏ���A�$� e�H�Z���~���џ�� ��؟�+��5�a�D� ��h�z�����ů�ԯ ���
�K�.�U���d� ������ۿ������ 5��*�k�N�uϡτ� �ϨϺ������1�� U�8�Jߋ�nߕ��ߤ� ���������%�Q�4� u�X�j�������� �����;��E�q�T� ��x����������� %[>e�t ������! E(:{^��� ���/�/A/$/ e/H/Z/�/~/�/�/�/ �/�/�/+??5?a?D? �?h?z?�?�?�?�?�? O�?
OKO.OUO�OdO �O�O�O�O�O�O_�O 5__*_k_N_u_�_�_ �_�_�_�_�_o1oo Uo8oJo�ono�o�o�d��tPARAM ��u�q ��	��jP�d9p��ht��pOFT�_KB_CFG � �c�u�sOPI�N_SIM  �{vn��p�p�RVQSTP_DSBW~r"t�Ht�SR Zy �� &!pINGS� EL_5SEM����vTOP_�ON_ERR  �uCy8�PTN �Zuk�uA4�R�_PR��D��`VCNT_�GP 2Zuq�!px 	r��ɍ����׏��wVD��ROP 1�i p� y��K�]�o������� ��ɟ۟����#�5� G�Y���}�������ů ׯ�����F�C�U� g�y���������ӿ� �	��-�?�Q�c�u� �ϙϫ���������� �)�;�M�_�qߘߕ� �߹���������%� 7�^�[�m����� ��������$�!�3�E� W�i�{����������� ����/ASe w������� +=Ovs� ������// </9/K/]/o/�/�/�/ �/�/�/?�/?#?5? G?Y?k?}?�?�?�?�?��?�?�?OO)�PRG_COUNT8v��k�GuKBENBĀ�FEMpC:t}O_U�PD 1�{T  
4Or�O�O�O __!_3_\_W_i_{_ �_�_�_�_�_�_�_o 4o/oAoSo|owo�o�o �o�o�o�o+ TOas���� ����,�'�9�K� t�o���������ɏۏ ����#�L�G�Y�k� ��������ܟן��� $��1�C�l�g�y��� ������ӯ����	�� D�?�Q�c��������� ԿϿ����)�;��d�_�q�=L_INF�O 1�E-�@ �2@����������� �ٽ`y�*�d�h'���¬��=`�y;MYSDEBU)GU@�@���d�If�SP_PASSUE�B?x�LOG � ���C���*ؑ�  ��A��?UD1:\�Ԙ���_MPC�ݵE&�$8�A��V� �A�?SAV !��������X���SV�Z�TEM_TIM�E 1"���@� 0  �X��X�X����$T1SVGUNS�@�VE'�E��AS�K_OPTION�U@�E�A�A+�_D�I��qOG�BC2_?GRP 2#�I�������@�  C����<Ko�CFG %z��� �����`��	�.> dO�s���� ���*N9r ]������� /�8/#/\/n/��Z+ �/Z/�/�/H/�/?�/ '??K?]�k?=�@0s? �?�?�?�?�?�?O�? OO)O_OMO�OqO�O �O�O�O�O_�O%__ I_7_m_[_}__�_�_ �X� �_�_oo/o�_ SoAoco�owo�o�o�o �o�o�o=+M Oa������ ���9�'�]�K��� o���������ɏ��� #��_;�M�k�}���� ����ß�ן��1� ��U�C�y�g������� ��������	�?�-� c�Q�s���������� Ͽ����)�_�M� ��9��ϭ�������m� ��#�I�7�m�ߑ� _ߵߣ���������� �!�W�E�{�i��� �����������A� /�e�S�u�w������� ������+=O�� sa������ �9']Km o������� #//3/Y/G/}/k/�/ �/�/�/�/�/�/?? C?��[?m?�?�?�?-? �?�?�?	O�?-O?OQO OuOcO�O�O�O�O�O �O�O__;_)___M_ �_q_�_�_�_�_�_o �_%oo5o7oIoomo �oY?�o�o�o�o�o 3!CiW��� ������-� /�A�w�e��������� �я���=�+�a� O���s�������ߟ͟ ��o�-�K�]�o�� ������ɯ���צ���$TBCSG_�GRP 2&ץ��  ��� 
 ?�  6�H�2�l�V���z����ƿ�������(~�d�E+��?�	 HC���>���G����?C�  A�.�e��q�C��>ǳ33D��S�/]϶�Y��=���� C\  B����B���>�̱��P���B�Y�zD��L�H�0�$��@��J�\�n�����@� Ҿ���������=�Z�`%�7����?3������	V3.�00.�	cr35��	*����
�`������� 3�|�4�   {��CT�v�}��J2��)������CFoG +ץ'�Y *������I�9���. <
�<bM�q� ������( L7p[��� ���/�6/!/Z/ E/W/�/{/�/�/�/�/ .�H��/??�/L?7? \?�?m?�?�?�?�?�?  OO$O�?HO3OlOWO |O�O����Oӯ�O�O �O!__E_3_i_W_�_ {_�_�_�_�_�_o�_ /oo?oAoSo�owo�o �o�o�o�o�o+ O=s�E���Y �����9�'�]� K�m�������u�Ǐɏ ۏ���5�G�Y�k�%� ��}�����ßşן� ��1��U�C�y�g��� ����ӯ������	� +�-�?�u�c������� ���Ͽ���/�A� S�����qϓϕϧ��� �����%�7�I�[�� �mߣߑ߳������� ���3�!�W�E�{�i� ������������ �A�/�e�S�u����� ���������� +aO�s��e� ����'K9 o]����� ��#//G/5/k/}/ �/�/[/�/�/�/�/�/ ??C?1?g?U?�?y? �?�?�?�?�?	O�?-O OQO?OaO�OuO�O�O �O�O�O�O___M_ �e_w_�_3_�_�_�_ �_�_oo7o%o[omo o�oOo�o�o�o�o�o !3�o�oiW� {������� /��S�A�w�e����� ��я�������=� +�M�s�a��������� ߟ�_	���_ן]� K���o�������ۯɯ ���#���Y�G�}� k�����ſ׿����� ���U�C�y�gϝ� ���ϯ��������	� ?�-�c�Q�s�u߇߽� ���������)��9� _�M����/����i� ������%��I�7�m� [��������������� ����EWi{5 �������� A/eS�w� ����/�+// O/=/_/a/s/�/�/�/ �/�/�/?'?��??Q? c??�?�?�?�?�?�? �?O�?5OGOYOkO)O��O}O�O�O�O�N  9�@S V_�R�$TBJOP_GRP 2,�E��  �?�V	-R4S.�;\��@|�u0{SPU >y��UT @�@�LR	 �C� ��Vf  C���xULQLQ>�33�UN�R����U�Y?�@�=�ZC��P���ͥR��P  �B��W$o/gC���@g�dDb��^���eeao�P&�ff�e=�7LC/kaB o�o�P���P�efb-C�p��^g`�d�o�P�L�Pt<�eVC�\  �Q@�'p�>`�  A�oL�`�_wC�BrD�S�^�]�_�S�`?<PB��P�anaa`C�;�`L�w�aQoxp�x~�p:��XB$'tMP@�PCHS��n���=�P����trd<M�gE�2pb� ���X�	��1��)� W���c���������� ��󟭟7�Q�;�I�(w���;d�Vɡ�U	V3.00RS�cr35QT*��QT�A�� �E�'E�i��FV#F"wq�F>��FZ� �Fv�RF�~M�F���F����F��=F����F�ъF��3�F���F�{�G
Gd�G�G#
��D��E'�
EMKE����E�ɑE����E��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF�u��<#�
<t%���ٵ=�_�:�V �R�p��V9� ]ESTPA�Rtp�HFP*SHR�\�ABLE 1/�;[%�SG�� (�W�G�G�G� WTQG�	G�
G�G�T��QG�G�GȜܱv�RDI~�EQ��ϧϹ�������W�O _�q�{ߍߟ߱���w�	S]�CS !ڄ��� ����������&�8� J�\�n����������� �� ]\�`��	�� (�:�����
��.�@��w�NUM  V�EEQ�P	P� ۰ܰw�_CFG� 0��)r-PIMEBF_TTb�p�CSo�,VERڳ�-B,R 11�;[ 8��Rd�@� �@&  � ������// )/;/M/_/q/�/�/�/ �/�/?�/?J?%?7? M?[?m?>�@�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_�y_�_�_l_�Y@�cY�MI_CH�AN8 c cDOBGLV��:c�X�	`ETHERA�D ?f�\`��?�_uo�oQ�	`oROUTV!	
�!�d�o�lSNM�ASKQhcba255.uߣ'9�ߣY�OOLOFS�_DIb��U;iO�RQCTRL I2		�Ϸ~T� ����#�5�G�Y� k�}�������ŏ׏鏀����.��R�V�PE_DETAI/h�|zPGL_CON?FIG 8�	����/cell�/$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c�u� ����(���ϯ��� ���;�M�_�q����� $�6�˿ݿ���%� ��I�[�m�ϑϣ�2� ���������!߰��πW�i�{ߍߟ߱�%} F�������/�A�C�i�H�Eߞ���� ������?��.�@�R� d�v������������ ����*<N`r ������ �&8J\n�� !�����/� 4/F/X/j/|/�//�/ �/�/�/�/??�/B? T?f?x?�?�?+?�?�? �?�?OO�?>OPObO�tO�O�O�O����User Vie�w ��}}1234567890�O �O�O_#_5_=T�P��]_���I2�I:O�_ �_�_�_�_�_X_j_�B3�_GoYoko}o�o�o o�op^46o�o@1CU�ovp^5�o �����	�h*�p^6�c�u����������ޏp^7R��)��;�M�_�q�Џ��p^8 �˟ݟ���%����F�L� l?Camera�J���������ӯ���E ~��!�3��OM�_�q�0�������y  e��Y z���	��-�?�Q��� uχϙ�俽���������>��e�5i��c� u߇ߙ߽߫�d����� �P�)�;�M�_�q�� *�<��i�������� �)���M�_�q���� ������������<�û ��=Oas��>� ���*'9 K]f�Q���� ���/�%/7/I/ �m//�/�/�/�/n <��^/?%?7?I?[? m?/�?�?�? ?�?�? �?O!O3O�/<׹��? O�O�O�O�O�O�?�O _!_lOE_W_i_{_�_�_FOXG9+_�_�_o o(o:o�OKopo�o)_ �o�o�o�o�o ��	g�0�oM_q� ��No����o� %�7�I�[�m�&l� n��Ə؏���� � �D�V�h��������� ԟ柍�g�ڻ}�2� D�V�h�z���3���¯ ԯ���
��.�@�R� ��3uF�鯞���¿Կ ������.�@ϋ�d� vψϚϬϾ�e�w��� U�
��.�@�R�d�� �ߚ߬���������� �*���w���v�� ������w����� c�<�N�`�r�����=� w��-�����* <��`r�����������  ��1CUgy��������   -/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_pE_W_i_�  
���(  �%( 	 y_�_�_�_�_ �_�_o	o+o-o?ouo�co�o�o�o�Z* �Q&�J \n������o� ��9�(�:�L�^� p���������܏�  ��$�6�}�Z�l�~� ŏ����Ɵ؟���C� U�2�D�V���z����� ��¯ԯ���
��c� @�R�d�v�����᯾� п�)���*�<�N� `ϧ����ϨϺ���� ����&�8��\�n� ���Ϥ߶��������� E�"�4�F��j�|�� ����������� e�B�T�f�x������� ������+�,> Pb�������� ��(o�^ p�������  /G$/6/H/�l/~/ �/�/�/�//�/�/? U/2?D?V?h?z?�?�/�`@ �2�?�?�?�3�7�P��!f�rh:\tpgl�\robots\�m20ia\cr�35ia.xml �?;OMO_OqO�O�O�Op�O�O�O�O ���O _(_:_L_^_p_�_�_ �_�_�_�_�O�_o$o 6oHoZolo~o�o�o�o �o�o�_�o 2D Vhz����� �o�
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟�ݟ�� &�8�J�\�n������� ��ȯߟٯ���"�4� F�X�j�|�������Ŀt־�8.1 �?�@88�?� ֻ�ֿ�3�5�G�i� ��}ϟ��ϳ������� �5��A�k�U�wߡ�����$TPGL_�OUTPUT �;�!�! ��������,�>� P�b�t������� ������(�:�L�^��p������������2�345678901�������� �"��BTfx�� 4�����
}$L^p��, >��� //$/� 2/Z/l/~/�/�/:/�/ �/�/�/? ?�/�/V? h?z?�?�?�?H?�?�? �?
OO.O�?<OdOvO �O�O�ODOVO�O�O_ _*_<_�OJ_r_�_�_ �_�_R_�_�_oo&o 8o�_�_no�o�o�o�o �o`o�o�o"4F �oT|����\��}�����0�B��T�e�@�������? ( 	 ��Џ ������<�*�L� N�`���������ޟ̟ ���8�&�\�J��� n���������ȯ���"�������*�X�j� F�����|�¿Կ��C� ��ϱ�3�E�#�i�{� 忇ϱ�S��������� �/ߙ�S�e�߉ߛ� y߿���;������� =�O�-�s���ߩ�� ]��������'���� ]�o������������ E�����5G%W }������g�� �1�Ug	w �{��=O	// �?/Q///u/�/��/ �/_/�/�/�/�/)?;? �/_?q??�?�?�?�? �?G?�?O�?OIO[O 9OO�O�?�O�OiO�O �O�O!_3_�O_i_{_�_�_�_�_�_�_�R��$TPOFF_L�IM >�op:���mqbN_S]V`  l�j�P_MON <�6�dopop2�l�aSTRTCHOK =6�f�� bVTCOMPA�T-h�afVWVA/R >Mm�h1d� �o �oop�`ba_DEFP�ROG %|j%�ZERO ZU�ZAUN	�j_D?ISPLAY`|n�"rINST_MSwK  t| ^z?INUSER�odt�LCK�|}{QUI�CKMEJp�"rS7CRE�p6��b?tpscdt�q���b*�_.�ST��jiRACE_C_FG ?Mi�du`	�d
?�u��HNL 2@|i����k r͏ߏ���'�9�K�]�w�I�TEM 2A��� �%$1234?567890����  =<��П�꓏  !���p ��=��c��^����� �����.���R��v� "�H�ί��Я���� ��*�ֿ���r�2ϖ� ����4�޿�ϰ���&� ��J�\�n���@ߤ�d� v��ς������4��� X��*��@���� �ߨ�������T��� x������l����� ���,�>�P������� FX��d����� �:�p"�� o�����F6 HZt~��N/t/ �/��// /2/�/V/ ?(?:?�/F?�/�/�/ j?�??�?�?R?�?v? �?QO�?lO�?�O�OO �O*O|O_`O _�O0_ V_h_�Ot_�O__�_ 8_�_
oo�_@o�_�_ �_Lodo�_�o�o4o�o Xojo3�oN�or�@�o��s�S��B���z�  �h��z ��C�:y
� P�v�]�����UD1:\������qR_GRP 1�C��� 	 @Cp���$��H�6�l�Z��|������f���˟���ڕ?�  
���<�*�`� N���r�������ޯ̯ ��&��J�8�Z����	�u�����sSC�B 2D�  �����(�:�L�^��pς��|V_CON?FIG E����@����ϖ�OUTP�UT F�������6�H�Z�l� ~ߐߢߴ��������� ���#�6�H�Z�l�~� ������������� �2�D�V�h�z����� ����������
�. @Rdv���� ���)<N `r������ �//%8/J/\/n/ �/�/�/�/�/�/�/�/ ?!/4?F?X?j?|?�? �?�?�?�?�?�?OO /?BOTOfOxO�O�O�O �O�O�O�O__+O>_ P_b_t_�_�_�_�_�_ �_�_oo'_:oLo^o po�o�o�o�o�o�o�o  $����!�bt �������� �(�:�-o^�p����� ����ʏ܏� ��$� 6�G�Z�l�~������� Ɵ؟���� �2�D� U�h�z�������¯ԯ ���
��.�@�Q�d� v���������п��� ��*�<�M�`�rτ� �ϨϺ��������� &�8�J�[�n߀ߒߤ� �����������"�4� F�W�j�|������ ��������0�B�S� f�x������������� ��,>Pa�t ��������(:L/x���k}gV�K ���//&/8/J/ \/n/�/�/�/W�/�/ �/�/?"?4?F?X?j? |?�?�?�?�/�?�?�? OO0OBOTOfOxO�O �O�O�?�O�O�O__ ,_>_P_b_t_�_�_�_ �O�_�_�_oo(o:o Lo^opo�o�o�o�o�_ �o�o $6HZ l~����o�� �� �2�D�V�h�z� �������ԏ���
� �.�@�R�d�v����� ����Ϗ�����*� <�N�`�r��������� ˟ޯ���&�8�J��\�n���������Ż��$TX_SCRE�EN 1G�g�}i�pnl/��gen.htmſ�*�<��N�`ϽPan�el setupd�}�dϥϷ����������ω�6�H�Z� l�~ߐ�ߴ�+����� ��� �2�߻�h�z� ������9�g�]�
� �.�@�R�d������ ����������}��� <N`r��; 1��&8� \��������QȾUALRM_�MSG ?��� �Ȫ-/?/p/ c/�/�/�/�/�/�/�/�??6?)?Z?%SEoV  -�6�"ECFG Iv��  ȥ�@�  A�1  w B�Ȥ
 [? ϣ��?OO%O7OIO�[OmOO�O�O�G�1G�RP 2J�; 0Ȧ	 �?�O �I_BBL_NO�TE K�:T?��lϢ��ѡ�0RDEFP�RO %+ (%N?u_Ѡc_�_�_�_ �_�_�_o�_o>o)o�boMo�o\INUSER  R]�O�o�I_MENHIS�T 1L�9  �(�0 ��)�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,1133,�1�oDVhz~��9 }9361� ����r�$�6�H� Z�l�~������Ə؏ ����� �2�D�V�h� z�	�����ԟ��� 
���.�@�R�d�v��� �����Я����� 9Rq��B�T�f�x��� ������ҿ����� ��>�P�b�tφϘ�'� 9���������(߷� L�^�p߂ߔߦ�5��� ���� ��$����Z� l�~����C����� ��� �2��/�h�z� ��������������
 .@��dv�� ���_�* <N�r���� �[�//&/8/J/ \/��/�/�/�/�/�/ i/�/?"?4?F?X?C� U��?�?�?�?�?�?�/ OO0OBOTOfO�?�O �O�O�O�O�O�O�O_ ,_>_P_b_t__�_�_ �_�_�_�_�_o(o:o Lo^opo�oo�o�o�o �o�o �o$6HZ l~i?{?���� ��2�D�V�h�z� ���-�ԏ���
� ���@�R�d�v����� )���П������� ��N�`�r�������7� ̯ޯ���&���J��\�n�����������$UI_PANE�DATA 1N����ڱ?  	�}����`�!�3�E�W� )Y� }�7�뿨Ϻ������� �i�&��J�\�C߀� gߤߋ������������"�4��X�7�� �q}�ϕ����� ����B����%�I�[� m������
������� ����!E,i{ b������l�ܳ7�<N`r ����-���/ /&/8/�\/n/U/�/ y/�/�/�/�/�/?�/ 4?F?-?j?Q?�?�? %�?�?�?OO0O�? TO�xO�O�O�O�O�O �OKO_�O,__P_b_ I_�_m_�_�_�_�_�_ oo�_:o�?�?po�o �o�o�o�oo�o sO $6HZl~�o� ������ �2� �V�=�z���s����� ԏGoYo�.�@�R� d�v�ɏ����П� �����<�N�5�r� Y�������̯���ׯ �&��J�1�n���� ���ȿڿ����c� 4ϧ�X�j�|ώϠϲ� ��+��������0�B� )�f�Mߊߜ߃��ߧ� ��������P�b� t����������S� ��(�:�L�^���� i�����������  ��6ZlS�w�'�9�}���"4FX)�}�� l�����/j '//K/2/D/�/h/�/ �/�/�/�/�/�/#?5?�?Y?��C�=��$U�I_POSTYP�E  C�?� 	 e?�?��2QUICKME/N  �;�?�?��0RESTORE� 1OC�?  �L?��!6OCC1O��maO�O �O�O�O�OuO�O__ ,_>_�Ob_t_�_�_�_ UO�_�_�_M_o(o:o Lo^oo�o�o�o�o�o �oo $6H�_ Ugy�o���� �� �2�D�V�h�� ������ԏ��� �w�)�R�d�v����� =���П������*� <�N�`�r������� �ޯ���&�ɯJ� \�n�������G�ȿڿ������7SCRE��0?�=uw1sc+@u2K�U3K�4K�5K�6K��7K�8K��2USE1R-�2�D�ksMì�U3��4��5��6���7��8���0NDO_CFG P�;�� ��0PDATE� ���N�one�2��_IN_FO 1QC�@��10%�[���Iߊ� m߮��ߣ�������� ��>�P�3�t��i����<-�OFFSET T�=�ﲳ$@ ������1�^�U�g� ��������������� $-ZQcu����?�
����UFRAME  �����*�RTOL_�ABRT	(�!E�NB*GRP �1UI�1Cz  A��~��~���������0UJ�9MSKG  M@�;N�%8�%��/�2V7CCM��V�ͣ#+RG�#Y�9���/j����D�BH�Yp71C���37f11?�C0�$MRf�2_�*S�Ҵ�	����~XC5G6 *�?�6����1$�5���A@v3C��. ��8�?��OOKOx1�FOsO�5�51���_O�O�� B����A2�DWO�O7O _�O8_#_\_G_�_k_ }_�__�_�_�_�_"op�OFoXo�%TCC�#A`mI1�i������� GFS��2a�Z; �| 2345678901�o �b�����o��!5�a�4BwB�`56 �311:�o=L �Br5v1�1~1�2��}/ ��o�a��#�G Yk}�p����� ��ُ�1�C�U�6� H���5�~���ߏ����	���4�dSELE�C)M!v1b3�VIRTSYNC��� ���%�SIO�NTMOU�������F��#bU���U�(u� FR:\H�\��A\�� ��� MC��LOG���   UD1懦EX����' B@ �����̡m��̡  OB�CL�1�H� ��  =	 1�- n6  -#������[�,S�A��`=��͗���ˢ��TRAIN�⯞b�a1l�
0d�$j�T2cZ; ( aE2ϖ�i��;�)� _�M�g�qσϕϧ���������	��F�ST�AT dm~2@�zߌ�*j$i߾���_GE�#eZ;�M`0�
� 02���HOMIN� fU��U� ~�(����БC�g�X����JMPERR 2=gZ;
  ��*j l�V�7���������� ����
��2�@�q�d��v�B�_ߠRE� h\Wޠ$LEX��iZ;��a1-e��VMPHASE  5�r�c&��!OFF/��F�P2n�j�0R�㜳E1@���0ϒE1!1?s33�����ak/�kxPk䜣!W�m[�䦲 �[����o3;� [i{ ����/� O�?/M/_/q/��/ ��//�/'/9/�/=? 7?I?s?�/�?�/�/�? �??Om?O%O3OEO �?�?�O�?�O�O�?�O �O�O__gO\_�OE_ �O�_�O�O/_�_�_�_ oQ_Fou_�_|o�o�_ �oo�o�o�o�o;oMo ?qof-�oI�� ���7�[P� ��������ˏ� �!�3�(�:�i�[�ŏ�g�}������TD__FILTEW�n��g �ֲ:���@� ��+�=�O�a�s��� ������֯������0�B�T�f�x���S�HIFTMENU� 1o[�<��% ��ֿ����ڿ���� I� �2��V�hώ��π�ϰ�������3�
��	LIVE/SN�AP'�vsflsiv��E����/ION * Ub�h�menu~߃���߰�ߣ���p���a	����E�.�50�s�P�@� ��AVɠB8z�z��}���x�~�P�� ����MEb�Կ�<�0���MO���q���z�WA�ITDINENDb������OK1N�OUT���SD���TIM����o�G���#���C����b������RELE�ASE������TM��������_AC�T[�����_DA�TA r��%�L����xRDIS�b�E�$XVR��s���$ZAB�C_GRP 1t��Q�,#�0�2\���ZIP�u'��&����[MPCF_G 1v�BQ�0�/� w�<�ɤ� 	�Z/  85�/�/H/�/l$?��+�/�/ �/?�/�/???r?�?  �D0�?�?��?�?�?�;���x��]hYLIND�֑y� ���? ,(  *VOgM�.�SO�OwO�O�M  i?�O�O^PO1_�OU_ <_N_�_�O�_�_�__ �_�_x_-ooQo8o�_0�o�oY&#2z� ���oC�e?@a?>N|�oq����q�A�$DSPHER/E 2{6M��_� ;o���!�io|W� i��_��,��Ï��� Ώ@��/�v���e�؏ ��p����������6ZZ�� �N