��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER� q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*�6��4OS ��DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� 0�BRE-  ? � �0�BB{F S{T� M�D|TRS$STD6XlQCWFA� 7X�QCW��"YV�"eS/ �A7 �  $�@TI�Nd@�0SULگ �R_@ g $}@ SW�@�RO�RR%	� �P�T� �@J�U� �SqFS4DN6
 �2P�0_@�cFOL[d!$�FIL� jjE�P��C�S�aDIG4R_C_SCA��c�INTTHRS�_BIdA�dSMA9L�bCOL�b9G�`� �� ��_IVTIM��$!0B"$S�?0xCCBDDN���-qI2wT2wDE�BUdA\!SCHN�"TOfa0�! �  Q0mr<0V� �;!�r~AUTTUN�� TRQa�uE�40N �qFS3A	XG  � 1eb}tj�rI�v
	"G_gr>7 l �!�3>@WEIGH�q�2� uS_5QF(�T�2�WA� 	pEsNTERVA�; -  Q�� S!�t�AS0S��$J-_STAF�p JQg���1(�U��2��3��W����� hqx��"COG+_X�Y�Z�ҁCM�p?�p�܂RSLT�4��D��D��	"_�p_�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDB	"I%�0 ,$M"Pp30f��� d��:pG p"��HCDv�GV�#GVY��Z�JDO5�,q���S��$R��E_�8@{٣�pAP�HBC��$VF6�P��2L��蘨@IL[����;����;�d@���RG���NGEW_���r�Q}�8��ڡ�5OBOA@fQY�sW2/�G<�	����ȴ\�2�E�KP��NUCNPRGOVp����@`d_TW�cj,�G�E^!NV2#�C�c0@�WTS�T�RL_SKI2!�$SJ�Q��NQpG�W��	"��7 �\ ;0FR]b� � CMDC���T0�b���TO?�� � �5گ���_�Ah �0 '��ALARM��_�*�TOT6�F#RZn l�,!Y 3�� X!��mӥ�X �Œ`X P�ʕ�U#��2��2
�8X#Z���FIX�8�ґF�"��IT�`IeB�PN_d��CH��%��_DFL _�B#F2N�ڶ�3����� ��3�"�����ʷ�� ����3��3p
��X��DIA����/#� ���%�����[1��g1�[� ��Z��#��!���%���$0�@
p��7F���D�� HA�pU��5����v�FSIW.6 �2PN@�`uR>!�PHMP�`HCK%���>0G�'�*#e A����pN�T��^H	��HUFARzs3��A��Ugv�Ca�$v0Q ����@p�@� � � SI0��P��5�IRT�U_��� %SV �2���   ��6>0]@]	xQ�EF@ ��oP�  @pP�� �//'/P9/K/U%@pd@p
m hK�/w/�/�/�(� �$��/� �/�/?.8 e"�/?J?\?r?8?�? |?�?�?�?�?�?�?>O 4ObOO�OTO�O�OjO |O�O�O�O_�O(__ \_f_�_B_�_�_�_�_  o�_$o�_Ho>oo^b �/�ot��%�/�o�o�k�	MC: 5�678  Af�sdt1 78901234q#^5w  	q 6x�z.Ops�'��j l�o�o���������,��5�DMM �)5�A ��x��������=���OR �2	Q� ���m��_� tuBo?)DN��S4D 
Q�!tY�d�!Ls|�q�`rƈ̀?�l�B�򴐠�$ ONFIoG �(�P� �� �������i!��� 2��,
Hand �guide��?��3���  �aX��с��ь�g#�=���A�� ύ�������p�ݯ �(��L�7�p�[����m*������ ʿܿ� ��$�6�H� Z�lɌ��ό��ϰ���@�����
�C�E�IW 2Q�(�0�C -�zՀ�Fտ��_`πB����d��C�  ��uq=#{�
_aNnk(���K����̥@�{�e��=D�����_a;����8I��_aIt$ ��$F�>����k"���Q�F��3]儢ѯǯ���x!�/�``+������.�����_a$�{����(4$��弥��>�E��B�<~w%�_a8E�=y5�;�jA������Q�>��]�_a?��m��箑��x��~u1�?�33��<��0�:�o�����0�����LSB ��~uq�ӻ��m��S]���8��� ���t�	eF|���]��߯����n���;�.����3�'	�����B���4* 2�/V��%D�DH  *%v�+��^-���
�/��/u/~u�J/l/�)AI��/�/8�?/ A��n5��p��4vO?;)�7 �?�?�o�?�8Jhq�?��?zyjG�_FSIW Q��9��O �O�Ou�