��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81s!�J3> �! � $SOFT��T_IDk2TOT�AL_EQs $̅0�0NO�2U SP?I_INDE]�5�Xk2SCREENu_(4_2SIGE0�_?q;�0PK_�FI� 	$T�HKYGPANE��4 � DUMM�Y1dDDd!OE4�LA!R�!R�	 � $TIT�!$I��N �Dd��Dd �Dc@�D5�F6��F7�F8�F9�G0 �G�GJA�E�GbA�E�G�1�G1�G �F�G2��B!SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C?CFS_UT~p0 "�1�3�#�ؗ`qX"�}R0  4F OIMCM�`O#S�` ��upi �_�p�EBA�!���M/� h�pIMPEE_F�N��N��0�@O��r�D_�~��n�Dy�F� dCCq_�r0  T� '��'�DI�n0"���p�P�$�I������F�t X� GRP0��=M=qNFLI�7��0UIRE��$g"~� SWITCH5��AX_N�PSs"C�F_LIM�� � �0EED���!��qP�t�`PJz_dVЦMODEh��.Z`�PӺ�ELBOF� ������p@� ���3���� FB�/��0�>�G�� �� WARNM��`/��qP��n�N�ST� COR-�0bFLTRh�TR�AT�PT1�� $ACC1a��N ��r$ORI�o"V��RT�P_S� C�HG�0I��rT(2��1�I��T�I1���� x pi#�Q��HDRBQJ; CQ�2L�3L�U4L�5L�6L�7L�T N�9s!��O`S <F +�=�O�x�#92��LLECy�}"MULTI�b@�"N��1�!���0T��w �STY�"�R`�=l�)2`��8��*�`T  |� �&$��۱m��P�̱��UTO���E��EXT����ÁB���"G2� (䈴![0������<�b+�� "D"���ŽQ��H<煰kcl�9�#���1��ÂM�ԽP���" '�3�$ �L� E���P<��`A�$JOBn�T����l�TRIG3�% dK�������<���\h��+�Y���_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`�0Z���0��P_�P��n@ ( @F RO.���&�t�IT�c�N�OM�
����S*��P`T)w@���bZ�P�d���RA�0଱2b"����
$T\����MD3�T�䢣`U31���p(5!H,Gb�T1�*E�7�c�KAb�WAb�cA4#�YNT���PDB�GD�� *(��P�Ut@X��W���AqX��a��eTAI^c�BUF��0!+� � 7n�PIVW�*5 P�7M�8�M�9
0�6F�7SI�MQS@>KEE�3PATn�^�a" 2�`#�"�L64FIX!, ���!d��bD�2Bus=CCI��:FPCH�P:BAD �aHCEhAOGhA]HW�_�0>�0_h@�f�A k���F�q\'M`#�"t�DE3�- l�p�3G��@FSOES]F gHBSU�IBS9WC���. ` ��MA�RG쀳��FAC<Lp�SLEWx`Qe�ӿ��MC��/�\pSM_JBM����QYC	g�ex��Д0 ā��CHN-�MP�#$G� Jg�_� #���1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�f�JR���rSEGF�R�PIO� ST�RT��N��cPV5���!41�r��
r�>İ�b�B�O�2` +�[���,q E`&�,q`y�Ԣ}t���yaSIZ%���t��vT�s� �z�y,qRSINF}Oбc��@�k��`��`�`L��8� T`7�CRCf�ԣCC/�9��`a�uah�ub'�MIN��uaD�s�#�G�D�YC��C �����e�q0��� �SEV�q�F�_�eF��N3�s�ah��X�a+p,5!�#1��!VSCA?� A䕖s1�"!3 � �`F/k��_�U��g��]���C�� a�s��R>�4� �����N����5a�R�HA;NC��$LG��P�6f1$+@NDP�t�AR5@N^��a�q���c��ME�18���}0f��RAө�AZ �𨵰�%O��FCT K��s`"�S�PFADIJ�OJ�ʠ� ʠ���<���Ր��qGI�p�BMP�dp�p�Dba��AES�@�	�K�W_��BAS��� �G�5  zM�I�T�CSX[@�@�!62�	$X����T9�{sC��N��`�a~P_HEIG9Hs1;�WID�0�aVT ACϰ�1�A�Pl�<���EXP�g���|��CU�0M�MENU��7�T[IT,AE�%)��a2��a��8 P�� a�ED�E  ��PDT��REM�.��AUTH_K�EY  ������ ��b�O	�!}1ERsRLH� �9 \� ��q-�OR�DB�_I�D�@l �PUN_O|��Y�$SYS0Ш�4g�-�I�E�E�V�#�`at(�PX�WO�� �: $�SK7!f2%�Td�T�RL��; �'AqC�`��ĠIND9�DJ.D��_��f1X��f���PL�A�R#WAj���SD�A���!+r|��UMM3Y9d�F�10d�&�d��J�<��}1PR�w 
3�POS���J�= �$�V$�q�PL~�>����SܠK�?����CrJ�@����ENE�@�T��A���S_�R�ECOR��BH� 5 O�@=$LA�>$~�r2�R�0�`�q�b`�_Du��0RO�@�aT[�Q��b�������! }У�P�AUS���dETU�RN��MRU��  CRp�EWM<�b�AGNAL:s2�$LA�!?{$PX�@$P�Fy A �Ax�C0 #ܠDO�`X�k�W��v�q�GO_AWA�Y��MO�ae����]�CSS_CCS;CB C �'N��CERI��гJ`u�QA0�}��@.�GAG� R�0�`���{`��{`OF��q�5��#MA���X��0&шL�L�D� �$ ���sU�D)E%!`��>�OVR10W�,��OR|�'�$ES�C_$`�eDSBIOQ��l ��B�VIB&� �c,��p���f�=pSSW�l��f!VL��PL��>�ARMLO
��`a����d7%SC ��bALspH�MP Ch �Ch �#h �#h 5�UU���C�'�C@�'�#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$�4�C�P3Wұ46�$VOLT37$$`�*�^1��$`�O1*�$o��0RQ�Y��2b4�0DH_THE����0SЯ4�7ALPH�4�`��D�7�@ �0�qb7�rR�5�88� ×����"��Fn�M�ӁVHBPFUAFL�Q"D�s�`�THR��i2dB�����G(��PVP���������
��1�J2�B�E�C�E�CPSu�Y@��Fb3 ���H�(V�H:U�G�@
X0��FkQw�[�Na��'B���C INHBcFILT���$ ��W�2�T1�[ ���$���H YАAF�sDO��Y�Rp�  fg�Q�+�c5h�Q0�iSh�QPL���W<qi�QTMOU�#c �i�Q\��X�gmb��vi��h�bAi�fI�aH!IG��ca	xO��ܰ4��W�"vAN-u!���	#AV�H!P�a8$P�ד#p�R_�:�A�a��B�N80�X�MCN���f1[1�qVE�p��Z2;&f�I�QO�u�rxZ�wGldDN{G|d���aF>!�9��aM�:�U�FWA�:�M l���X�Lu��$!����!l�ZO����0%O�blF�s�13�DI�W�@��Q���_�|�!CURVA԰&0rCR41ͰZ�C<� r�H�v���<�`��<�(�f�CH�QR3�S����t���Xp�VS_��`�ד�F��ژ����?NST�CY_ E L����1�t�1��U��U24�2B�NI O7�x�����DEVI|� F��$5�R�BTxSPIB�P����BYX����T���HNDG��G H tn���L��Q�C���5��Lo0 H���f��FBP�{tFE{�5�t��T��I�DyO���uPMCS�v�>�f>�t�"HOT�SW�`s�
?ELE��J T���e�2���25�� O� ��HAA7�E��344�0?ܘ�A�K �� MD�L� 2J~PE ��	A��s��tːÈ�s�JÆG!��rD"��0������\�TO��W��	��/��SLAV��L  �0IN�Pڐ���`%ن_C�Fd�M� $n��ENU��OG��`b�ϑ]զP�0`�<��]�IDMA�Sa��\�WR�#��"]�sVE�$a�SKI�S!Ts��sk$��2u���J�������	��Q����_SVh�EXC�LUMqJ2M!ONLD��D�Y��|�PE �ղI_V�APPsLYZP��HID-@�Y�r�_M�2��VRFY�0��r�1�c�IOC_f�� 1�������O��u�LS����R$DUMMKY3�!���S� L_TP/Bv�"����AӞ�ّ N ����RT_u��� Ґ�G&r[�O{ D��P_BA�`g�3x�!F R��_5���H���?���� �� P $<�KwARGI��� ~q�2O ��wSGNZ�Q �~P/�/PIGNs�l��$�^ sQANNUN�@�T<�U/�ߴ�LAzp]	Z��d~��EFwPI��@ R @�F�?IT�	$TOTA%��d���!��M�NIY�!S+���E�A[�
oDAYS\�ADx��@��	� �EF_F_AXI?�TI�̈0zCOJA ��ADJ_RTRQ
��Up��<P�1D ��r5̀Ll�T �0? ]P�"p��mtpd��V 0w�G�h�������SK�S�U� ��CTRLw_CA�� W��TRANS�6PI?DLE_PW���!h��A�V��V_��l�V �DIA�GS���X� /�$2�_SE�#TAC���t!�!0z*@&��RR��vPA���p ; SW�!�!� � ��ol�U��oO�H��PP� ��I9R�r��BRK'#��"A_Ak���x 2x�9ϐZs2��%l�W��0t*�x%RQDWf�%MSx�t5AX�'��"��LIFECAYL���10��N�1 {"�5Z�3{"dp5�Z�U`}�MOTN°Y�$@FLA�cZO3VC@p�5HE	��SUPPOQ�ݑAq�� Lj (C�1_XT6�IEYRJZRJWRJ��0TH�!UC��6�XZg_AR�p��Y2�H�COQ��Sf6AN��w$���ICT�E�Y `��CACHE�C9�M��PLAN��UFFIQ@�Ф0<�1�	��6
��MSW��EZ 8�KEY�IM�p��TM~�S@wQq�wQ#�����OCVIE� �[; A�BGL��/�}�?� 	�?��D�\p�ذST��!�R� �T� �T� �T<	��PEMAIf�ҁ���_FAUL��]�Rц�1�U��� �TRE�?^< $Rc�u�S�% IT��BU!FW}�W��N_� 'SUB~d��C|��8Sb�q�bSAV�e�b�u �B��� �gX�^P �d�u+p�$�_~`�e�p%yOTT����s�P��M��OtT�LwAX � ��X~`9#�c�_G�3
�YN_1�_�D��1 �U2M���T��F��H@ g�`� 0p��Gb-s7C_R�AIK���r�t�RoQ�u7h�q'DSPq��rP��A�IM�c6�\����s2��U�@�A�sM*`I�P���s�!DҐ6�T!H�@n�)�OT�!6��HSDI3�ABSC���@ Vy���� �_D�CONVI�G���@3�~`	F�!�pd��psq�SCZ"���sMER�k��qFB��k��pEiT���aeRFU:@�DUr`����x�CAD,���@p;cHR�	A!��bp�ՔՔV+PSԕC���	C��pN�ғSp�_cH *�LX� :cd�Rqa�| ����W� �U��U��U�	�U�TOQU�7R�8R�9R���0T�^�1k�1x�1���1��1��1��1*��1ƪ2Ԫ2^�k�U2x�2��2��2��U2��2��2ƪ3Ԫ%3^�3k�x�3���To���3��3��3ƪ54Ԣ%�XTk!0�d <� 7h�p�6�p�O��p����NaFDR^Z$eT^`V��Gr����䂴2REMr� Fj��BOVM�z�A�TROVٳDT�`-�MX<�I�N��0,�W!IND�KЗ
w�׀�p$DG~q36��P�5�!9D�6�RIV���2��BGEAR�IO�%K�¾DN�p��J��82�PB@�CZ_MCCM�@�1��@U���1�f ,②a?� ���PI�!�?I�E��Q�U��H�am���g� _0Pfq�g RI9e���bE�TUP2_ h � �cTD�p����! a�����BAC�ri T�P�b�`Z�) OG��%�8��p��IFI�!�p0m�>��	�PT�"���FMR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4��@C��Uk���� T�FS#p�Tl� P���e�qP�p�$EX_���1PM2��2� 3�5�s�G ���m ���֍�SW�eOe6DE�BUG���%GRt���pU�#BKU_��O1'� �@P�O�I5�5M�S��OOfswSM���E�b�Q�0�0_E n �0��P_�TERM�o��`�ORI+�p<��P�SM_���br�q��0�TA��r���UP>�Rs� -�1�2�n$�' o$S�EG,*> ELTO���$USE�pNFIAU"4�e1��|�#$p$UFR����0ؐO!�0����OT��'�TAƀU�#N;ST�PAT��P��"PTHJ����Ep�P rF�V"ART�`�`%B`�abU!REL<:�aSHFT��V!\�!�(_SH+@M$�D��� ��@N8r�����OVRq��rSH�I%0��UN� �aAGYLO����qIl�����!�@��@ERV ]��1�?:�¦'�2`��%��5�%�RCq��EASYM�q�EV!#WJi'��}�E���!I�2��U@D��q�%Ba��
5Po��0�p6�OR�MY� `GR��t2b5n� � p��UPa�Uu Ԭ"�)���TOCO!S�1POP ��`�p(C�������Oѥ`KREPR3��aO�P,�b�"ePR�%WU�.X1��e$PWRf��IMIU�2R_	S��$VIS��#(AUqD���Dv" v���$H���P_AD+DR��H�G�"�Q��Q�QБR~pDp1�w H� SZ�a��e`�ex�e��SE�l�r��HS��MNv?x ���%Ŕ��OL���p<Px��-��ACROlP<_!QND_C��גx�1�T �ROUPT���B_�VpQ�A1 Q�v��c_��i���iр�hx��i���i��v�AMCk�IOU��D�g�fsu^d�y $|�P_D��VB`b�PRM_�b?�H�TTP_אHaz{ (��OBJEr�l�P��$��LE�#��s`{ � \��u�AB_x�T~��S�@�DBGL�V��KRL�YHIoTCOU�BGY �LO a�TEM���e�>�+P'�,PSS�|�P�JQUERY�_FLA�b�HW(��\!a|`u@�3PU�b�PIO��"��]�ӂ/dԁ=dԁ�� _�IOLN��}�����CXa$SL�Z�$INPUTM_g�$IP#�P��L'���SLvpa~���!�\�W�C-�B?�I�O�pF_ASv��$L ��w �F1"G�U�B0m!���0HY��ڑ����UOPs� ` ������[�ʔ[�і"�[PP�SIP�<�іI��2��0�IP_MEsMB��i`� X��cIP�P�b{�_N�`����R�����bSP��p$FO�CUSBG�a~�U=J�Ƃ �  � �o7JOG�'�DI�S[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A���APHIb�Qt�]�D� J7J\����� _KEYt�� �KՀLMO�Na���$XR���ɀ��WATCHa_��3���EL��b}Sy~���s� f �!V�g� �CTR�3򲓥��LG�D�� �R��I�
LG_SIZ���J�q XIƖ�I�FDT�IH� _�jV�GȴI�F�%S O���q �Ɩ���v������K�S����w�kR�N����E�@�\���'�*�U�s�5��@L>�4�DAUZ�EA�pՀ�Dp�f��GH�B�ᢐBOO>��� C���P�IT���� ��RE=C��SCRN�����D_p�aMARG f�`��:���T�L���S�s��W�Ԣ�I�JGMO�MNC�H�c��FN��R�Knx�PRGv�UF���p0��FWD��HL.��STP��V��+�X��Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28�����Gh�0PO��������M8�Ģ��EX��TUIv�I��(�4�@� t�x�J0J�~�P��J0r��N�a�#ANA���O"�0VAIA��dC�LEAR�6DCS�_HI"�/c�O��O�SI��S��IGN_�vpq��uᛀT�d� DEV�-�LLA �°BUTW`��x0T<$U�EM��Ł�����0�A�R���x0�σ�a�@OS1*�2�3�a�`� �ࠜh�AN%�-���-�IDX�DP��2MRO��Գ!�S�T��Rq�Y{b! _�$E&C+��p.&A&���`� L��ȟ%Pݘ��T\Q�UE�`�Ua��?_ � �@(���`�����# �MBG_PN@ R`r��R�w�TRIN��P���BASS�a	6IR�Q6��MC(��{ ��CLDP��> ETRQLI��!D�O9=4FLʡh2�A�q3zD�q7��LD8q5[4q5ORG�)� �2�8P�R��4/c�48=b-4�t� �rp[4(*�L4q5S�@TO0Qt��0*D2FRCLM�C@D�?�?RIAt,1I�D`�D� d1��R�QQprpDSTB�
`� �F�HA�XD2���G�LEXC#ES?R+2�AMhPa�͠�BD4�ёB�qj`�`�F_A�J��C[�O�H� K���# \���bTf$� ���LI�q�SREQU7IRE�#MO�\�a^�XDEBU��� uL� M䵔 �p`���P�c�AA�� N��
Q�q�/�&���f-cDC��B�IN�a�?�RSM�Gh� N�#B��N�a,1aPS}T9� � 4��7LOC�RI���;EX�fANG��A^,1ODAQ䵗�@c$��9�ZMF�� ���f��"��%u#Ю�VSUP�%aF�X�@IGGo�� �rq�"��1��#B��$���p%#by��rx����vbPDATA�K�pE;���Ρ��M܋�*� t�`MD
�qI��)�v� �t�A��wH�`��tDIA<��sANSW��t(h���uD��)�bԣ�(@$`� PCU�_�V6�ʠ�d�PLODr�$`�R���B��B�p�����+2RR}2�E�  ���V�A/A d$C'ALI�@��G~��2��!V��<$R��SW0^D"��A�BC�hD_J2SqE�Q�@�q_J3M�
G�1SP�,��@	PG�n�3m�u�3p�@���JkC���2'AO�)IMk@{BCSKAP^:ܔ9�wܔJy�{BQܜ�����`�_AZ.B��?�ELx��YAOCMP�c|A)��RT�j���c1�ﰈ��@1���t����Z��SMG��pԕ� ER!����AINҠACk�@p����b�n _��������D�/R�f�DIU��CDH�@t
�#a�q$V�lFc�$x�$�� �`@���b��̂�E��H �$BE�LP����!ACCE�L���kA°IR�C_R�pG0�T<!�$PS�@B2L  ����W3�طx9� ٶPATH���.�γ.�3���p�A_@��_�e�-B�`C�_MG�$D�D��ٰ��$FW��@�p����γ����D}E��PPABN�ROTSPEEu�����O0��DEF�>Q����$USE)_��JPQPC��J�Y����-A 6qYN��@A�L�̐�L�M�OU�NG��|�O9L�y�INCU��a��¢ĻB��ӑ�AENCS���q�B�����D�IN�I�����p�zC�VE�����2�3_U ��b�LOWL���:�O0��0�Di�B�PҠ� ��rPRC����MOS� �gTMOpp�@-GPE�RCH  M�OVӤ �����!3�yD�!e�]�6�<�� ʓA����LIʓdWɗ��p:p3�.�I�TRKӥ�AY����?Q^����m�b��`p�CQ�� MOM�B?R�0u��D����y�0Â��D�UҐZ�S_BCKLSH_C����o� n��TӀ���
c��CLALJ��A8��/PKCHKO0��Su�RTY� �q���M�1�q_
#c�_�UMCP�	C���SsCL���LMTj��_L�0X����E �� �� ���m�`h���6��PC��B��H� �P�ŞCN@�"XT����CN_b��N^C�kCSF����V6����ϡj����nCAT�SH s�����ָ1���֙�0��������PA���_P���_P0� e�`��O1u�$xJG� �P{#�OG���TORQU(�p�a�~�����Ry������"_W ��^�����4t�
5z��
5I;I ;Iz�F��`�!��_8�1��VC"��0�D�B�21�>	P8�?�B�5JRK�<�2��6i�DBL_SMt�Q&BMD`_DLt�&BGRV4
Dt�
Dz��1H_���31�8J�COSEKr�EHLN �0hK�5oDt�jI��jI <1�J�LZ1�5Zc@y���1MYqA�HQBTH|WMYTHET09�NK23z�/Rn�r@[CB4VCBn�CqPASfaYR<4gQt�gQ�4VSBt��R?UGT	S���Cq��a��P#x���Z�C$DUu  ��R䂥э2�Vӑ��9Q�r�f$NE�+p!Is@�|� �$R�#Q�A'UPeYg7EBHBALCPHEE.b�.bS�E �c�E�c�E.b�F�c�j�FR�VrhVghd��lUV�jV�kV�kV�kUV�kV�kV�iHrh@�f�r�m!�x�kH�kUH�kH�kH�kH�i�OclOrhO��nO��jO�kO�kO�kO*�kO�kO�FF.bTQ𰉔E��egSPBA�LANCE��RLmE�PH_'USP���F��F��FPFULC�3��3��E��{1�l�UTO_p ��%T1T2t���2NW�����ǡ��5�P`�擳�T�OU�|��� INSEG���R�REV��R���D3IFH��1���F�1�;�OB��;C���2� �b�4LC�HWAR��;�AB�W!��$MECH`]Q�@k�q��AXk��P��IgU�i�� �
���!����ROBF��CR��ͥ*��C��_s"T �� x $WEI3GHh�9�$cc�2� Ih�.�IF ќ�'LAGK�8SK��nK�BIL?�OD��LU��STŰ�P�@; �����������
�Ы�L��  2y�`�"�DEBU.��L&�n��PMMY�9��NA#δ9�3$D&���$��� �Q �DO_:�A��� <	����~��L�BX�P�ND��+�_7�L�t�OH  �� %��T���ѼT������TICK/�C�T1"��%������N��c�Ã�R L�S���S�|����PROMPh��E� $IR�� X�~ ���!�MA�I�0��j���_9�����t�l�R�0C�OD��FU`�+�I�D_" =�����G�_SUFF<0 �3�O����DO ��ِ��R��Ǔن�S�����!{������	�Hn)�_FI��9��7ORDX� ����C36��X������GR9�S��ZDT�D��v�ŧ4{ *�L_NA4����K��DEF_I [�K���g��_���i�`�Ɠ�š���IS`@i �萚����e�D���4�0i�Dg�(���D� O��LOCKEA!uӛ�`�Ͽ���{�u�UMz� K�{ԓ�{ԡ�{���� }��v�Ա��g��� ���^���K�Փ� ����!w�N�P'���^���,`�W\�[R�	7�TEFĨ� �OULOM�B_u�0�VI]SPITY�A�!}OY�A_FRId���(�SI���R�������3���WB�W��0��0_,�EAS%��!�P& "���4p�G;�_� h ��7ƵCOEFF_Om����m�/�G!%�S.�߲CA5����u��GR` � �G $R� �X]�TME�$R�s�Z�/,)�ER�T;�:䗰7�  ]�LL��S�_SV�(�$~����@����{ "SETU��MEA��Z�x0�u�|����� � � 6�� ȰID�"���!*��&P���*�F�	'����)3���#���"�5;`*�N�REC���!7��SK_��� �P	�1_USER���,��4���D�0��VEL,2�0���2�5S��I��0�MTN�C�FG}1�  ���Oy�NORE���3��2�0SI��1�� ��\�UX-��ܑPDE�A _$KEY_�����$JOG<EנS�VIA�WC�� 1DS�Wy���
��CMULT�GI�@@C��2?� 4 �#t�+�z�XYZ��쑡����z� �@_ERR���� ��S L�-����@��s0BB$B�UF-@X17ࡐM�OR�� H	�CU�A3�z�1Q�
��3<���$��FVI��2SbG��� � $SI�@ G�0VO B`נ�OBJE&�!FAD�JU�#EELAYh' ���SD�WOU��p�E1PY���=0Q�T i�0�W�DI�R$ba�pےʠD#YN�HeT�@���R�^�X����OP�WORK}1�,>�SYSBU@p 1�SOP�aR�!�jUĔk�PR��2�ePA`�0�!�cu� 1OP��EUJ��a'�D�Q/IMAG�A	��`fi�IMACrIN,��bsRGOVRD=a�b�0�aP�`sʠ�� �^uz�LP�B��@��!PMC_E(,�Q��N@�M�rǱb��1Ų7�=qSL&��~0���$OVSAL\G*E��*E2y�Ȑ�_=p�w��>p�s@���s	����y��t�#}1� @�@;���MOE�RI#A��
N���X�s�f�����PL�}1�,RTv�m�AT�USRBTRC_T(qR��B �����$� �Ʊ��,�~0� D��`-CSALl`�SA0���]1gqXE���%���C��J�
���cUP(4����PX���؆�q��3�w� ��PG�5� $SUB�������t�JMPWAITXO��s��LOyCFt�!D=�CVF	ь�y�⻑R`�0��CC_�CTR�Q�	�IG�NR_PLt�DB�TBm�P��z�BW�)����0U@���IG��a��Iy�TNLND��Z�R]aK� N��B�0�PE�s���r���f�SPD}1� L�	�A�`gఠ�S��U!N�{���]�R!�B�DLY�2���sRP�H_PK�E��2RETRIEt��2�b�5����FI�B� ����8� 2���0DBGLV�L�OGSIZ$C�K%TؑUy#u�D7�_��_T1@�EM�@C\1A����R��D�F�CHECKK�R�)P�0����@&�(b�LEc�" PA9�T(���P�C߰PN�����ARh�0������PO�BORMATTnaF�f1h���02�S��UXy`	���LB��4� { rEITCH���7�9PL)�AL?_ � $��XPRB�q� C,2D�!���+2�J3D���{ T�pPDCKyp���oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYLOYA��m�_1t�2t���J3AR��؀�x�֏�laTIA4��u5��6,2MOMCP@�����������0Bϐ�AD��������PUBk`R��;���;�������z4�` I$PI\Ds�oӓ1�yՕ�w�2�w�Z��I
��I��I���p����n���y�e`�9S|)bT�SPEED� G��(�Е��/���Е �`/�e�>��M��ЕSAMP�6V��/���ЕMO�@ 2@�A��QP���C��n� ����������LRf`kb`�ІE9h�EIN0 9��7S.В9
yxPy�GAMM%�S���D$GETH)bP�cD]��2
��IB�q�I�G$H�I(0;A��LRE�XPA8)LW VM8z)��tg���C5�CHKKp4]�0�I_��h` eT��n�q��eT�,���� �$^�� 1�iPI� RCH_D�313\��30LE�1�1\�o(�Y�7 �t�MSWFuL �M��SCRc��7�@�&��%n�f�SV���PB``�'��!�B�sS_SAV�&0ct5B3NO]�C \�C2^�0�mߗ�u� �a��u���u:e;��1���8��D�P����� ����)��b9�� e�GE�3��V�7���}Ml�� � ��YL��QNQS RlbfqXG�P�RR#@dCQp� �S:AW70��B�B[�CgR:AMxP�KCL�H���W�r��(1n�g�M�!o��� �F�P@}t$W P�u�P r��P5�R <�RC�R��%�6�`���� ��qsr X��O�D�qZ�Ug�ڐ>D�[ ��OM#w� J?\?n?�?�?��9�b"��2�L]�_��� |��X0��bf��qf@��q`�ڏgzf��Eڐ(�>j�"�ܰ��Fd�PB��PM�QU��� � 8L�Q�COU!5�QTH�I�HOQBpHYSfY�ES��qUE�`t�"�O���  �1P�@\�UN���C�f�O�� P���Vu��!����OGSRAƁcB2�O�t�VuITe �q:pINFO�����{�qcB��e�OI�r� (�@SLEQS��q���p�vgqS����{ 4L�ENABDR>Z�PTIONt���p��Q���)�GCF��G�$J�q^r�� R���U�g������_ED����ѓ �F��PK���E'NU߇وA�UT$1܅COPY������n�00MNx���PRUT8R� �Nx�OU���$G[rf�d�RGAkDJ���*�X_:@�բ$�����P��W��P��} ��)�}�[EX�YCDR|��NS.��F@r�LG�O�#�NYQ_FREQR�W� �#�h�TsLAe#������ �CRE� s��IF��sNA���%a�_Ge#STA�TUI`e#MAIL�����q t��������ELEM��� �/0<�FEASI?�B��n�ڢ�vA�]� � I�p��`Y!q]�t#A�ABM����E�p<�VΡY�BCASR�Z��S�UZ��0$q���RMS_TR;�qb  ���SY�	�ǡ��$����>C�Q`	� 2� _�TM�� ����̲�@ �A��)ǜ��i$DOU�s]$NLj���PR+@3���r�GRID�qM�BA�RS �TY@��O�TO�p��� Hp_"}�!����d�O�P/��� � �p�`P�OR�s��}���SReV��)����DI&0T����� #�	�#�U4!�5!�6!�7!�I8�e�F�2��Ep?$VALUt��%���ֱ��/��� !;�1�q�����(F_�AN�#�ғ�Rɀ|(���TOTAL��,S��PW�Il��REGEN�1�c�X��ks(��a���`T1R��R��_S� ��1ଃV�����⹂Z�E��p�q��Vr���7V_H��DA�S�����S_Y,1�R4�S�� AR�P2� >^�IG_SE	s��d��å_Zp��C_��~��ENHANC�a�� T ;�8������INT�.���@FPsİ_OVRsP�`p�`��Lv�҂o��7�}��Z�@�SSLG�AA�~�2 5�	��D��S�BĤ�DE�U�����T�E�P���� !�Y��
�J��$2�IL_MC�x r#_��`TQ�`��q���'�B5V�C�P_� 0ڽM�	V1�
V1��2�2�3�3
�4�4�
�!���`� � m�A�2IN~VIBP���1�U2�2�3�3�4�4�A@-�C2�p� MC_YFp+0�0L	1(1d���M50Id�%"FE� S`�R/�@�KEEP_HNA�DD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0�#i�.�#REM�"�$�P�½%�!�(U}�e�$�HPWD  �`#SBMSK|)G��qU2:�P	�COLLAB� �!K5��B�� ��g��pI�TI1{9p#>D� �,�@FLAP��$�SYN �<M�`C�6���UP_DL�YAA�ErDELAh�0ᐢY�`AD�Q�	��QSKIPN=E� ���XpOfPcNTv�A�0P_Xp �rG�p�RU@,G��:I +�:IB1:IG�9JT�9J@a�9Jn�9J{�9J9<���RA=s� X����4�%1�QB� N�FLIC�s�@J�Ux�H�LwNO_H�0X�"?��RITg��@�_PA�pG�Q�S ��^�U��W���LV�d�NGRLT �0_q��O�  " ��OS���T_JvA V	�A�PPR_WEIG=H�sJ4CH?pvT�OR��vT��LOO��]�+�tVJ�е�ғaA�Q�U�S�XOB'�L'�@aJ2P���7�X�T�<a43DP=`�Ԡ\"<a�q\!��RD�C��L� �рR"��R�`� �RV��j8r�b�RGE��*��cN�FLG�a�Z��ΒSPC�s�UM�_<`^2TH2N�H��P.a 1� mm`EF11��� lQ �!#� <�p3AT� g�S�&�Vr �p�tMq�Lr����HOMEwr�t2'r�-?Qcu�
�w3'r����(���w4'r�'�9��K�]�o����w5'r뀤���ȏڏ����w6'r�!�3�E�W�i�{�
�w7'r힟��ԟ(����w8'r��-� ?�Q�c�u��uS$0�q��p�� sF��`�la�!`P����0�`/���-�IO[M��I֠��*�POW=E�� ��0rZa*��� �5ވ�$DSB GNAL���0Cp���1�RS2323�� Ɍ~`��� / ICEQP��PEp��5PsIT����OPBx0ޣ�FLOW�@TR`vP��!U���CU�M��UXT�A��w�ERFAC�� Uv��kbSCH��'� tQ  _��>�f�Q$����OM���A�`T�P#UP%D7 A�ct�T��U�EX@�ȟ�U EFqA: X"�1RSPT�N����T ��PPaA�0o񩩕`EXP��IOS���)ԭ�_`���%��C�WR�A���ѩD�ag֕`ԦF�RIENDsaC2U�F7P����TOOLΫ�MYH C2LE�NGTH_VTE��I��Ӆ$S�E����UFINV�_���RGI��{QITI5B��X�v��-�G2-�G1@7�w�SG�X��_��UQQD=#���AS�Äd~C�`��q�� ��$$C/�S�`������ �  }��VERSI� ������5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����� ����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT��C��  ��DI�N�O�A�Dq�EXE��HPV_��AT�Qz
��LARM�RECOV ��RgLMDG �*�5�OLM?_IF *��`d�O�_�_�_�_j�_�'o9oKo]onm, 
��odb��o�o�o0�o^��$� z, �A   2D{�P�PINFO u[ �Vw��������`����� ��*��&�`�J���n�����DQ���� 
��.�@�R�d�v���𚟬���a
PPLI7CAT��?�P���`Ha�ndlingTo�ol 
� 
V�8.30P/40�Cpɔ_LI
8�83��ɕ$ME�
F0G�4�-
?
398�ɘ��%�z�
7�DC3�ɜ
�No+neɘVr���ɞ_@6d� ~Vq_ACTIVU���C죴�MOD�P���C�I��HGA�PON���O�UP�1*�� Ai�m����Қ_��6��1*�  �@��������Q����Կ�@�
���=�� ���5��Hʵl�K�HTTHKY_��/�M� SϹ���������%� 7ߑ�[�m�ߝߣߵ� ���������!�3�� W�i�{�������� ������/���S�e� w��������������� +�Oas� ������ '�K]o��� �����/#/}/ G/Y/k/�/�/�/�/�/ �/�/�/??y?C?U? g?�?�?�?�?�?�?�? �?	OOuO?OQOcO�O �O�O�O�O�O�O�O_ _q_;_M___}_�_�_��_�_�_�_kŭ�TO�p��
�DO_CL�EAN9��pcNM  !{衮o�o��o�o�o��DSP�DRYRwo��HI��m@�or��� ������&�8�J���MAXݐWdak�H�h�XWd�d��>�PLUGGW�Xg\d��PRC)pB�`E�kaS�Oǂ�2DtSEGF0�K � �+��o�or�����p�����%�LAPO b�x�� �2�D�V�h� z�������¯ԯ�+�TOTAL����+�_USENUO�\�� e�A�k­�RGD�ISPMMC.�2��C6�z�@@Dr\��OMpo�:�X�_S�TRING 1	~(�
�M!��S�
��_ITwEM1Ƕ  n� �����+�=�O�a� sυϗϩϻ����������'�9�I/�O SIGNAL���Tryou�t Modeȵ�Inpy�Simu�lateḏO�ut��OVE�RRLp = 10�0˲In cy�cl�̱Pro?g Abor��̱�u�Status�ʳ	Heartb�eatƷMH �Faul	��Aler�L�:�L�^�p����������� ScûSaտ��-�?� Q�c�u����������� ����);M_q��WOR.�û� �����+ =Oas��������//'.PO����M �6/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�?8�?�?H"DEVP.�0 d/�?O*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8_J_\_n_PALT	��Q�o_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o8�o�_GRIm�û 9q�_as��� ������'�9� K�]�o�������'�R	�݁Q����)� ;�M�_�q��������� ˟ݟ���%�7�I�ˏPREG�^���� [�����ͯ߯��� '�9�K�]�o�������෿ɿۿ�O��$A�RG_� D ?	����0���  	]$O�	[D�]D���O�e�#�SBN_�CONFIG �
0˃���}�C�II_SAVE � O�����#�T�CELLSETU�P 0�%  ?OME_IOO�O�%MOV_H������REP��J��UTOBACK�����FRwA:\o� Q�,o���'`��o����� ��  f�o�����*�!�3�`��Ԉ��f���� ������o�{��&�8� J�\�n���������� ��������"4FX j|�������끁  ��_�i�_\ATBCK�CTL.TMP �6.VD GIF? .TP D_8q��NLQ���.f�INI�P�Օ��c�MESSAG�����8��ODEC_D����z��O�0��c�PAUSM!!��0� (783�U/g+(Od/�/ x/�/�/�/�/�/�/? ??P?>?t?1�0$: ?TSK  @-��<T�f�UPDT���d�0
&XWZD�_ENB����6S�TA�0��5"�XI�S��UNT 2|0Ž� � 	�0���b ��� ���pv�~^io�:UA M   �D����uK�Oo�}C/�#���쀴şO� _�O$_�7AMET�߀2CMPTA@��\w@^��@��Ã@q�@W��%@C
]5�5�~4�15�*u5� �4���4�ff8]�SCRDCFG }1�6��	��Ź�_�_oo (o:oLo��o�Q���_ �o�o�o�o�o�o]o �o>Pbt���o9�i�GR<@M/��s/NA�/�	�i��v_ED�1��Y� 
 �%{-5EDT-��'�GETDATAU�o�9��?�j�H�o�f�\��A�^�  ���2�0&�!�E���:IB����~�ŏ׏m����3 ��&۔��D��ߟJ� ����9�ǟ�4��� ϯ�(����]�o�����5N������(��w��)�;�ѿ_��6 ϊ�gϮ�(�CϮ���ϝ�+��7��V�3� z�(��z�����i���B�8��&���~�]����F�ߟ�5����9~������]����`Y�k�����CR� !ߖ���W�q���#�5����Y��p$�NO_D�EL��rGE_U�NUSE��tIG�ALLOW 1���(*S�YSTEM*S�	$SERV_G�R�V� : REGƟ$�\� NU�M�
��PMU|B ULAYNP�\PMPA�L�CYC10�#6 $\UL�SU�8:!��Lr�BOXOR=I�CUR_���PMCNV��10L�T4�DLI�0��	�� ��BN/`/r/�/�/�/�/�/���pLAL_?OUT �;����qWD_ABOR�=f�q;0ITR_�RTN�7�o	;0NgONS�0�6 
H�CCFS_UTI�L #<�5CC�_@6A 2#; h ?�?�?O#O6]�CE_OPTIO�c8qF@RI'A_Ic f5Y@�25�0F�Q�=2qz&}�A_LIM��2.� �K �&]B��KXK QY�2O�Q��B�r
�qFK Q5T1)T�R�H�_:JF_P�ARAMGP 1�<g^&S�_�_��_�_�VC�  C�d�`�o!o`U�`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?퀗2HE ONFqI� E?�aG_P�;1#; �� �o1CUgy��aKPAUS�19�yC ,��� ������	�C� -�g�Q�w���������hя���rO�A�O��H�LLECT_b�B�IPV6�EN. �QF�3�NDE>�� �G�712�34567890���sB�TR����%
 H�/%)���� ���W���0�B���f� x���㯮���ү+��� ��s�>�P�b����� �����ο��K��@(�:ϓ�^�|��B!F�� �I|�IO ##��<U%e6߰'�9�K���TR�P2$��(9X�t�Y޼`�%�̓ڥH��_M[OR�3&�=�K XB��a��A �$��H�6�l�~���D~S��'�=�r_A?�a�a`��K K��R�d�P��)F�ha�A-�_�'�9�%
� k��G� ��%Z�%���`K c.�P�DB��+���c?pmidbg��	��`:�K ` ��QU��p��N � �K ���)X���]�K �sX<�^�K �s�g�$� �sf�l�q��ud�1:��:J��DE�F *ۈ��)��c�buf.t�xt����_L�64FIX , ������l/[Y/�/}/ �/�/�/�/
?�/.?@? ?d?v?U?�?�?�?�?��?�?,/>#_E -���<2ODOVOhOXzO�O6&IM��.o�=YU>���d�
�6IMC��2/���ñdU�C��20�M��QT:Uw�Cz  B��i�A���A����A@��B3��*CG�B<�=w�i�B.���B���B����B�$�D�%�B���ezVC�q��C�v�C�n��D-lE\D�n�j�0�Bl9"��22o�D|���0�0 GC�ZC����
�xObfi�D4cdv`D��`�/�`v`s]E�D �D�` E4��F*� Ec���FC��u[F����E��fE��f�Fކ3FY��F�P3�Z��@��33 ;��>LS���Aw�n,a@�0@e�5Y���a����`A��w�=�`<#����
��?�ozJR�SMOFST �(�,bIT1��D2 @3��
д����a���;��bw?���<�M�N/TEST�1O�CER@�4��>VC5`#A�w�Ia+a�aOR�I`CTPB�U�C��`4���r�0:d�����qI?�5���qT_�PROG ��
�%$/ˏ�t���NUSER  �U������KEY_TBL  �����#a��	
��� !"#$%&�'()*+,-.�/��:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s������LCK�x
����STAT/���s_AUTO_D�O �	�c�IN?DT_ENBP���1Rpqn�`�T2�����STOr`���XCΔ� 26���8�
SONY XC�-56�"b�����@��F( А{�HR50w����>�P�7b�t�ACff����ֿ� Ŀ ����C�U�0�yϋ� fϯ��Ϝ���������-ߜ�TRL��LE�TEͦ ��T_�SCREEN }��kcs�����U�MMENU� 17�� < ܹ���w������ ���K�"�4��X�j� ������������5� ��k�B�T�z����� ����������. g>P�t��� ���Q(: �^p����/ ��;//$/J/�/Z/ l/�/�/�/�/�/�/�/ 7?? ?m?D?V?�?z? �?�?�?�?�?!O�?
O WO.O@OfO�OvO�O�O�(y��REG 8�y����`�M�ߎ�_MANUAL��k�DBCO��RI�GY�9�DBG_E7RRL��9�ۉqa��_�_�_ ^Q�NUMLI�pϡꘀd
�
^QPXW�ORK 1:����_5oGoYoko}oӍD�BTB_N� ;T�����ADB_AWAYfS��qGCP 
�=�p�f_AL�pR��bBbRY�[�
�WX_�PW 1<{y�n�,��%oc�P��h_M&��ISO��k@L��s�ONTIMX��&
���vy
��2sMOTNEND��1tRECORD ;1B�� ���sG�O�]�K��{�b ��������V�Ǐ�]� ���6�H�Z����� ����#�؟������ 2���V�şz������� �ԯC���g��.�@� R���v�寚�	���п ���c�χ�#ϫ�`� rτϖ�Ϻ�)ϳ�M� ��&�8ߧ�\�G�U� ��߶�����I������4�� �p7�n�� �ߤ��������� "���F�1���|���� ����[�����i����BTf���bTO�LERENC�dB��'r�`L��^PC�SS_CCSCB' 3C>y�`IP�t}�~�<�_ `r�K�����/�{��5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O �O�O�O�O�O_�~�kLL� D��&q�ET�c�a C�[C�`ZP^r_ +A� p� �sp���QGPt[	 A�p�Q�_�[? �_�[4oU�p��p�pSB�V�c�(a�P�Woio{h+�o�X0�o�oY��[	r��hLU�NH���8yn�d���2ܘ��c���aD@VB���|�G����+��K�  �otGhXGr�So����eB   /=��Ͷa>�tYB�� �pC�p�q�aA"�H�S�Q-��q����ud�v�����AfP� ` 0���DX^P��p@�a
�Q�XTHQ����a DaW>� �a9P��b �e:�L�^�h�Hc�́PQ�RFQ�PU�z� ֟�o\^��-�?��`c�u����zCz㎉ů�b2�Щ�RDw��(��}�ҁ� ��S̡0��]�0�.��@���EQ�p��F� X�ѿUҁп�VS���NSTCY 1)E��]�ڿ�� K�]�oρϓϥϷ��� �������#�5�G�Y��k�}ߏߒ��DEV�ICE 1F5� MZ�۶a��	� � �?�6�c���	{䰟����_HNDGD G5�VP���R�LS 2H�ݠ�� /�A�S�e�w����� Z�PARAM I��FgHe�RBT� 2K��8р<X��WPpC�C��,`E¢P�Z�z��}%{�C*  �2��jMTLU,`"nPB, s��M� }�0gT�g��
B��!�bcy�[2Dc hz����/�x�/gT#I%D���C�` b!�R��A���A,��B_d��A��P��_cC4kP�!2�C��$|Ɓ�]�ffA�À_��B�� �| a���/�/�T (�P 54a5�}%/7/d? /M?_?q?�?�?�?�? �?O�?OO%O7OIO �OmOO�O�O�O�O�O �O�OJ_!_3_�_�_3 �_�_�_�_�_o�_(o oLo^oЁ=?k_IoS_ �o�o�o�o�o�o�o #5G�k}� ������H�� 1�~�U�g�y�ƏAo� Տ���2�D�/�h�S� ��go����ԟ����ϟ ���R�)�;���_� q����������ݯ� <��%�7�I�[�m��� ������}�&��J� 5�n�YϒϤϏ��ϣ� ѿ������F��/� Aߎ�e�w��ߛ߭��� ������B��+�x�O� a����������� ,���%�b�M���q��� ������������ L#5�Yk}� �� ��6 1CUg���� ����	//h/�� �/w/�/�/�/�/�/
? �/.?@?I/[/1/_? q?�?�?�?�?�?�?�? OO%OrOIO[O�OO �O�O�O�O�O&_�O_ \_3_E_W_�_?�_�_ �_�_�_"ooFo1ojo E?s_�_�om_�o�o�o �o�o0f=O a������� ���b�9�K���o� ��Ώ��[o��(���L�7�I���m�������$DCSS_SL�AVE L����ё~��_4D  љ���CFG M�ѕ�������FRA:\Đ�L-�%04d.C�SV��  }�� m���A i�CHq�z������|�����  �����Ρޯx̩ˡҐ-��*�����_CRC_OU/T N�������_FSI ?>њ ���� k�}�������ſ׿ � ����H�C�U�gϐ� �ϝϯ��������� � �-�?�h�c�u߇߰� �߽���������@� ;�M�_������� ��������%�7�`� [�m������������ ����83EW� {������ /XSew� ������/0/ +/=/O/x/s/�/�/�/ �/�/�/???'?P? K?]?o?�?�?�?�?�? �?�?�?(O#O5OGOpO kO}O�O�O�O�O�O _ �O__H_C_U_g_�_ �_�_�_�_�_�_�_ o o-o?ohocouo�o�o �o�o�o�o�o@ ;M_����� �����%�7�`� [�m��������Ǐ�� ����8�3�E�W��� {�����ȟß՟�� ��/�X�S�e�w��� �����������0� +�=�O�x�s������� ��Ϳ߿���'�P� K�]�oϘϓϥϷ��� ������(�#�5�G�p� k�}ߏ߸߳����� � ����H�C�U�g�� ������������ � �-�?�h�c�u����� ����������@ ;M_����� ���%7` [m����� ��/8/3/E/W/�/ {/�/�/�/�/�/�/? ??/?X?S?e?w?�? �?�?�?�?�?�?O0O +O=OOOxOsO�O�O�O��O�C�$DCS_�C_FSO ?�����A? P �O�O _?_:_L_^_�_�_�_ �_�_�_�_�_oo$o 6o_oZolo~o�o�o�o �o�o�o�o72D Vz����� ��
��.�W�R�d� v������������ �/�*�<�N�w�r��� ������̟ޟ��� &�O�J�\�n������� ��߯گ���'�"�4� F�o�j�|�������Ŀ ֿ������G�B�TϾ�OC_RPI�N _jϳ����ς��O��`��1�Z�U��NSL��@&�h߱��������� "��/�A�j�e�w�� ������������ B�=�O�a��������� ��������'9 b]o����� ���:5GY �}������ ///1/Z/U/g/y/ �/�/�/�/�/�/�/	? 2?-???Q?z?u?��� �߆?�?�?�?OO@O ;OMO_O�O�O�O�O�O �O�O�O__%_7_`_ [_m__�_�_�_�_�_ �_�_o8o3oEoWo�o {o�o�o�o�o�o�o /XSew� �������0� +�=�O�x�s������� ��͏ߏ���'�P��K�]�o����� �PR�E_CHK P�۪�A ��,�8�2��� �	 8�9�K��� +�q���a�������ݯ �ͯ�%��I�[�9� ���o���ǿ��׿�� �)�3�E��i�{�Y� �ϱϏ��������� ��-�S�1�c߉�g�y� ���߯����!�+�=� ��a�s�Q����� ���������K�]� ;�����q��������� ����#5�Ak {����� �CU3y�i ������/-/ G/c/u/S/�/�/�/ �/�/�/??�/;?M? +?q?�?a?�?�?�?�? �?�?�?%O?/Q/[OmO O�O�O�O�O�O�O�O _�O3_E_#_U_{_Y_ �_�_�_�_�_�_�_o /ooSoeoGO�o�o=o �o�o�o�o�o= -s�c��� ����'��K�]� woi���5���ɏ���� ����5�G�%�k�}� [�������ן�ǟ� ���C�U�o�A����� {���ӯ����	��-� ?��c�u�S������� Ͽ῿�����'�M� +�=σϕ�w�����m� �����%�7��[�m� K�}ߣ߁߳��߷��� �!���E�W�5�{�� �ϱ���e�������	� /��?�e�C�U����� ����������= O-s����] ����'9] oM������ �/�5/G/%/k/}/ [/�/�/��/�/�/�/ ?1??U?g?E?�?�? {?�?�?�?�?	O�?O ?OOOOuOSOeO�O�O �/�O�O�O_)__M_ __=_�_�_s_�_�_�_ �_o�_�_7oIo'omo o]o�o�o�O�o�o�o !�o1W5g� k}������ /�A��e�w�U����� ��я��o����	� O�a�?�����u���͟ �����'�9��]� o�M���������ۯ�� ǯ�#�ůG�Y�7�}� ��m���ſ�����ٿ �1��A�g�E�wϝ� {ύ�������	�߽� ?�Q�/�u߇�e߽߫� ���������)��� _�q�O�������� ������7�I���Y� �]������������� ��!3WiG� �}����%� A�1w�g� �����/+/	/ O/a/?/�/�/u/�/�/ �/�/?�/9?K?�/ o?�?_?�?�?�?�?�? �?O#OOGOYO7OiO �OmO�O�O�O�O�O_ �O1_C_%?g_y__�_ �_�_�_�_�_�_o�_ +oQo/oAo�o�owo�o �o�o�o�o);U_ _q����� ���%��I�[�9� ���o���Ǐ����� ۏ!�3�M?�i��Y� ������՟�ş�� ��A�S�1�w���g��� �������ӯ�+�=���$DCS_SG�N QK�c���7m� 12�-FEB-19 �15:15   |O�l�4-JANt��08:38}������ N.D������������h�x�,rWf*σ��^M��  O�VE�RSION �[�V3.5.�13�EFLOG�IC 1RK���  	����P�?�P�N�!�P�ROG_ENB � ��6Ù�o�U?LSE  TŇ��!�_ACCLI�M����Ö���WRSTJNT��c��K�EMO�x̘��� ���INIT S.�G�Z����OPT_SL ?�	,��
 	�R575��Y�74j^�6_�7_�50��1��2_�@ȭ��<�TO  Hݷ���V�DEX��d�c����PATHw A[�A\��g�y��HCP_CLNTID ?��6� @ȸ�����IAG_GRP� 2XK� ,`����� �9�$�]�H������1234567�890����S�� |�������!�� ��H���;�dC�S���6�� ���.�R v�f��H�� //�</N/�"/p/ �/t/�/�/V/h/�/? &??J?\?�/l?B?�? �?�?�?�?v?O�?4O FO$OjO|OOE��O y��O�O_�O2_��_�T_y_d_�_,
�B^ 4�_�_~_`Oo�O &oLo^oI��Tjo�o.o �o�o�o�o �O'�_ K6H�l��� ����#��G�2�`k�V���B]�?�BS��;�.����� �D|Ρ@�YD�!���Ƈ�����(��L�B\ډ�4?  6(�:��� 6��������؟����CT_CONFI/G Y��Ӛ��egU���STBF_TTS�ǁ
��b����Û�u��O�MAU��|��M_SW_CF6�Z���  �OCVI�EW��[ɭ������-�?�Q�c�u� G�	�����¿Կ��� ���.�@�R�d�v�� �ϬϾ�������ߕ� *�<�N�`�r߄�ߨ� ����������&�8� J�\�n���!���� ���������4�F�X��j�|����RC£\�e��!*�B^�������C2g{�SB�L_FAULT �]��ި�GPM�SKk��*�TDI�AG ^:�ա�I��UD1:� 6789012�345�G�BSP �-?Qcu�� �����//)/P;/M/tJ��
@q���/$�TRECP��

��/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O�BOi/{/xO�/UMP_OPTIONk����ATR¢l��	λEPMEj��OY_�TEMP  ß��3B�J�P�9AP�DUNI��m��Q��YN_BRK� _ɩ�EMG?DI_STA"U�alQSUNC_S1`ɫ� �FO�_�_�^
�^dpOoo%o7oIo [omoo�o�o�o�o�o �o�o!3EWi {�E�����y�Q ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d��z� ������˟���� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i���������ÿ ݟ�����/�A�S� e�wωϛϭϿ����� ����+�=�O�a�{� iߗߩ߻�տ����� �'�9�K�]�o��� ������������#� 5�G�Y�s߅ߏ����� i�������1C Ugy����� ��	-?Qk� }��������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?u?�?�? �?��?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ m?w_�_�_�_�?�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9Ke_W�� ��_�_����#� 5�G�Y�k�}������� ŏ׏�����1�C� ]oy��������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;���g�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�_�i�{ߍߟ߹��� ��������/�A�S� e�w��������� ����+�=�W�E�s� �����ߧ������� '9K]o�� ������# 5O�a�k}�E�� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-?GYc? u?�?�?��?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_Q?[_m__�_�? �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/I_S ew��_���� ���+�=�O�a�s� ��������͏ߏ�� �'�A3�]�o���� ���ɟ۟����#� 5�G�Y�k�}������� ůׯ�����9�K� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� �ߑ�C�M�_�q߃� ���߹��������� %�7�I�[�m���� �����������!�;� E�W�i�{��ߟ����� ������/AS ew������ �3�!Oas ��������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?+ =G?Y?k?!?��?�? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�O �O�O	_#?5??_Q_c_ u_�?�_�_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o -_7I[m�_�� ������!�3� E�W�i�{�������Ï Տ����%/�A�S� e�q�������џ� ����+�=�O�a�s� ��������ͯ߯�� ��9�K�]�w����� ����ɿۿ����#� 5�G�Y�k�}Ϗϡϳ� ���������'�1�C� U�g߁��ߝ߯����� ����	��-�?�Q�c� u����������� m��)�;�M�_�y߃� ������������ %7I[m�� ������!3 EWq�{���� ���////A/S/ e/w/�/�/�/�/�/�/ �/�/+?=?O?i_? �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O��O�O�O�O�O? ��$ENETMOD�E 1aj5��  0�054_F[PRR�OR_PROG %#Z%6�_�YdU�TABLE  #[t?�_�_�_gdR�SEV_NUM �2R  ��-Q)`dQ_AUTO_ENB  PU�+SaT_NO>a �b#[EQ(b  �*��`��`��`��`4`+�`�o�o�oZd�HIS%c1+PSk_�ALM 1c#[� �4�l0+ �o;M_q���o�_b``  #[�aFR�zPTCP_�VER !#Z!��_�$EXTLO�G_REQ�f�Qi,�SIZ5�'�SkTKR�oe�)��TOL  1D�z�b�A '�_BWD�p��Hf��D�w_DI�� dj5�SdDT1KRņS�TEPя�P��O�P_DOt�QFA�CTORY_TU�N�gd<�DR_G�RP 1e#YNad� 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ�ԟ� ��1��U�@�y�d�v������ӯ����LW
 Jg��,��t�ۯ�j�U���y�B_�  B୰����$  A@��s�@UUUӾ��������E�� E�`F?@ F�5U/�,���L���M���Jk�Lzp��JP��Fg�=f�?�  s���9�Y9}��9��8j
��6��6�;���m���y� �!� �� Q�(������[FEATURE� fj5��JQ�HandlingTool �� "
PE�nglish D�ictionar�y�def.�4D St�ar�d�  
! h�Analog� I/OI�  !�
IX�gle _ShiftI�d��X�uto Sof�tware Up�date  rt� sѓ�matic Backupӿ3\st��g�round Ed�it��fd
�Camera�`�Fd�e��Cnr�RndIm���3��Common �calib UI��� Ethe�n���"�Monito�r�LOAD8�t�r�Reliab�y�O�ENS�Dat�a Acquis�>��m.fdp�iagnos��]�i��Document? VieweJ���870p�ual� Check S�afety*� c�y� �hanced7 Us��Fr�����C �xt. D�IO :�fi�� �m8���end��ErrI�L��S�������s  t Pa��r[�� ���J�944FCT�N Menu��v�e�M� J9l�TPw InT�fac{�_  744��G���p Mask E�xc��g�� R8�5�T��Prox�y Sv��  1�5 J�igh-wSpe��Ski
� R738Г��mmunic��o{ns�S R7���urr�T�d�022���aю�conne�ct 2� J5އ�Incr��st�ru,Қ�2 R�KAREL C�md. L��ua޷�R860hRu�n-Ti��Env�L�oa��KU�el� +��s��S/W�ѹ�7�Licen�se���rodu�� ogBook(System)��AD pMA�CROs,��/Ogffs��2�NDs�#MH�� �����MMRC�?��OR�DE� echSt�op��t? � 8�4fMi$�|� 13dx��]е�׏���Modz�witchI�VP��?��. sv��2O�ptm�8�2��fCil��I ��2g� 4 !+ult�i-T�����;��PCM funY�Po|���4$�^b&Regi� r .�Pri��FK+7����g Num S[elW  F�#>�� Adju����60.��%|� fye���&tatu�!�$6���%��  9� J6RDM� Robot)�s�cove2� 56�1��RemU�n�@� 8 (S�F3Servo�ҩ��)SNPX yb�I�\dcs�0�}�Libr1��H'� �5� f�0���58��So� t�r�ssag4%G 91�p ��&�0���p/I��  �(ig TMILI�B(MӋ�Firm�����gd7���s�A�cc����0�XAT9X�Heln��*L�R"1��Spa�c�Arquz�im'ulaH��� Q���7Tou�Pa��I���T��c��&��e�v. f.svUSB po���"�iP�a��  �r"1Unexcept��`0i$/���׷H59� VC&�r��[6���P{��R�cJPRIN�V�; �d T@�TSP OCSUI�� r�[�XC��#Web sPl6�%d -c�1R�@4d�����I�R66?0FV�L�!�FVGridK1play C�lh@��,��5RiR�R.@���?R-35iA�>��Ascii���"���� 51f�cUspl� � (T����S��@rityAvoidM �`6��CE��rk�gCol%�@�GuF� 5P��j}P����
 �B�L�t� 120
C C� o�І!J��P"��y��� o=q�b� @DCS b ./��c��O��q��`Ң; ���qckpa3boE4�DH@�O�TШ�main N���1.�H��an.���A> aB!FRL�M���!i ���MIo Dev�  (�1�� h8j��spi�JP��� �@��Ae1/Ⱦr���!hP� M�-2� i��߂^0i��p6�PC�� � iA/'�Pas�swo�qT�RO#S 4����qeda�;SN��Cli�����G6x Ar�� 4�7�!���5s�DE�R��Tsup>Rt<�I�7 (M�a�T�2DV�
�3D Tri-���&���_8;�
�A�@Deaf?����Ba: odeRe p 4t0@��e�+�V�st�64MB DRA�M�h86΢FsRO֫0�Arc� GvisI�ԙ�n�՞7| ), �b�Hgeal�wJ�\h��OCell`��p� �sh[��� Kqw�c� - �v��бp	VCv�tyy�s��"Ѐ6�ut@��v�m���xs ���TD_0��J�m�`� 2��a[�>R t{si�MAILYk��/F2�h��ࠛ 90 H��F02]�eq�P5'���T1C��5����FC��U�=F9�GigEH�S�qt�0/A� if�!�2��boF�driz=c �OLF�qS����" H5k��OPT ��49pf8���cro6���@��l�ApA�S�yn.(RSS)# 1L�\1y�rH�L�� (2x5�5�d�pCqVx9����est�$�SР��> \pϐSuSF�e$�tex�D o���A�	� BqP���a�(R00�QGirt��:���2)��D��1�e�VKb@l/ Bui, n��W�APLf��0��Va�kT�XCGM��D��qL����[CRG&La�YBU��YKf�L��pf��k�\sm��ZTAf�@�О�Bf2�и��V#�s���2� r���CB����
f���WE��!��
���T�p��D"T�&4 Y�V�`���EH����
�61Z��
�R=2�
�E (Np��F�V�PK�B���#��Gf1`?�G���H�р?I2�e ����LD�L��N��7\s@����`���M��del�a<,��2�M�� "L[P��`?��_�%�����S��-�F�TSO�W�J;57��VGF�|�wVP2֥ 5\b� `0&�cV:���T;qT� �<�ce,?�VPD��$
�T;F��DI)�<IN�a\so<��a-�6Jc6s6�4L�M�V91R�h���Tri�� ���5�` �f�@�������P
� ����`���Img PH�[ll��I/A  VP"�S��U�Ow��!�%S�Skastdpn�)ǲt�� SWIM�EST�BFe�00��-Q� �_�PB�_��Rued�_�T�!��_�S ��_bH57�3o2c2��-oNbJ!5N�Iojb)�Cdo�cxE��o�_�lp��o�T dP�o�c�B�or�2�.rٱ(Jsp�EfrS�Eo�f1�}�r3 9RGoeELS��sL����s�����B`	��S\ $�F�ryz&�ftl�o~�g�o�� �������?�����AP  �n�&�"�l � �T�@<�^��Y��e��u8Z���alib ��Γ��ɟ3���埿�3\v ��e\c�6��Z�f�T�v�R V�W���8S��UJ91`����i�ů[c91+o�w8���847 �:��A4�j��Q��tx6�m���vrc.��`��HR���ot�0�ݿ��  ��8�ޯ�460�>eS0L�97���U�Є���60.� g�н�+� �'�ܠ�Ϻ�8co��DM߱U"������2�pi�߲T! ��na;�� ���u%��ⅰI��loR�0d��1a59gϱ�L����95�ϔ�R����1��?��o�#��1�A�/���vt{�UWaeǟ���ￇ73[�r��7�ρ�C W&��62K�=fR���8��������d����2�ڔ����@��@" "http �����t7 �� vg R7��78�����4�� ��TTP�T�#	��ePC�V4/v߀�j�Q�F�a7��$N�0�/2�r�IO�)/;/M/6.s�v3�64i�oS�l? torah?*�|`�?��AM/�?
??.?80�k/��1 JO��� ,O�tro���[P��OB4c.K?�g'��)�24g?�� (B��Od�\iOA5s1b�?U_�?vi�/i��/�/Wn��`�o%�Fo�4l�$of��o�XF I)xo�cmp�\7��mp���du�C��lh����o(A �_Bt� �o]6P��m�`I?�w�@���naO��4*O0wi�%P�?"�bsg?�]7�HYEM���8woVJ�/fե11?o��DMs&�BC��7J�\����(�52�XFa A�P�ڟ<�v�`/şa�qs����/Of$��1�9�V�RK���ph�քH5�+�=�IN/¤Sk1iW�/�IF��_�%��fs�I�O�	l����"<𜿚$�`����\jԿz5bO�v'rouς�3(�ΤH (DϮ��?sG�� |��F�Ou�������D)O��*�3P$�FӀ��k��ϻ���럴� ��PL��ʿ��pbo�x�ߦebo���SIh �>�R.�0wT{����fx6��P���D��3��#_I\m$;YEe�OԆM�hx�W�=Ete,���dc#t\���O$kR�������Xm*���ro`3��D�l�j9���V'�  FC ���|@�ք f?6�KARE0�_�~ c(Kh��.cf����WpoO�_K�u�p��a���H/j#-g Eqd/�84���$qu�o��/ o2o�?Vo<�7C�)�s�N�JԆ�|?�3l\s�y�?�40�?Τwi0o�u]?�w58�?,FÀ$OJ�
?Ԇ"i$o�!�V��u&A��3PR�ߩ5, s��v�1\  �H552B�Q21|p0R78P�510.R0  �nel J6�14Ҡ/W�ATUP��d8P5�45*�H8R6��9�VCAM�q9�7PCRImP\1tPU�IF�C8Q28  ingsQy0��4P P�63P @P PSC�H��DOCV8ڀD �PCSU���0�8Q0=PqpVE�IOCr��� P54�Pupd�PR69�aP���PSET�ptC\hPQ`Qt�8P7`Q~�!MASK��~(PPRXY���R7B#POCO _ \pppb36����PR�Q��b1Pd6�0Q$cJ539.eH�sb��vLCH�-`(�OPLG�q\bPQ0]`��P�(`HCR��4`S�aund�PMCS�IP`e0aPle5=Ps�p(`DSW� �  q�Pb0`�aPa��(`PR�Q`Tq�RE`(Poa60�1P<cPCM�PHcR=0@q\j23b�V�`E`�S`UPvis�P`E` c�`UPcPsRS	a�bJ69E`�sFRDmPsRM;CN:eH931PHc�SNBARa�rHLB�USM�qc�Pg;52�fHTCIP0cTMIL�e"P�`e�J �PA�PdSTP�TX6p967PTEL�p��P�`�`
Q8P8$Q48>a"PPX��8P95�P`[�95�qqbUEC-`F
PUFRmPfahQ�CmP90ZQVCO��`@PVIP%�5�37sQSUIzVS9X�P�SWEBIP�SwHTTIPthrQ#62aP�!tPG���c�IG؁�`c�PG�S�eIRC%��cH76�P�e Q�Q|�9Ror��R51P s�:P�P,t53=P8u8=Py�C�Q6]`�b��PI��q52]`sJ�56E`s���PDsC�L�qPt5�\rdf�q75UP cR8��r�u5P sR55]` ,s� P8s��P�`CP��PP�SJ77P0\o�6��cRPP�cR6�ap�`�QtafT�79P`�64�Pfd87]`�d90P@0c��=P,���5�9ta�T91P� ��1P�(S���Qpai�P0]6=P- C�PF��T	���!aLP PTS\�pL�CAB%�I �БIQ` ;�H�UPP�aintPMS�Pap��D�IP|�STY%�ot\patPTO�pb�P�PLSR76�`b�5�Q��WaNN�P7aic�qNNE`��ORS�`�cR68�1Pint'�FCBD�P(�6x�-W`M�r���!(`OBQ`pl�ug�`L�aot ��`OPI-���PS\PZ�PPG�Q7�`�73ΒPRQa�d�RL��(Sp��PS��n�@�E`��� �PTS-��� W��P�`apwp�`��P`cFVR�P�lcV3D%�l�PB�VI�SAPL�Pc�yc+PAPV1�p�a_�CCGIP -� U��L�Prog�+PCCR�`�ԁB��P �PԁK=�"L��P��p��(h�<�P���h�̱�@g�Bـ�
TX�%���CT�C�ptp��2��P927"0ҝPs2�Qbv��TC-�rmt;�6	`#1ΒTC9`Hc�CTE�Perj�E.IPp.p/�E�P�c\��I�use��Fـ�vrv�F%���TG��P� CP��%�d -�h�H-�Tra�PC�TI�p��TL� TRS���p�@נ���IP�PTh�M%�le�xsQTMQ`ver, �p�SC:���F���Pv\e�PF�IPS�V"+�H�$cj�ـtr�aCTW-���CP�VGF-��SVP2�mPv\fx���pc��b��e��bVP4�f�x_m��-��SVP�D-��SVPF�P_Kmo�`V� cV���t\��LmPoveq4��-�sVPR��\|�tPV�Qe5.W`V6�*u"��P}�o`8���`��CVK��N�IIP��CV����I{PN9�Gene�� �D��D�R�D���� � ��f谔�pos�.��inal��n���DeR���`��d̔P��omB���onA,���R�D�R��\���TXf��D$b��omp�� "N��P���m���! ��=C�-f����=FXU8�����g F��(��Dt II��r�D��u�� "����Cx_ui X������f2��h	Cral2��D,r9ui�|Ԣ� it2c��0co��e"���{�ا(.)� ����� ���� IQnQ ��I[ ��_=� wo��,bD�� ��|G{G� ������4 �e�� vʷ� ��{&� 2��Z �uz������� ��TW&q~�q 5�׷&�o{? ;0�� � �2� �yݻ ���W&�{�� ?�3� �A��e�/>� �\�3&T���� 77߸ ����� ����� ֵ��&���8 �l1��S{�) ���d �*J� F's� ~��� 6:�0� ��,��s��- Q�v�� ��� �,{�T �ZBLx6����6 ��6�;��Par ���s>�E��j�6dsq��F  �������ЁDhel����<�ti-S�� �Ob��Dbcf�O������t OFT��P <A�_�V�ZI��D���V\�qWS��= odtle�Ean��(bzd��titv��Z�z�Ez XWO� H6�6���5{ H�6H691�E14܀TofkstF�. Y682�4�`�f7804�E91�g�`y30oBkmon_�E�eݱ�� qlm���0 J�fh��B��_  ZDTfL�0�f(P7�Eck�lKV� �6|��D858��ّ�m\b����xo�k�ktq��g�2.g���yLbk�LVts��IF�b�k������Id I/f��GR� �han�L��Vy��%���%ere�����i�o�� ac�- �A�n�h���cueACl�_�^ir���)�g��	.�@�& G<��R630���p� v�p�&H�f��un��R57v�OJ�avG�`Y��owc��-ASF��O0��7���SM������
af��ra)fLa�vl�\
F c�w a���?VXp�oV �30��NT "L�FFM��=�����yh	a�G-�w�� �m2.�,�t���̹�6ԯ��s�d_�MC'V����D����fslm�i�sc.  �H5522��2�1&dc.pR�78����0�7�08J614�Vip AT�Uu�@�OL�545�ҴINTL�6�t8 (VCA����sseCR1I��ȑ��UI���r7t\rL�28g�зNRE��.f,�6q3!��,�SCH�d{ Ek�DOCV��D�p��C,�<�L�0Q�wisp��EIO���xE,�54����9ށ�2\sl,�SE�T���lр�lt2��J7�ՌM�ASK��̀P'RXY҇��7��зOCO��J6l�3x�l�� (SVl��A�H�L�@Օ��53�9Rsv���#1κ�LCH���OP�LGf�outl�0���D��HCR
s�vg��S@�h��C1Sa�!�{�50��D��l�5!�lQ��DSWº�S����̀��OP4����7��PR���yL�ұ�(Sgd����PCM���R0 \s��5P՝���a0���n�q� AJ��1��N�q�2��PR�Sa���69�� (AuFRD��<���RMCN����93A�ɐCS�NBA�F9� HL	B��� M��4����h�2A�95z�HTyCaԈ�TMIL6��j95,��857�.,PA1�ito޻�TPTXҴ JNK�TEL��piL��� XpL�80�I)���.�!��P;�J95��s "N���H��UEC��7\csF�FR��<Q��C��w57\{VCOa�,,���IP1jH��wSUI�	CSX1�>�AWEBa���HTTa�8�R62���m`��GP%�I�G %tutKIP�GSj�| RC1_;me�H76��7P�ws_+�?x�wR51�\iw��N���H�53!��wrL�8!�h�R66�� H���Ԡ���@;J56��1���N0���9�j��L���R5(`%�A|�5q�r�`,�18 5��{165!��@��"5��H84!�2!9��0��PJ���wn B[�J77!���R6�5h3n���y36P��3R6��-`;�� Ԩ@��exe�KJ87��#J90!�stu+�~@!䷬��k90�k�op�B����@!�p�@|BA�g*�n@!��QF��06!�@[�F�F�aP�6��́,�TS�� NC[�CAB�$iͰl1I��R7���@q�y�CMS.1�rog+QM�� ��� TY$x�CTOa�nv\+��1�(�:,�6�con�~0v��15��JNN�%�e:��P��9ORS�%x���8A�815.[�FCBaUnZQ�P�!��p{��CMOB6��"G��OL��x�wOPI�$\lr[��SŠ�T	D7�U��C7PRQR9RL��ӁS�V�~`���K�ETS�$1��0���3��Ԩ�FVR1�L�ZQV3D$ ���B�Va�SAPL1�C�LN[�PV��	rCcCGaԙ��CL��3CCRA�n "�W!B�H�CSKQn\0�p��)�0CTPn�ЌQe��\�p!$bCt�aT0U�pCTC�yЋR�C1�1 (�s��t�rl,�r��
TXv��TCaerrm�r��MC"�s��#C�TE��nrr�RE�a�XPj�^��rm�c�^�a"�P�QFp!$���$p "�rYG1�tTG$c8�r�QH�$SCTI�w! s��CTLqd�ACK�Rp)��rL.a�R82��M��YPk�.���OF��.���e�{�CN���^�1�"M�^�a�С�Q`UPS��!$��M�QW�$�m�VGF�$R �MH��P2�� H�5� ΐq��ΐ�$([MH[�VP�uoY�����$)��D��hg��VPF��"MH�G̑`e!�+�V/vpcm�N��ՙ�N��$��VPRqd)��C	V�x�V� "�X�,��1�($TIa�t\muh��K��etpK��A%Y�VP%ɠ�!PyN���GeneB�rip����8��extt���Y�m�"�(��HB ���)��x��������Ȣ�res!.�yA�ɠn����*���p�@M�_�NĀ6L������yAvL�Xr��̈2��"R;�Ƚ\r�a��	P�� h86���Gu+ʸ�Ͽ�SaeLɨm�9�69�P��Ȩr�Ȩ2�ɹ1��n	2�h� �0L�XR}�RI{�e� L�x���Ac�Ș���N�vx�8L��"��2\r�]�N�82�d���b�� �a��y1��/�k�@���A��ruk�ʘ L��sop��H�}�ts{�����s��9��oj965��Sc��<h��5 J9�{��
�PL�J	een���t I[
x�co�m��Fh�L�4 J���fo��DI�F+�6�Q����ra#ti|��p��1�0�
R8l߾�M���Ȅ�P��8� �j�m�K�X�HZ����N$�oڠ��3�q��3vi���80�~�l Sl�yQ��tpk�xb�j�.�@� R�d������,/n(��8�8�0���
:�O08�<�Q}�CO���P]T��O (��.��Xp|�~H���?�v� �wv��8�2q2�pm���722��j7�^�@ƙ���3cf�=Yvr���vcu���O�O�O �O_#_5_7�3Y_��gwv4{_�_w�ʞ��ust_�_�cus�_�Z��oo,o�>oPo�io��nge���(pLy747�jWcelʨHM47ZK�Eq {���[m�M3FH�?�(wsK�8�J�n���o��fshl;��wmf�ڢ�? :�}(4	<gs J{��II)̏rމw��X�774k�L��/7ntˏ݊e+�f��se�/�aw��H8�ɐ��EX \�!+:� �p��~�00��n�h�,:Mo+�xO��1g "K�O��\a��#0��.8���{h�L?8�j+�mon�:�͙t�/�st�?-�w �:���)�;��(=h�;
d Pۻ�{:o  ��� �J�0��re�����STD�!tre?LANG���<81�\tqd���x����rch.�������htwv��WWָ� R7�9��"Lo�51 (�I�W�h�Ո�N4�aww� չvy �623c�h; a?�cti�֘!H�X�iؠ�t ��n,�։����yj��"AJP@�L3p�vr{�H�6�׽!��- SeT� �E3�) G�J934���LoW�4 (S������� <���911 ��8!4�j9�所�+���y�
��	�bt.N�ite{�R �� I@Ո�����P��������	 ����Z�vol��X ��9�<�I�pئ��ld*���F�8C64{��?��K��	�k扐�֘1�wmsk��M�q�Xa��e����p���0RBT�1ks.OPTN�q�f�U$ RTCamT��y��U��y@��U��UlU6L��T�1Tx����SF�q�Ue�6T��USwP W�b DT�qT2h�T�!/&+p��TX�U\j6&��U U�UsfdO&�&ȁT����662DPN��bi��%�Q�%62 V��$���%�� �#(��(6To6e St�%��#5y�$�)5(To�%tT0�%5��W6T���%�#�#orc��#I���#���%�cct�6ؑ?�4=\W6965"p6}"�#\j536���4�"�?kruO O,IAm?Np�C �?t�0<<O�;�e �%����?
;gcJ7 "AyV�?�;avsf�O0__&_8WtpD_V_"0GT�F|_:UcK6�_r�_r�O�3e\s�Or2^y`O:�migxG�vgW! m�%��!8�%T�$E A{6�p�o6��#37N�)5R!5_2E���$0���$Ada�Vd���V�?�;Tz7�_�e7DDTF9���#8�`�%���4y�ted `Z@�A}�@�}�04N�`}�}���}�dc& $}����u 6�v�8�v1�u1\b�u$2x}���}� R83�u�"}��"}�valg���Nrh�&�8��J�Y�o�ue��� j�70�v=1��MIG�uerfa��{q����E�N�ء��EY=E�ce A���� ���pV�e�A!���2Յ@�Q�%��u1�e�i�@���H�e����J0� �'��b��T��E In�B�  W�|���537g����(M%I�t�Ԇr��ݟ��am���nеv!4g�U -�v J߆8�`��F���P�y�ac��p�2���Rɏ jo�<�2�� djd�8r}� og\k�0���g��wmf�F;ro/� Eq'�4"�}�3 J8��oni[��ᅩ}Ĵ��� o� ��ʛ��m$@�R�e��{n�Д��V�o������  �����裆"�POS\����ͯ �menϖ�⑥OM�o�43��� �(Coc� An[�t����"e�a\�vp��.ރ�cflx$�le���8�hr�tr�NT�� CF+�x E�/�t	qi�M�ӓxc��p�f�lx����Zċcx��
0 h��h�8��mo��=� Hع��)� (�vSE�R,���g�0߆0\r�vX�= ��I �7 - �ti��Hv��VC�828��5��L"�RC��n# G/���w�P�y�;\v�vm "o�l�@��x`��=e�ߠ-�R-3?������vM [�AX/2�)�S��rxl�v#�0��hy8߷=� RAX춡A�����9�H�E�/Rצ����h߶"�RXk��F�˦8�5��2L/�xB8�85_�q�Ro�0i9A��5\rO�9� K��v����8����.�n "�v��88��8s�i ?�9 ���/�$�y O�MS�"���&�9R Hq74&�`�745��	p��p��ycr0�C�c�hP0� j�-`�a%?o��6D950R7�trl��ctl�O�APC���j�uqi"�L���  �����^棆!�A���qH��&-^7����� ��6196C�q�794h��Ƙ� M�ƔI��9�9��(��$�FEAT_ADD ?	���Q�%P  	 �H._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n���������TDEMO� fY   WM_�� ������// %/R/I/[/�//�/�/ �/�/�/�/�/?!?N? E?W?�?{?�?�?�?�? �?�?�?OOJOAOSO �OwO�O�O�O�O�O�O �O__F_=_O_|_s_ �_�_�_�_�_�_�_o oBo9oKoxooo�o�o �o�o�o�o�o> 5Gtk}��� �����:�1�C� p�g�y�������܏ӏ ���	�6�-�?�l�c� u�������؟ϟ��� �2�)�;�h�_�q��� ����ԯ˯ݯ���.� %�7�d�[�m������� пǿٿ���*�!�3� `�W�iϖύϟ����� ������&��/�\�S� eߒ߉ߛ��߿����� ��"��+�X�O�a�� ������������� �'�T�K�]������� ����������# PGY�}��� ���LC U�y����� �/	//H/?/Q/~/ u/�/�/�/�/�/�/? ??D?;?M?z?q?�? �?�?�?�?�?
OOO @O7OIOvOmOO�O�O �O�O�O_�O_<_3_ E_r_i_{_�_�_�_�_ �_o�_o8o/oAono eowo�o�o�o�o�o�o �o4+=jas �������� 0�'�9�f�]�o����� ����ɏ�����,�#� 5�b�Y�k��������� ş����(��1�^� U�g������������ ���$��-�Z�Q�c� �������������  ��)�V�M�_όσ� �ϯϹ��������� %�R�I�[߈�ߑ߫� ����������!�N� E�W��{������ �������J�A�S� ��w������������� F=O|s ������ B9Kxo�� ����/�/>/ 5/G/t/k/}/�/�/�/ �/�/?�/?:?1?C? p?g?y?�?�?�?�?�?  O�?	O6O-O?OlOcO uO�O�O�O�O�O�O�O _2_)_;_h___q_�_ �_�_�_�_�_�_o.o %o7odo[omo�o�o�o �o�o�o�o�o*!3 `Wi����� ���&��/�\�S� e������������ ��"��+�X�O�a�{� ���������ߟ�� �'�T�K�]�w����� �����ۯ���#� P�G�Y�s�}������� �׿����L�C� U�o�yϦϝϯ����� ���	��H�?�Q�k� uߢߙ߫�������� ��D�;�M�g�q�� ���������
��� @�7�I�c�m������� ��������<3 E_i����� ��8/A[ e������� �/4/+/=/W/a/�/ �/�/�/�/�/�/�/? 0?'?9?S?]?�?�?�? �?�?�?�?�?�?,O#O 5OOOYO�O}O�O�O�O �O�O�O�O(__1_K_ U_�_y_�_�_�_�_�_ �_�_$oo-oGoQo~o uo�o�o�o�o�o�o�o  )CMzq� �������� %�?�I�v�m����������ُ���;�  2�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������|'9  : >Ugy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ������������ �%�7�I�[�m���� ������������! 3EWi{��� ����/=C6Yk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ ASew���� ���+=O as������ �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/��A��$FEAT_�DEMOIN  �E��q��>��Y�INDEXf��u��Y�ILECO�MP g�����t�T����SETUP2 �h����� � N ܑ��_AP2BCK 1i��?  �)B��"�%�C�>���1� n�E����)���M�˯ �������<�N�ݯr� �����7�̿[��� ��&ϵ�J�ٿWπ�� ��3�����i��ύ�"� 4���X���|ߎ�߲� A���e�����0�� T�f��ߊ�����O� ��s�����>���b� ��o���'���K����� ����:L��p�� ��5�Y�}� $�H�l~� 1��g�� /2/ �V/�z/	/�/�/?/ �/c/�/
?�/.?�/R? d?�/�??�?�?M?�?�q?O�?O<O���P�� 2�*.cVRCO�O�0*�O��O�3�O�O�5w@PC��O_�0FR6:D�O=^�Oa_�KT�� �_�_&U�_�\h�R_�_�6*.FzOo�1	(SoEl�_io�[STM �b�o�^+P�o�m�0iPe�ndant Pa'nel�o�[H�o ��g�oYor�ZGIF|��e�Oa��ZJPG �*��e�0��z��JJS������0@���X�%
J�avaScriptُ�CSʏ1��f��ۏ %Cas�cading S�tyle She�ets]��0
AR�GNAME.DT���<�`\��^����Д៍�АDISP*ן���`$�d���V�e��CLLB�.ZI��=�/`:\Ҩ�\�����Co�llabo鯕�	?PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V�9������$�4i���V���z����!ߘ�TPEIN�S.XML(�@�:�\<����Cust�om Toolb�ar}��PASS�WORD���>F�RS:\��� %�Passwor�d Config ��?J���C��"O�� 3�����i����"�4� ��X���|�����A� ��e�����0��T f�����O� s��>�b� [�'�K��� /�:/L/�p/��/ #/5/�/Y/�/}/�/$? �/H?�/l?~??�?1? �?�?g?�?�? O�?�? VO�?zO	OsO�O?O�O cO�O
_�O._�OR_d_ �O�__�_;_M_�_q_ o�_�_<o�_`o�_�o �o%o�oIo�o�oo �o8�o�on�o�! ��W�{�"�� F��j�|����/�ď S�e���������T� �x������=�ҟa� �����,���P�ߟ� �����9����o�� ��(�:�ɯ^����� #���G�ܿk�}�ϡ� 6�ſ/�l�����ϴ� ��U���y�� ߯�D� ��h���	ߞ�-���Q����߇��,��$F�ILE_DGBCK 1i������ �( �)
SUMMARY.DG,���MD:`�����Diag S?ummary����
CONSLOG���y����$���C�onsole l�og%���	TPA'CCN��%g������TP Acc?ountinF����FR6:IPKDMP.ZIP�����
��)����Exception-�����MEMCHECCK�����8��Memory D�ata��LN{�)�RIPE�p��0�%�� Packet 9LE���$Sn�STAT*#�� %LSt�atus�i	F�TP�/�/��:�mment T�BD=/� >)�ETHERNE��/o�/�/��E�thernU<�figuraL��'!?DCSVRF1//�)/B?�0 ve�rify all�E?�M(5DIFF:? ?2?�?F\8diff�?}7o>0CHGD1�?�?�?LO �?sO~3&�
I2BO)O;O�O� bO�O�OGD�3�O�O�OT_ ��O{_
VUPDA�TES.�P�_���FRS:\�_�]���Updates� List�_��P�SRBWLD.C	Mo���Ro�_9��PS_ROBOW�EL^/�/:GIG���o>_�o�Gi�gE ��nost�icW�N�>��)�aHADOW��o�o�ob�Sh�adow Cha�nge��*8=+"rNOTI?=�O��Noti�fic�"��O�{A�PMIO�o���h��f/��o�^U�*�UI3�E�W�L�{�UI������ B���f��_������� O���������>�P� ߟt������9�ί]� 򯁯�(���L�ۯp� �����5�ʿܿk� � ��$�6�ſZ��~�� wϴ�C���g���ߝ� 2���V�h��ό�߰� ��Q���u�
���@� ��d��߈��)��M� ��������<�N��� r����%�����[��� �&��J��n� �3��i�� "�X�|� �A�e�/�0/ �T/f/��//�/=/��/�/�$�$FIL�E_�PPR�P���� �����(MDONL�Y 1i5�  
 �z/Q?�/u? �/�?�?t/�?^?�?O �?)O�?MO_O�?�OO �O�OHO�OlO_�O_ 7_�O[_�O_�_ _�_ D_�_�_z_o�_3oEo �_io�_�oo�o�oRo �ovo�oA�oe w�*��`�����&�O��*VI�SBCK,81;3�*.VDV�����FR:\o�ION?\DATA\��/���Visio�n VD filȅ��&�<�J�4� n������3�ȟW�� ����"���F�՟�|� �����m�֯e����� �0���T��x���� ��=�ҿa�s�ϗ�,� >���b���ϗϼ� K���o��ߥ�:����^����ϔ��*MR2_GRP 1j;��C4  B�}�	 71�������E�� E� � F@ F�5�U������L����M��Jk��Lzp�JP�ߣFg�f�?��  S����9�Y�9}�9���8j
�6���6�;��A��  ���BH��B-���B���$��������������@UUU#�����Y�D� }�h����������������
C��_CF�G k;T �M���]�NO� :
F0�� � \�RM_C�HKTYP  B0�}�000��{OM_MIN	�x���50X�� SSBdl5:0��bx�Y����%TP_DEOF_OW0x�9>�IRCOM���$GENOVR/D_DO*62��THR* d%d��_ENB� ^�RAVC��mK�� ��՚�/3ĩ/��/�/�� ��M!OUW s���}��ؾ��8�g�;?�/7?Y?[?o  C��0�����(7�?�<B�?B�����2��*9�N SM�TT#t[)��X�4��$HOSTCd1=ux���?��� MCx��;�zOx�  27.�0�@1�O  e �O�O	__-_;Z�O^_�p_�_�_�LN_HS	a�nonymous@�_�_�_oo1o yO��FhFk�O�_�o�O �o�o�o�oJ_'9 K]�o�_��� ��4o�XojoG�~ �o^�������ŏ� ����1�T���y� ����������,�>� @�-�t�Q�c�u����� ����ϯ���(�^� �M�_�q�����ܟ�  �ݿ��H�%�7�I� [Ϣ�ϑϣϵ���� l�2��!�3�E�Wߞ� ��¿Կ����
����� ��/�v�S�e�w�� ������������ +�r߄ߖ�s������ �����������'9 K]������� ��4�F�X�j�l> ��}����� �//1/T��y/��/�/�/�/.D\AEN�T 1v
; P�!J/?  � �/3?"?W??{?>?�? b?�?�?�?�?�?O�? AOOeO(O�OLO^O�O �O�O�O_�O+_�O _ a_$_�_H_�_l_�_�_ �_o�_'o�_Koooo 2o{oVo�o�o�o�o�o �o5�oY.��R�v��zQUICC0���3���t14��"����t2���`�r�ӏ!ROUTERԏ��#�!PCJOG$����!192.�168.0.10���sCAMPRT,t�P�!d�1m�����RT폟�����$NAME !�*?!ROBO����S_CFG 1u��) ��Auto-sta�rtedFTP&��=?/֯s ����0�B��f�x� ��������S����� �,���������ϼ� ޯ���������ʿ'� 9�K�]�oߒ�ߥ߷� ��������(: ~�k�Ϗ������� ������1�C�f��� y������������,� >�R�?��cu� �`�����( �$M_q���� �� /H%/7/ I/[/m/4�/�/�/�/ �/�~/?!?3?E?W? i?����?�/�?/ �?OO/O�/�?eOwO �O�O�?�ORO�O�O_ _+_r?�?�?�?�O|_ �?�_�_�_�_o�O'o 9oKo]ooo�_o�o�o �o�o�o�oF_X_j_ ~ok�_����� �o���1�TU���y���������U�)�_?ERR w3�я��PDUSIZ � g�^�p����>�WRD ?�r�Cq�  ?guestb�Q��c�u�������"�SC�DMNGRP 2�xr�����Cqg�\�b�K� �	P01.00� 8(q   e�5p�5pz�5p�B  �{ ����H����L��L��L�����O8�����l������a4� x��Ȥ�Zx��8���\����)�`�;�������d�.�@�R��ɛ_GROUېy*�����	ӑ����QUPD  d?u����İTYg�����TTP_AUTH 1z��� <!iPeOndan��-�l����!KARE�L:*-�6�H�K�C]�m��U�VI�SION SET ���ϴ�g�G�U����� �R�0��H�Bߏ�f��x��ߜ߮���CTRL {����g��
S�FFF9�E3��AtFRS�:DEFAULT�;�FANUC� Web Server;�)����9� K��ܭ����������߄WR_CONF�IG |ߛ �;��IDL_C_PU_PCZ�g�sB�Dpy� BH_��MINj�)�}�GNR_IO��g����a�NPT_SIM�_D_�����STAL_SCRN��� ���TPMOD�NTOL������R�TY��y���� �E�NO���Ѳ]�OL_NK 1}��M� �������eMASTE��ɾe�SLAVE ~���c�O_CFGٱBUO�O@CYCLEn>T�_ASG 1ߗ+�
 ���� //+/=/O/a/s/�/��/�/�/��NUM���
@IPC�H�^RTRY_CNZ���@�������� @kI��+E�z?E�a�P�_MEMBERSg 2�ߙ� $���2���ݰ7�?�9�a�SDT_ISO�LC  ����$J23_DSM�+�3JOBPRsOCN��JOG���1�+�d8�?��+�O�/?
�LQ�O__�/_�OS_e_w_�_`��O Hm@��E#?&BP�OSREQO��KANJI_���a~[�MON ����b�yN_goyo�o�o��o�Y�`3�<� �0�e�_ִ��_L���"�?`EYLOGG+INLE��������$LANGU�AGE ��<eT� {q�LGa2Y�	�b���g�xP���  ��Rg�'��b���>��MC:\RSC�H\00\<�XpN�_DISP ��+G�J��O�O߃LO�Cp�Dz���A�sOGBOOK ������󑧱����X�����ϏᏀ���a�*��	p�����!�m��!����=p_BUFF [1�p��2F�๟���՟D� C�ollaborativǖ���F�=� O�a�s�������֯ͯ ߯���B�9�K����DCS �z� =���'�f��?ɿ�ۿ���H@{�IO ;1�� ~?9����9�I�[�mρϑ� �ϵ����������!� 3�E�Y�i�{ߍߡ߱���������E��TMNd�_B�T�f�x�� ������������� ,�>�P�b�t��������L��SEVD0�.�TYPN1�0$6���QRS"0&|��<2FL 1�"�J0�������0�GTP:pO�F�NGNAMp1D�mr�tUPS��GI"5�aO5�_�LOADN@G �%�%TI�pZ�UZAUN#�(MAXUALRM�'p���(��_PR"4�F0d��1�B_P{NP� V 2�C�	MDR07�71ߕ�BL"8�063%�@ ��_#?�ߒ|/�C�A�z�6��/���/Po@�P 2��+ ��ɖ	T 	t  ��/�%W?B? {?�k?�?g?�?�?�? O�?*OONO`OCO�O oO�O�O�O�O�O_�O &_8__\_G_�_�_u_ �_�_�_�_�_o�_4o oXojoMo�oyo�o�o �o�o�o�o0B% fQ�u���� ����>�)�b�M� ����{��������Տ ��:�%�^�p�S��������D_LDX�DISApB�M�EMO_APjE� ?C
  �,�(�:�L�^�p�������� 1�C ����4�����૟4��X���C_M?STR ���w��SCD 1��� L�ƿH��տ���2� �/�h�Sό�wϰϛ� �Ͽ���
���.��R� =�v�aߚ߅ߗ��߻� ������<�'�L�r� ]���������� ����8�#�\�G���k� ��������������" F1jUg�� �����B -fQ�u����h�MKCFG 񓆽�/�#LTAR�M_��7"�0�0N/V$� MEgTPUᐒ3�����ND� ADCOLxp%� {.CMNT�/s �%� �����.E#>!�/4�%PO�SCF�'�.PR�PM�/9ST� 1���� 4@��<#�
1�5�?�7 {?�?�?�?�?�?�?)O OO_OAOSO�OwO�O��O�O�O_�A�!SI�NG_CHK  ��/$MODAQ�,#����.;UDE�V 	��	M�C:o\HSIZE�ᝢ��;UTASK� %��%$12�3456789 ��_�U9WTRIG +1���l3%%��9o���"ocoFo5#�VYP�QNe��:SEM_�INF 1�3'� `)�AT&FV0E0�po�m)�aE0V�1&A3&B1&�D2&S0&C1�S0=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o '��K������ ��я:�L�3�p�#� 5���Y�k�}������ $�[�H���~�9��� ��Ưد��������ӟ �V�	�z�������c� Կ����
��.��� d��)�;��Ͼ�q��� ����˿<���`�G� �ߖ�IϺ�m�ϑϣ� ���8�J��n�!ߒ��M�������h_NIwTOR� G ?�[�   	EX�EC1�/�25�3�5�45�55��P7�7*5�85�9�0�� ��4��@��L��X� ��d��p��|�������2��2��2���2��2��2��2���2��223ʡ�3��3@�;QR_�GRP_SV 1ݚ�k (�5W�r3��������MO�Q_�D��^�PL_N�AME !3%�,�!Defa�ult Pers�onality �(from FD�) �RR2� �1�L6(L�?�,0	l d �������� //(/:/L/^/p/�/��/�/�/�/�/�/ZX2 u?0?B?T?f?x?�?�?�?�?\R<?�?�? O O2ODOVOhOzO�O��O�OZZ`\RD�?�N
�O_\TP�O :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo _)_~o�o�o�o�o�o �o�o 2DVh z�[omo���� 
��.�@�R�d�v����������Џ� �Ef  Fb� gF7�����!��d�?�Q�6� t���������ʜ8����� ݘ� ���"�@�F�d���� �"𩯹�� A� � ϩU[�$n��B�E ��� � @D��  �?�� �?x�@��A@�;f�|�FH� ;�	l,��	 |��j��s�d�>��� ���� K(��Kd�$2K ��J7�w�KYJ���ϜJ�	�ܿ��� @I���_f��@�z��f��γ�N�������	Xl�������S�Ľ�Ô��X������5���  �����A?oi#��;���� � �l� �Ϫ�-���ܛ�G�G����@�n�@a   �  ��ܟ*��͵	'� � �H�I� � � �Рn�:����l�È=������@�ߚЕ����/�����̷yNP�  ',����-�@
�@����?=�@A�~��B�  Cj�a�Be�Ci��@#��Bи�T J� ,ee��^^ȹBР��P�����̠�����ADz ՟�n�3��C�i�@��R�R�Yщ��  ��@� ���  =��?�ff������n� ɠ#�@y9G
(���I�(�@uP~����t�t����>����;�Cd;���.<߈<��g�<F+<AL�������,�d�|,�̠?fff?���?&&��@���@x��@�N��@���@T� H�ِ�!-�ȹ�| ��
`������ �//</'/`/r/]/�/��eF���/�/ �/�/m?��/J?�(�E��G�#�� FY�T?�?P?�?�? �?�?�?O�?/OO?O eO�ħO�IQOG�? �O1?�OmO_0_B_T_"������A_�_@	_�_�_�_ o��A��aAn0 bФ/o C�_pUo�_�Op��؃o��o�o�o���W������oC�E�  q�H�d��؜a@q���e�F�BµWB�]�NB2�(A���@�u\?��D�������b��0�|�uR�Ｃ�
x~������Bu*�C��$�)`��$ ���GC�#���rA�U����1��eG�D�I�m�H�� I:��I�6[F����C�I��J��:\IT�H
~QF�y���p�*J�/ �I8Y�I��KFjʻCe�o�� s�����Џ���ߏ� *��N�9�r�]����� �������۟���8� #�\�G�����}����� گů���"���X� C�|�g�����Ŀ��� ����	�B�-�f�Q� ��uχ��ϫ������ ��,��P�b�M߆�q� �ߕ��߹�������(� �L�7�p�[����������s(la��33:����$�le�3���d�,�4���@�R�wa����l�~�wa���ex����wa4 �{�� ����(L:ue%P�P~�A�O�������	����G2W} h������/����O�O7/m/[(d =�s/U/�/�/�/�/�/ ?�/1??U?C?y?�=  2 Ef9g�Fb��77�9fBX)aa)`C9A`�&`w`@-o�?9de�O-OOQOpn�?�?�O�O��O�O9c?�0�A7hJldw`w`!w`xn
 �O9_K_ ]_o_�_�_�_�_�_�_��_�_o#ozzQ ���h��G���$�MR_CABLE� 2�h ��a�T� @@��0�Ae��a�a�a���`��0�`C�`�aO8�tB����a�=��"R�`E5����F�o�f�#���0��0�DO�5��`�,��M�qQ D������o�ho8  ���C�0]7�d4�`�����&z��bEM3�q"4��`y`�By`C�p�bHE���`�br�ڰ�5Dg�9Hv��Ҡ`��0�q�p�b0�z�`���	��T D�g+�y/o�c -���H� �2���V��� ��������'�"��� D���^q��o��\ ��������������w*,�** \c�OM �ii����ŋ��P%�% 234567O8901i�{� f�H����������1�����
��`��not sent� 5���;��TESTFECS�ALGR  eg�`��1d.�š�a�`� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.x�ml��ֿkqY��DEFAULT�-�i4\bGRP 2�M�  �E�7�E�  �%For�ce�sor c?heck  ���b��z��p����h5-���ϻ��������%�!1st cle�aning of� cont. v��ilation��}�Rߗ+��[��Дߦ߸���me;ch�cal`������0��h5k�@�R�d�v����>(�rolle_Ƶ����/���(��:�L��Basi�c quarte�rly�������,�������������M��:(�"GpP(�X_h5�������#C���M"��{Pbt�|��Suppq�?grease���?/&/8/J/�\/��C+ ge��./ batn�y`/��/h5	/�/�/�/?� ?_�ѷen'�v��/�/��/��?�?0�?�?�?�G=?O�qp"CrB1O��0 �/`OrO�O�O�O�t$,��Lf��C-(��A�O:�OO$_6_H_Z_�l_�t*cabl,�O(���S<(��Q�_:�
_�_�_oo�0oo)(Ӂ/�_�_����_�o�o�o�o�o��O@hau1�l�2r x(�<qC:��op������_ReplaW�fU��2�:�._4�F�X�j�|�(�$%���ߟ ����#���
��.�@� ��d���ŏ׏����П ����U�*�y����� r���������	�q�� ?�߯c�8�J�\�n��� ϯ�����ڿ)���� "�4�Fϕ�jϹ�˿�� ����������[�0� ϑ�fߵϊߜ߮��� ��!���E�W�,�{�P� b�t����߼��� ��A��(�:�L�^��� ������������  $s�H������q �����9] o�Vhz��� U�#�G/./@/ R/d/��/�/��// �/�/??*?y/N?�/ �/�?�/�?�?�?�?�? ??Oc?u?JO�?nO�O��O�O�O+Jkb	 H �O�O__6M2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o�*<ND@ ̾bA?�  @!Q _���Fwp�� �H* �** @A>F�pRT��f�x�:�������ҏ��eO^C7�Տ#�5� G�	�k�}���ُ��� c�����W��C�U� g���ß)�����ӯ� ��	��-�w�����9� ������m�Ͽ��=��O�E!Q�$MR�_HIST 2��>EN�� 
 \�
B$ 2345678901^�f�#�
�]�9O���φ� ��O�)�;����q� �ߕ�L�^߬����ߦ� ���7�I� �m�$�� ��Z���~������!� ��E�W��{�2������h�����:�SKCF�MAP  >EKQ��r5�!P�����ONREL7  .�3����EXCFENB�8
��QFNC�XJJOGOVL�IM8dNá ��K�EY8��_�PAN7����R�UN����SFSPDTYPx<C��SIGN8J�T1MOT�G���_CE_GRP7 1�>EV� �@�����/Ⱥ ��/�/U//y/ 0/n/�/f/�/�/�/	? �/???�/c??\?�? P?�?�?�?�?�?O)O�OMO,���QZ_E�DIT5 )TC�OM_CFG 1����[�O�O�O }
�ASI �yB3�
__+[_�O_��>O�_bHT__ARC_U.���	T_MN_MO�DE5�	UA�P_CPL�_gN�OCHECK ?��� ��  o.o@oRodovo�o�o �o�o�o�o�o*�!NO_WAITc_L4~GiNT�A����EUwT_E�RRs2���3��@ƱJ�����>_�)��|MO�s��}x�:Ov���8�?������ l��rP�ARAM�r�����j���5�5�G� = ��d�v�~� X������������֟0�0����b�t������SUM_RSPACE�����Aѯ�ۤ�$ODRDS�P�S7cOFFS?ET_CARt@�_��DIS��PE?N_FILE:�7��AF�PTION�_IO��q�M_�PRG %��%�$*����M�WOR�K �yf ���춍��� N  "�������	 �������It��RG_D?SBL  ��C��{u��RIEN�TTO7 �C�� A �UT__SIM_Dy����V�LCT ���}{B �٭��_�PEX�P=��RA-T�W dc���UP ���`����e�w�]ߛߩ���$�2r�L6�(L?���	l d������&� 8�J�\�n����� ���������"�4�F�X���2�߈��������������*�< w�Tfx��������J`[ˣG���Tz��Pg����� �/"/4/F/X/j/|/ �/�/�/���/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?�/�/,O >OPObOtO�O�O�O�O �O�O�O__(_:_��O��y_�]2ӆ��_�^�_�_�W^]^] ��/ooSog��Hg rohozo�o�o�o�o�o�F`�#|`�A��  9y����OK�1��+k�+�����<�E�A�nq @D��  �q����nq?���C��s�q1� �;�	l��	 �|�Q�s�r�q�>��u �sF`H�<zH~�H�3k7GL�zHpG�99l`7�k_B�T�F`C4��*k�H���t��-�Ae����k������s���  ���������EeBVT����dZ=�3��ڏ ��@�q-�Fk�y�{FbU��= n@6�/  ���z�Fo���Be	'� �� ��I� ��  �:p܋=����ڟ웆�@����B�,���B�Ȇ�g�AgN����  a'|���g��B��p�BӀC׏����~@  #�Bu��&�ee�^^މB:p2���>�`m�6p�Z�=Dz?o }�܏������׿�������Ǒ��� f�  O� �M���*�?�ff�_8�J�ܿC 3pϑ�ñ8=  �ϵʖq.·�(= �ŁP���'��s�tL�>���/�;�Cd;���.<߈<��g�<F+<L  ��^oiΚrd@��r�6p?fff?�?�&�п�@��@�x��@�N�@���@T싶� Z���ћtމ�u�߈w 	�x��ti�>�)�b�M� ��q���������� ���:�%�^��������W���S�E�  G��=F�� F k���������1U @yd����� �q��	��{�A���h�����a��ird��A{/w/PJ/5/n/	�A��A���":t�/ C^/�/Z/< ލ?���/�/X1??���W����:g��pE� ~1�?�04�0
1�1@I�Ӏ��BµWB�]�NB2�(A���@�u\?����������b��0�|�uR�Ｃ�
�>������Bu*�C��$�)`���? ���GC�#���rA�U����1��eG���I�m�H�� I:��I�6[F����C4OI��J��:\IT�H
~QF�y�O�l@�*J�/ �I8Y�I��KFjʻC��-?�O �O__>_)_b_M_�_ �_�_�_�_�_�_o�_ (oo%o^oIo�omo�o �o�o�o�o �o$ H3lW�{�� �����2��V� h�S���w�����ԏ�� �����.��R�=�v� a�������П����ߟ ��<�'�`�K�]��� ������ޯɯ��&��8�#�\��3(J���33:a������J��3��c4�����������������ڿ�n����ex��n�4 �{2� 2�r�`ϖτϺϨ��%%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ����� �����3��W�B�{�f�4���������d �A����!��1�3�E� {�i�������������  2 Ef�7�Fb�7��6BX�!�!� C9� �� n�@�/`r������#x���+=�3?, V�8Jv�n�n��n��.
 D�� ���//%/7/I/�[/m//�/�:� ���ֻ�G���$�PARAM_ME�NU ?2���  �DEFPULS�E�+	WAIT�TMOUT�+R�CV? SH�ELL_WRK.�$CUR_STY�L� 4<OPT�JJ?PTB_?Y2C�/?R_DECSN  0�Ű<�?�?�?�?�? OO?O:OLO^O�O�O�O�O�O�!SSREL_ID  .�����EUSE_P�ROG %�*%8�O0_�CCCR0�B���#CW_HOST7 !�*!HT�_�=ZT��O_�Sh_zQ��S�_<[_TIME�
2�FXU� GDE�BUG�@�+�CGI�NP_FLMSK�o5iTRDo5gPG�Ab` %l�tkCyHCo4hTYPE�,� �O�O�o# 0Bkfx��� ������C�>� P�b���������ӏΏ �����(�:�c�^��p�����7eWORD� ?	�+
 	�RSc`n�PNeS��C4�JOv1΃�TE�P�CCOL�է�2��gLP� 3��n��OjT�RACECTL �1�2��! ���> ?�Қ�q�DT Q��2�Ǡ��D �o :����3Ԡ�Ԡ�@�}�ׯ���;�4��4��4��� ;�u:�q:�8����;�	8�
8�8�*8�8�8�8��@*:�8�8���P� ���ٱ޴���ؿ�$�6���
ϸl�~�(� *8�+ +��(��)���� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������'
 ,�>�P�b�t������� ��F�X�С�*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6@ub t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀�V �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�?��1�$PGTRA�CELEN  ��1  ����0��6_UP ����A�@�1����1_�CFG �E��3�1
@�<D�0<DZO<C�0uO$B�DEFSPD e�/L�1�0��0�H_CONFIG� �E�3 ��0�0d�D��2 	�1�APpDsA�A�0ۂ�0IN'@TROL �/MOA8pE�QPE�E��G��A<D�AILI�D(C�/M	bTGR�P 1ýI �l�1B  ������1A�33�FC� F8� _E�� @eN	�A��AsA�Y�Y�A�@�� 	RO�Hg�_ ��8cokB;`baBo�,o>oxobo�o�1>�?��?B/�o�o�~�o =%<��
C@y d��"����<��  Dz@�I� @A0�q� �������ˏ ���ڏ���7�"�4�@m�X���|���Ú)ґ�
V7.10b�eta1HF �@����Aq���Q  �?M� �BܠP�p ��C��&�B�EQA���Q�P�Q��� ß[�m����<CA ��0�b�@���f����'��ҡ�R�ܣ�R�љ���1�i�=�����t<B!C�eQKNOW_M � lE7FbTSV ĽJ�BoC_� b�t�����������࿨�1�]aSM�SŽK� ���	NB�0���ĿK���-�bb��A�R P����0�Ŗ��VbQMR�S��T�i�N���d���V]STކQ1 1�K
 �4MU�iǨj�  K�]�oߠߓߥ߷��� ����2��#�h�G�Y� ��}�������
���(���,�27�I��1G�<t�H��P3^�p�����,�4��������,�5(:,�A6Wi{�,�7����,�8�!�3,�MAD�6 �F,�OVLD  �KD�xO.�PARNUM  ��MC/%�SCH� �E
9'!G)�3Y%U�PD/��E�/P�_CMP_��0@�0�'7E�$ER_CHK�%5H�&�/�+�RS���bQ_MOȤ+?=5_'?O�_R/ES_G6��:�I� o�?�?�?�?O�?O 7O*O[ONOOrO�O�O�{4]��<�?�Oz5 ���O__|3 #_B_ G_|3V b_�_�_|3�  �_�_�_|3� �_�_o�|3Oo>oCo|2V �1�:�k1!�@c�?�=2THR_ICNRc0i!}�o5d�foMASS�o Z�g�MN�o�cMON_�QUEUE �P:�"�j0��O�N� �U1Nv�+DpENqDFqd?`yEXEo�`u� BEnpPAsO�PTIOMwm;DpP�ROGRAM %$z%Cp}o(/Br?TASK_I��~OCFG �$x��K�DATA�M�T���j12/ ď֏������+�=� O�a����������͟^��INFO�͘��3t��!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w�����Θ� '��FJ�6a K_N��T��˶ENBg ڽw1��i2��GN�2�ڻ� P(O�=����]ϸ�@�<��v� �u�u���dƷ_EDIT ��T�����G�WE�RFL�x�c)�RG�ADJ Ҷ�A�  $�?j00��a��Dqձӆ5O�?��ʨ�<u�)%e������FӨ��2�R��	H;plR�G�b_�>�pAodw�t$�*�=/� **:�j0�$�@�5Y�T���^��q�߈b~�L�� \�n��������� ������4�F�t�j� |�������������b LBT�x� ���:��$ ,�Pb���/ ����/~/(/:/ h/^/p/�/�/�/�/�/ �/V? ??@?6?H?�? l?~?�?�?�?.O�?�? OO O�ODOVO�OzO �O_�O�O�O�O�Or_ _._\_R_d_�_�_�_�_�_�_�f	g�io�p Wo�o{d�o�~o�o�zoB�PREF� �Rږp�p
~�IORITY�w�[���MPDSP�q��pwUT6�����ODUCT3������OG��_�TG��8��ʯrTO�ENT 1׶�� (!AF_I�NE�p,�7�!�tcp7�_�!�udN���!iccmv��ޯrXYK��ض���q)� 0,�����p��&� 	��R�9�v�]�o��� ��П������*��$N�`�*�sK��9}�߸����Ư ,�/�6쒯�����خ�A~t�,  �Hp ��P�b�t����u�w��HANCE �R��:�wd��连��2s�9Ks��PO�RT_NUM�s�p���_CARTREP{p�Ω��SKSTA�w nd�LGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_�a_seiban �o\��olߒ�}߶ߡ� ��������"���X� C�|�g�������� �����	�B�-�f�Q� ��u����������� ��,<bM�q �������(�L�VERSI�yp�w} disabledWSAVE ߾z�	2600H7K68S?�!ؿ0����/ 	5(�r$)og+^/y�e{/�/�/�/�/�*�,/?� �p���_�p 1��Ћ� �����Wh?z?�W*p/URGE��B�p}vlgu,�WF�0DO�v�Ʋ�vW%��4(�C�W�RUP_DELA�Y �\κ5R_?HOT %Nf�q�׿GO�5R_NORMAL&H�r6O�OZGSEMIjO�O�O(q_QSKIPF3��W3x=_98_J_\_ ]�_�_{_�_�_�_�_ �_�_	o/oAoSoowo eo�o�o�o�o�o�o�o +=aOq� �������'� �7�]�K�������)Eo�$RA{���K�/�zĀÁ_PAR�AM�A3��K �@.�@`�61�2�C<��y��C��6$�BÀBTI�F�4`�RCVTMkOUu�c��À�DCRF3��I ��+QBG���D�}�D	�N��1@�3�8<���]�YE2ޅ�����*��2S�_��k_ �;�Cd;��.�<߈<�g��<F+<L�� �Ѱ��d�u�L��� ����ϯ����)��;�M�_���RDIO�_TYPE  �M=U�k�EFPOS�1 1�\�
 x4/�����+�$/ <��$υ�pϩ�D��� h��ό��'������ o�
ߓ�.ߤ�Rߌ��� ����5���Y���i� ��*�<�v���r���� �����U�@�y���� 8���\������������?��c����2 1�KԿX�Tx�x��3 1�����nY�S4 1�'9K��/�'/�S5 1���/�/�/�/>:/S6 1�Q/c/�u/�/-??Q?�/S7 1��/�/
?D?�?��?�?d?S8 1� {?�?�?�?WOBO{O�?�SMASK 1����L��O�D�GXNO����F&�^��MOT�EZ�Ż��Q_ǁ��%]pA݂��PL_�RANG!Q]�_QO�WER �ŵ��P1VSM_DRY�PRG %ź%�"O�_�UTART ��^�ZUME_�PRO�_�_4o��_�EXEC_ENB�  J�e�GSP�D`O`WhՅjbTD�Bro�jRM�o�hI�NGVERSIOoN Ź#o��)I_AIRPU�RhP �O(�MMKT_�@T�P#_À�OBOT_ISO�LC�NTV@A'q^huNAME�l��o��JOB_ORD_�NUM ?�X�#qH768w  j1Zc@�r�
�rV�s��r�?�r�?�r�pÀPC_OTIMEu�a�xÀoS232>R1��� LTEA�CH PENDA1Nw�:GX�!O� Mainte�nance CoKnsj2����"���No Use B�׏������1�C�y�V�NPO�P@�YQ��cS�CH�_L`�%^ �	�ő��!UD1�:럒�R�@VAI�L�q@�Ӏ�J�QS�PACE1 2�ż ��YRs�i��@Ct�YRԀ'{��8�?��˯� ���"���7�2�c�u� ����G���߯ѿ򿵿 �(��u�AC�c�u� ����Ͻ�߿���ϵ� �(��=�_�qσϕ� C߹������߱��$� �9�[�m�ߑߣ�Q� �����߭��� ���	� W�i�{���M����� ��5���.S�e� w�����I������ �*?as� �E�����/ &//;/]o��� ���/2/�/?"?�/ 7?Y/k/}/�/�/O?�/ �/�?�?�?O0OOK�A��*SYPpM�*�8.3026�1 yB5/21/�2018 A ��WPfG|�H�_T�X`� !$CO�MME�$�USAp $ENABLEDԀ�$INN`QpIO�R�B�@RY�E_SOIGN_�`�AP�AsIT�C�BWRK�B=D<�_TYP�CRINDXS�@W�@�%VFRI{�_GR�PԀ$UFRAyM�rSRTOOL\V�MYHOL�A$�LENGTH_V{TEBTIRST�T�  $SEC�LP�XUFINV_�POS�@$M�ARGI�A$WgAIT�`�ZX2�\��VG2�GG1�AI �@�S�Q	g�`_WR�B�NO_USE_DyI�BuQ_REQ�B�C�C]S$CUR�_TCQP�R"a^f ��GP_STAT�US�A @ `�A3`�BLk�H$zcy1�h�P ��@}_�FX �@�E_MLT_CTf�CH_�J�`CO�@�OL�E�CGQQ$�W�@w�b#tDE�ADLOCKuD�ELAY_CNT��a3qGt�a$wf _2 R1[�1$X<�2[2�{3[3$Zwy�q%Y�y�q`%V�@�c�@�b$V�`�RV�UV3oh>b�@ � �d�0ar'MSKJ�LgWaZ��C`NRK�PS_RATE�0$���S
`�Q�TAC��PRDH���e�S*��a4�At�0�DG�A 0�P��flp bquS2�ppI�#`
`�P �
�S\`  }�A�R_ENBQ� �$RUN?NER_AXI�<`�ALPL�Q�RU�TH�ICQ$FLI�P7��DTFERE�N��R�IF_CH�SU�IW��%V)�G!1����$PřA�Q�P�ݖ_JF�PR�_P�	�RV_D�ATA�A  {$�ETIM����$VALU$��	�OP_  � �A  2� �SC*��	� �$ITPa_!�SQ]PNPOU}��o�TOTL�o�DS}P��JOGLIb�N�PE_PKpc�Of�ji��PX]PTAS��$KEPT_M#IR��¤"`M�b�APq�aE�@�y�`q�g@١c�q�PG��BRK6�x���L�I��  ?�SJ�q��P�ADEz�ܠBS{OCz�MOTNv�DUMMY16Ӂ�$SV�`DE_�OP��SFSPDO_OVR
���@�LD����OR��T-P8�LE��F����6��OV��SF��F����bF�d�ƣ&c)��fQc�LCHDLY>��RECOV���`���W�PM��gŢ�R�O������_F�?�� @v�S �NVE�R�@�`OFS�PC,�CSWDٱc�ձ��X�B����TRG�š��`E_FDO��MOB_CM}���B���BLQ�¢	�Q�̄V�za�BUP�g��G
��AM���@`K�̊�e�_M!�d�AMxf�Q��T$CA����DF���HBKXd�v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�3�A��ATIO�0��͠��US����WaAB��R+c�`tá`xDؾA��_AUXw�?SUBCPUP���S�`����3Եжc���3�FLA�B�HW_Cwp"�Ns&�]s�Aa��$UNI�TS�M�F�ATT�RIz�Z�CYC=L�CNECA����FLTR_2_F�I��TARTUP`Jp����A��LP�������_SCT*cF�_F�F_P���b�FqS��+�K�CHA/Q���*�d�RSD���Q����Q���_T�H�PROr���հE#MPJ���G�T�� �Q�DI��@y�RAILAC4/�bMX�LOf�xS��ځ���拁���+PR#�S`app��C� 	��F�UNC���RIN�`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ng�DAQ�B�rkL�D�र&q�M�K���TI���j���$�@RIA_S�W��AF��Pñ�#��%%�p9r1��MsOIQ���DF_~P�(�PD"LM-�F�A�PHRDY�DORG�H; _QP�>s%MULSE~Pz�T��*�� J��Jײ���FAN_AL�MLVG��!WRN�%HARDP��Uc�O�� K2$SHADOW]�kp�a02���� STOf�+�_,^�w�AU{`R��eP_SBR�z5����:F�� �3MPINF?�\�4��3gREGV/1DG�b+cVm �C�CFL(��?�DAiP��ҌZ`�� �����Z�	� �P(Q$�A�$Z�Q V�@�[�
o� ��EG��o���kAAR���㌵�2�axG��AXEROB��RED���W�QD�_�Mh�S�YA��AF��FS�GW�RI�P~F&�STRP����E�˰EH�)�$�D�a\2kPB6P��t=V��Dv�OTO�19)���ARYL�tR0�v�3���FI&�ͣ?$LINKb!\�J�Q�_3S���E���QXYZ2�Z5N�VOFF���R�RJ�XxPB��d0s�G�cFI�03g��������_J ��'�ɲ�S&qR0LTV[6���aTBja�"�b�C���DU�F7.�TUR� X��eĂQ�2XP�ЊgFL��E���x@�`�U9Z8����� 1	)�K��Mw��F9��劂����ORQj��G;W3���#�Ґd ���uz����1�tOVE�q_�M��ё?C�uEC �uKB�v'0�x-�wH� �t���& `��qڠ �B�ё�u�q�wh�EC�h����ER��K	B�EP����AT�K�6e9e�W����AXs�'��v�/� �R ����!�� � �P��`��`�3p�Yp�1�p�� ��  �� (�� 8�� H��  X�� h�� x�� ����ޙ�DEBU�$�%3�I��·RAB����ٱ�sV��� 
d�J、��@� ��������Q���a�� �a��3q��Yq+$�`%"\<�cLAB0b�u�'�GRO���b<��B_s��"Tҳ *`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθ0uݸ��PNT0��?�SERVE �Z@� $`EAV�!�PO����nP�!�P@�$!Y@ � $>�TRQ"�b
=��BG�K�%"�2\��� _ � l��5�D6ER)RVb(�I��V0`;�N��TOQ:�7�L�@P
�R��e G�%�Q��� <�50F� ,h�`�z�>�RA�? 2 d!�����S�  M��p0xU ����OCuG��  ��CO�UNT6Q��FZN�_CFGF� 4#��6��TG4�_�=�����(���VC ���M �"��$06��q ��FA E� &��X�@������$�A����AP��P@�HEL�0��� 5b`B_BA�S��RSR�6"�CSH����1�Ǌ�U2��3��4��5��6��7��8��}�R�OO����P�PNL�EA�cAB)ë ��A[CKu�INO�T���(B$UR0� =�_cPU��!0��OU+�Pd�8j��� V���TPFWD_KA1R��� ��RE(ĉ qP�P�>QUE�:�RO�p�`r0P1I � x�j�P�f��6�Q�SEM��0��� An��STYL�SO j�DIX�&������S!_TMCMANsRQ��PENDIt�$KEYSWI�TCH���kH}E�`BEATM83PE{@LE��>]�J�U��F��Sp�DO_HOM# Ol�@�EF�pPRaPB�A#PY�C� O�!<���OV_M|b<0 IOCM�dFQ��h�HKYA# D�Q�7��UF2���M���p�cFOR�C�3WAR�"�O}M|@  @S�T#o0U)SP�@1�2&3&4E���TЕO��L���8U�NLOv�D4K$E}DU1  �SY��HDDNF� ~M�BLOB  p��SNPX_AS�� 0@�0�о81$SIZ�1�$VA{���MUL�TIP-��# A�� � $ ��� /4`�BS��0�yC���&FRIFB�O�S���3� NF�ODBUP߰�%�@3;9(��ҋ�Z@ mx��SI��TEs\�r�cSGL�1T�R�p&�Н3B��@�0S'TMTq�3Pg@V�BW�p�4SHOWܾ5@�SV��_Gv�� 3p$PCJ�XPИ���FB�PH�SP AW�EP@V�D�0WC� ���A00��PB XG@ XG XG$ XG5VIU6VI7VI8VI9VIAVIBVI�XG�YF��0XGFVH��XbI1�oI1|I1�I1�I1��I1�I1�I1�I1��I1�I1�I1�I1�Y1Y2UI2bI2*oI2|I2�I2�I�`��X�I2p�X�I2�I2��I2�I2�I2Y2PY�p�hbI3oI3|IU3�I3�I3�I3�IU3�I3�I3�I3�IU3�I3�I3Y3YU4�i4bI4oI4|IU4�I4�I4�I4�IU4�I4�I4�I4�IU4�I4�I4Y4YU5�i5bI5oI5|IU5�I5�I5�I5�IU5�I5�I5�I5�IU5�I5�I5Y5YU6�i6bI6oI6|IU6�I6�I6�I6�IU6�I6�I6�I6�IU6�I6�I6Y6YU7�i7bI7oI7|IU7�I7�I7�I7�IU7�I7�I7�I7�IU7�I7�I7Y7TրVP� UD��y"ՠ��
<A62��t�R��CMD� ��M5�Rv�]��Q_h�R���e�����<�YSL���  � �%\2��+4��'��W�BVA�LU��b��'���F�H�ID_L���H�I��I���LE_���㴦�$0C�S�AC�! h ��VE_BLCK���1%�D_CPU5ɧ 5ɛ ������C�� ��R " � PWj��#06��LA�1SBћ������RUN_FLG�Ś����ĳ ����������H���ХĽ�TBC2��#/ � @ B��e ��S�8=�FTD	C����V���3dՆQ�THF�����R��L�ESERVE9��F��3�2�E�|�Н�X -$��LEN9��F��f�cRA��W"G�W_5��b�1��д2�MO$-�T%S60U�Ik�0�`ܱF����[�DEk�21LACEi0�CqCS#0�� _MA� pj��z��TCV����z�T�������.B i�'A�z�'AJh�#E�M5���J��@@i�V�z���2Q �0&@�o�h��JK��VK�9��{���щ�J0l����JJ��JJ��AAL���������e4��5�ӕ N1��P����.�LD�_�1�* �CF�"%{ `�GROU��(�1�AN4�C�#m ?REQUIR���EBU�#��6�$Tk�2$���z�܏ #�& \�AP�PR� C� 0�
$�OPEN�CLO�S�St��	i�
\��&' �Mf�p����W"-_MG߱7CB@�A���B�BRK@NOLD|@�0RTMO_5�H�p1J��P�� ������������6��1�@ �)!�#�(� ������'��+#PATH''@!6#@!��<#� � '��1SCaA���6IN�ңUCJ�[1� C0@UM�(Y ��#�"������*���*��� PAYwLOA~J2LؠOR_AN^�3L���91�)1AR_F�2LSHg2B4LO�4�!F7�#T7�#ACRL_�%�0�'�$r��H��.�$HA^�2FLEX��J!�) P�2�D��߽���0��* :����z�FG]D��`��z���%�F1]A �E�G4�F�X�j�|���BE���������� ��(��X�T*�A���@�XI�[�m�\At�T$g�QX<�=��2TX ���emX���������� ��������+	�J>+ �-�K]o|�٠AT�F�4�CELFPѪs�J� �*� JEmCTR��!�ATN�vzH�AND_VB.���1��$, $8`Fi2Av���SWu�	#-� $$M*0.�]W�lg��PZ����A��� 1�����:AK��]A�kAz��LN�]D*kDzPZ G��C�CST_K�lK�N}DY��� A����0 ��<7]A<7W1�'��d�@g`�P��������"
"J"�. M�2D%"p�H���~�ASYMj%0��� j&-��-W1�/_ �{8� �$�����/�/�/�/ 3J<�:p9�/�89�D_VI��v����V_UN!I�ӛ��cD1J���� ╴�W<��n5Ŵ�w=�4��9��?�?<�uc$�4�3�%�H����/�j��0�DIzuO���k�>�0 �`��I��A ��#���@ģ���@����IPl� 1 �[ /�ME.Qph��9�ơT}�PT� ;pG �+ Gt� ����'��T�0 �$DUMMY1���$PS_�@RMF�@  G b�'7FLA@ YP(c|���$GLB_T P�ŗ���9 P�q���2 X� z!SuT9�� SBRM �M21_V�T$_SV_ER*0O�pL����CL����AGP�O��f�GL~�EW�>�3 4H �$YrZrW@�x�A1B+�A���"j� �U&�4 8`NZ�"�w$GI�p}$&�� -� �Y�>�5 qLH {��}$F�E��NEAR(PN��CF��%PTANC��B	!JOG�@� �6.@$JOI�NTwa?pd�MSE]T>�7  x�E��HQtpS{r��up>�8�� �pU.Q?��� LOCK_F�OV06���BGLV��sGLt�TEST�_XM� 3�EMP������_�$1U&@%�w`24� Y�B��5��2�d��3���CE- ���� $K�AR�QM��TPD�RA)�����VECXn@��IU��6��{HEf�TOOL�C�2V�DRE IS�3ER6��@AC)H� 7?Ox ӦQ�29Z�H I� � @$RAIL__BOXEwa�oROBO��?��?HOWWAR�1�<_�zROLMj���:qw�jq� �@ O{_Fkp! d�tl>�9�� �R �O8B: �@�,	""�OU�;�Һ��3ơ�r�q_�$PIP��N&`H�l��@��#@CORD�EDd�p >f�fpO��� < D ��OB⁴sd����Kӕ���qSYS��ADR��f��T�CHt� = ,�8`ENo��1Ak�_�{�-$Cq_�f�VW�VA��> � � &��PREV�_RT�$ED�ITr&VSHWRBkq�֑ &R:�v��D��JA�$�a$HEAD�6�� ��z#KE:�E�CPwSPD�&JMP��L~��0R*P��?���1%&I��S�rC��pNE; �q�wTICK�C��M�13�3{HN��@ @�8 1Gu�!_GPp6���0STY'"xLO��:�2l2?�A tk 
m G3%%$R!�{�=��S�`!$@��w`���ճ���Pˠp6SQU��E��u��TERC�0��T=SUtB ����@hw&`gw�Q)�pOЌ���@IZ��{��^�PR�kюB1XsPU���E_DO���, XS�K~�AXiI�@���UR�p�GS�r� ^0�&��p_,) �ET�BPm��Jo��0Fo��0A|����Rԍ��a�;�SR�Cl >@P��b_�yUr��Y�� yU��yS��yS���UЇ �U���U���U�]��U@l[��Y�bXk�]Cm`�����YRSC��� D h�DS�~0��Q�SP���eA	Tހ���A]0,2NҿADDRES<B�} SHIF{s��_W2CH���I�Ю=q�TVsrI��E�"���a�Ce�
��
�;�VW�A��F \��q��0l|\A@�rC�_B"R{zp�ҩq��TXSCREE��Gv��1TIN!A���t{����A�b?�H T1�ЂB �����I��A��BE�y RRO������� �B��D��UE4I ��g�!p�S��R�SM]0�GUNEX0(@~Ƴ�j�S_S�ӆ@��Á։񇣣�ACY򼯂0� 2H�pU�E;�J�����@G+MT��Lֱ�A�нO	�BBL_| W�8���K ��0s�OM��LE/r��� �TO!�s�RIGHΓ�BRD
�%qCKsGR8л�TEX�@|����WIDTH��� �B[�|�<��I�_��Hi� L 	8K���_�!=r���R:�_��Yґ��)O6q�Mg0紐�U��h�Rm��LUqMh��FpERVwD �P���`�N���&�GEUR��F4P)�)� LP��(R	E%@�a)ק�a�!���f �5�6�7�8Ǣ#B�É@���t�P�fW�S@M��USR&�O �<����U�Qs�FsOC)��PRI;Q�m� :���TRIP>�m�UN����Pv��0��f%��'8���@�0 Q���.�AG �0T� �aL>q�OS�%�RPo���8�R/�A�H�L4����U¡�S�U�g��¢5��OF�F���T�}�O�� 1R����ĝS�GUN��>6�B_SUB?���N,�SRTN�`TUg2���mCOR| D�R�AUrPE�TZ�#'��VCC��	3V �AC36MFB1�f$OPG �W �(#��ASTEM�0����0PE��T3�G�X �\ ��M�OVEz�<���AN��� ���M���LIM_X��2��2�� 7�,�����ı�
��VF�`E�� }��04Y��IB�7���5S��_Rp� 2���/ WİGp+@���}СP��3�Zx# ���3����A�ݠCZ�DRID����Vy08�90�� De�MY_UBYd���6��@��!q��X��P_S���3��L�KBM,��$+0DEY(#EX�`�����UM_MUb� X����ȀUS��� ���G0`PACI���а@��:��:0,�:����RE/�3qDL�+��:[��/TARG��P�rr��R<�\ d`�H�A��$�	��AR��#SW2 ��-��@�Oz�%qA7p�yRE�U�U�01�,�HK�2]g0�qP�� N� �EAM0GW�OR���MRC]V3�^ ���O�0M�C�s	���|�REF_���x (�+T� ������p���3_RCH 4(a�P�І�hrj�NA8�5��0�_ ��2�����L@��n�@@OU ~7w6���Z��a2[��RE�p�@;0�\�c�a'2K�@S+UL��]��C��0�3^��� NT��L� 3��(6I�(6q�(3� L��Q5��Q5I�]7q��}�Tg`4D`�0|.`0�AP_HUCv�5SA��CMPz��F�6�5�5�0_�aR ��a�1I\!X�9|"�GFS��ad ���M��0p�UF�_x��B� �ʼ,RO`��Q��'����UR�3#GR�`.�3IDp���)�D�;��A��~�IN��H{D��V@AJ���S͓UW mi=�����TYLO*�5�����bt +�cPA�� �cCACH �vR�UvQ��Y��pj�#CF�I0sFR�XqT���Vn+$HO����P!A3�XBf`�(1 ���$�`VPy<� ^b_SZ313he6K3he12J�eh �chG�chWA�UMP\�j��IMG9uP�AD�iiIMRE��$�b_SIZ�$P���0 ��ASYN�BUF��VRTD�)u5tqΓOLE_C2DJ�Qu5R��C���U��vPQuEC;CUlVEMV �U<�r�WVIRC�aIuVTPG���rv1s��5qMPLAqa��v��V0�c��� C/KLAS�	�Q�"��d  �ѧ%ӑӠ�@}¾�$�Q���Ue� |�0!�rSr�T@�#0! �r�iI���m�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f � >֦3�@Sp��SLOW>�RO��ACCE���!� 9�VR�#���p:���cAD�����PAV��j�� D����M_qB"���^�JMPG ��g:�#E$SS�C��x&�vPq��h$ݲvQS�`qVN��wLEXc�i T`��sӂ��Q�FLD6 �DEsFI�3��02���:��VP2>�Vj� �A���V�4[`MV_PI s��t���A�@��FI��|�Z��Ȥ������A���A��~�GA�ߥ1 LOO��1 JCB���Xc��^`�#PLANE��R��1�F�c�����pr�M � [`�噴��S���� f����Af��R�Aw�״rtU��pRKE��d�VANC�A��.�� k���ϲ��BR_AA� l���2� ��p�#��m# h�@��O K�$��d����kЍ0OU&Aʞ"A�
p�pSK��TM@FVIEM 2�l ��P=���n� <<��dK�UMKMYK1P��`mD�ȟ�CU��z#AU��o $���TIT�$P�R����OP����VSHIF�r�p`J�Qsԙ�fO�xE$� _R�`U �#����s��q����@��G�"G�޵'�T��$�SCO{D7�CNTQ i�l�>a�-�a� ;�a�H�a�V���1�*+�2u1��D�����  � SMO"�Uq��a�JQ���K��a_�R[�r�n�*@LIQ�AA/`/�XVR��s�n�yTL���ZABC�Ct�t�c�
LїZIP��u���L�VbcLn"���M�PCFx�v:�$��� ���DMY_�LN�������@y�w� Ђ(a�u� MC�M�@CbcCART�_�DPN� '$J71D��=�NGg0Sg0�BUX�W� ��UXEUL|ByX����	�����x �	���m�YH�D>b  y 80�֞�0EIGH�3n�?�(� H����$z� ���|�����$B� Kd'��_��L3��RVS�F`���OVC�2'�$|�>PD&��
q���5D��TR�@ �Vc��SsPHX��!{ ,� �*<�$R�B2 2 ���C!��  ���V+L�b*c%Rg!`+g"�`V*~�,8�?�V+ �/V.�/�/?�/�/V(7%3@/R/d/v/�/6? �/�/�?�?�?O4OOION;4]?o?�?�?�? SO�?�?�O_�O0_Q_8_f_N;5zO�O�O�O �Op_�O_o8o�_MonoUo�oN;6�_�_�_ �_�_�oo%o4U j�r�N;7�o�o �o�o�o� BQ�r�@5���������N;8� ����Ǐ=�_�n����R���ş��ڟN;Gw � џ
�
����?���W� i�{�������ï�.��������A��d W�<�N�|�������Ŀ ֿ�ޯ���0�B� _�R�d�꿤϶����� ��������*�L�^� �rτ�
��������� ���&�8�J�l�~�w `ҟ @�Ѐ�����ߩ��-� ���&�,���9�{� ����a����������� ����A'Y� ������� �a#1�
���N;_MODE  y��S ��[�Y�B���
/�\/*	|/�/R4CW�ORK_AD�	��
T1R  ����� �/� _I�NTVAL�+$���R_OPTIO�N6 �q@V�_DATA_GR�P 27���D��P�/~?�/�?�9� �?�?�?�?OO;O)O KOMO_O�O�O�O�O�O �O_�O_7_%_[_I_ _m_�_�_�_�_�_�_ �_!ooEo3oioWoyo �o�o�o�o�o�o�o /eS�w� ������+�� O�=�s�a�������͏ ���ߏ��9�'�I��o�]�����$SA�F_DO_PUL�S� �~������C?AN_TIM�����ΑR �+�+Ƙ�"��5�;#U!P"�1!��� �?E�W�i� {�����.�ïկ���X��'(~�T"2F���dR�I�Y��2�o+@a얿�����)�u��� k0ϴ���_ ��  �T� � �2�D�)�T D��Q�zό� �ϰ���������
�� .�@�R�d�v߈ߚ�/<V凷������߽��R�;��o �W�p��
�?t��Diz$�~ �0 � �T" 1!�������� ����������*�<� N�`�r����������� ����&8J\ n���������"4FX �� ࿁������ �/`4�=/O/a/s/ �/�/�/�/�/�/�!!/ �0޲k�ݵu�0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ ok $o6oHoZolo~o�o�o �o�o1/�o�o 2 DVhz�/5?�� ������&�8� J�\�n���������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u��� ���`Ò�ϯ ����)�;�M�_� q���������˿ݿ�� ����3� ����&2,��	12345678v��h!B!�U�2�Ch���0� �ϵ����������!� 3�9ѻ�\�n߀ߒߤ� �����������"�4� F�X�j�|�h�K߰��� ������
��.�@�R� d�v������������� ��*<N`r ������� &��J\n�� ������/"/ 4/F/X/j/|/;�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �/�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_�?L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o=_�o �o�o�o�o�o 2 DVhz�����h������u�o�.�@�R���Cz � B��   ����2&� � �_�
���  	�_�2�Տ���,�_�p������ďi�{�������ß ՟�����/�A�S� e�w���������N�� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�_�����<v�_��$SC�R_GRP 1
�+� +�� �t ��� ���	 ��������� �������_�����Ϝ)�a����&�DE� DW8���l��&�G�CR-3�5iA 9012�34567890���M-20��8~��CR35 ��F:�
��������������:֦�Ӧ��G���&������	���]�o����:���H���>�����������&���ݯ:��j����g�X�����B�t�����������A����  1@�`��@� (' ?�=��Ht�P�
��F@ F�`z�y����� � �$H���Gs^p��B� �7��/�0// -/f/Q/�/u/�/�/�/�8���P�� 7%?�����"?W?-2?<�	���-<@H�1�?t�ȭ7�������?-4A, �&E@�<�I@G�B-1 3OZOlO-:HA�H�O�O.|O P�B(�B�O��O_��EL_DE�FAULT  ~����`�SHOTSTR�#]A7RMIPOWERFL  i�z/UYTWFDO$V� /URRVENT 1�����NU L!DU�M_EIP_-8��j!AF_IN�E#P�_-4!FT$�_->�_;o!��`o� �*o�o!RPC_MAIN�o�jh�vo�o�cVIS�oii��o!TMPpPU�Yd�k!
PMON_�PROXYl�Ve Z�2r��]f���!RDM_SR�V��Yg�O�!�R��k��Xh>���!%
�`M��\i����!RLSYNC��-98֏3�!gROS�_-<�4"���!
CE4pMT'COM���Vkn�˟{!	��CONS̟��Wl���!��WOASRC��Vm�vc�!��USBd��XnR���Noӯ��� ����!��E��i�0����WRVICE_�KL ?%�[ �(%SVCPR#G1��-:Ƶ2ܿ�"˰3�	�˰4,�1�"˰5T�Y�˰6|ρ�˰7�ϩ�˰�����	9����ȴf�!�˱ οI�˱��q�˱ϙ� ˱F���˱n���˱�� �˱��9�˱��a�˱ ߉��7߱��_��� �����)���� Q����y��'��� O����w����� ����˰��İd �c������ =(as^�� ����/�/9/ $/]/H/�/l/�/�/�/ �/�/�/�/#??G?2? k?V?}?�?�?�?�?�? �?O�?1OCO.OgORO �OvO�O�O�O�O�O	_��O-_��_DEV ��Y�MC�:5Xd�GTG�RP 2SVK ���bx 	� 
+ ,�PK 5_�_ �T�_�_�_o�_'o9o  o]oDo�ohozo�o�o �o�o�o�o5{�_ g������ ����?�&�c�u� \�������Ϗ���J \)���M�4�q���j� ����˟ݟğ��%� ��[�B��f����� �ٯ�������3�� W�i�P���t���ÿ�� �ο���A�(�e� L�ί��RϿ��ϸ��� ��� ��O�6�s�Z� �ߩߐ��ߴ������ '�~ϐ�]���h�� ������������5� �Y�@�R���v����� ����@�	��?& cu\����� ���;M4q X�������/ �%//I/[/B//f/ �/�/�/�/�/�/�/�/ 3??W?�L?�?D?�? �?�?�?�?O�?/OAO (OeOLO�O�O�O�O�O��O�O�O_iV �N�Ly�6 * �		S=>��+�c"_VU@Tn_Y_B����B�2�J�j~Q´~_g_�_��Q%JOGGI�NG�_�^7T(?Vj�Z�Rf��Y���/e�_%o7e�Tt�]/o�o{m�_�o�m ?Qi�o�o;)Kq%��o�}os ������9�{ `��)���%���ɏ�� �ۏ�S�8�w��k� Y���}���ş���+� �O�ٟC�1�g�U��� y�������'���� 	�?�-�c�Q���ɯ�� ��w���s����;� )�_ϡ���ſOϹϧ� ��������7�y�^� ��'ߑ�ߵߣ����� ���Q�6�u���i�W� ��{������=�� M���A�/�e�S���w� ����������� =+aO������ u���9' ]���M��� ���/5/w\/� %/�/}/�/�/�/�/�/ =/"?4?�/?�/U?�? y?�?�?�??�?9?�? -OO=O?OQO�OuO�O �?�OO�O_�O)__ 9_;_M_�_�O�_�Os_ �_�_o�_%oo5o�_ �_�o�_[o�o�o�o�o �o�o!coH�o{ ������;  �_�S�A�w�e��� ����я���7���+� �O�=�s�a������ П�����'��K� 9�o�������_���[� ɯ���#��G���n� ��7���������ſ�� ��a�Fυ��y�g� �ϋϭϯ�����9�� ]���Q�?�u�cߙ߇� ����%���5���)�� M�;�q�_���߼��� �������%��I�7� m������]������� ����!E��l�� 5������� _D�we� ����%
//� ��=/s/a/�/�/�/ ��/!/�/??%?'? 9?o?]?�?�/�?�/�? �?�?O�?!O#O5OkO �?�O�?[O�O�O�O�O _�O_sO�Oj_�OC_ �_�_�_�_�_�_	oK_ 0oo_�_co�_so�o�o �o�o�o#oGo�o; )_Mo����o ����7�%�[� I�k���������� ُ���3�!�W���~� ��G�i�C����՟� ��/�q�V������w� �������ѯ�I�.� m���a�O���s����� ��߿!��E�Ͽ9�'� ]�Kρ�oϑ����� Ϸ����5�#�Y�G� }߿Ϥ���m���i��� ���1��U��|�� E���������	��� -�o�T������u��� ��������G�,k� ��_M�q��� ����%[ Im���	� ��//!/W/E/{/ ��/�k/�/�/�/�/ 	???S?�/z?�/C? �?�?�?�?�?�?O[? �?RO�?+O�OsO�O�O �O�O�O3O_WO�OK_ �O[_�_o_�_�_�__ �_/_�_#ooGo5oWo }oko�o�_�oo�o�o �oC1Sy�o ��oi����� 	�?��f�x�/�Q�+� ��Ϗ�����Y�>� }��q�_�������˟ ���1��U�ߟI�7� m�[�}����ǯ	�� -���!��E�3�i�W� y�ϯ��ƿ������ ��A�/�eϧ���˿ UϿ�Q��������� =��dߣ�-ߗ߅߻� ���������W�<�{� �o�]������� ��/��S���G�5�k� Y���}����������� ����C1gU� �����{���� 	?-c���S ������/;/ }b/�+/�/�/�/�/ �/�/�/C/i/:?y/? m?[?�??�?�?�??  O??�?3O�?COiOWO �O{O�O�?�OO�O_ �O/__?_e_S_�_�O �_�Oy_�_�_o�_+o o;oao�_�o�_Qo�o �o�o�o�o'ioN `9���� ��A&�e�Y�G� i�k�}�����׏��� =�Ǐ1��U�C�e�g� y����֟���	��� -��Q�?�a���ݟ�� ퟇��ϯ��)�� M���t���=���9��� ݿ˿��%�g�Lϋ� ��mϣϑϳ����� ��?�$�c���W�E�{� iߟߍ߯������;� ��/��S�A�w�e�� �����������+� �O�=�s������c� ����������'K ��r��;���� ���#eJ� }k�����+ Q"/a�U/C/y/g/ �/�/�//�/'/�/? �/+?Q???u?c?�?�/ �?�/�?�?�?OO'O MO;OqO�?�O�?aO�O �O�O�O__#_I_�O p_�O9_�_�_�_�_�_ �_oQ_6oHo�_!o�_ io�o�o�o�o�o)o Mo�oA/QSe�����%{,p��$SERV_MA_IL  +u!���+q�OUTPU]T�$�@��RV 2�v  $� (�q�}���SAVE7�(�TO�P10 2W�� d 6 *_�π(_������ #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽݷ毅YP��'�FZN_CFG �u'$�~����?GRP 2�D�� ,B   A�[�+qD;� B�\��  B4~��RB21��HELL��u��j��k�2�����%RSR�������
�C� .�g�Rߋ�v߈��߬߀����	���-�?�Q�_�  �_�%Q���_���,p�����ޖ�g�2�,pd����HK ;1�� ��E� @�R�d����������� ������*<e�`r���OMM ������FTOV_ENB�_����HOW_REG_�UI�(�IMIO/FWDL� �^�^)WAIT���$V1�^�NT�IM���V�A�_)_UNI�T����LCT�RYB�
�MB�_HDDN 2W� 2�:%0  �pQ/�qL/^/�/�/�/��/�/�/�/�"!ON�_ALIAS ?5e�	f�he�A? S?e?w?�:/?�?�?�? �?�?OO&O8OJO�? nO�O�O�O�OaO�O�O �O_"_�OF_X_j_|_ '_�_�_�_�_�_�_o o0oBoTo�_xo�o�o �o�oko�o�o, �oPbt�1�� �����(�:�L� ^�	���������ʏu� � ��$�Ϗ5�Z�l� ~���;���Ɵ؟��� �� �2�D�V�h���� ����¯ԯ���
�� .�ٯR�d�v�����E� ��п���ϱ�*�<� N�`�r�ϖϨϺ��� w�����&�8���\� n߀ߒߤ�O������� ����4�F�X�j�|� '����������� �0�B���f�x����� ��Y��������� >Pbt��� ���(:L �p����c� � //$/�H/Z/l/ ~/)/�/�/�/�/�/�/�? ?2?D?V?]3�$�SMON_DEF�PRO ����1 �*SYSTE�M*0m6REC�ALL ?}9� ( �}tp�disc 0=>�147.87.1�49.40:11�304 4 �>0�632 �1�951�72]?O+M}t�pconn 0 ��?�?�?�?�O�O4G
�xyzrate 61 JO\OnO�O_d#_6E�G�=28�@��O�O_�_�_�L11 GMY_k_}_o o3_E_@�_�_�_�o�o1J�? Sh\ono�o#6O�o �o�o�o���_�QJ \n��#�6oHoZo ��������AJ�\��n����#�6�H�9548ݏ�������oK� \�n����#�6�ȟڟ�������4�8�copy frs�:orderfi�l.dat vi�rt:\tmpback\ǟ[�y�
���/�/��mdb:*.*ԯ�����l��7�3x��:\H� ɰZ�[�s����(�;�4��aǿٿV���� �ϩϼKJ�\�nπ���#�6�H�6284  ����ߓߥ߸J�\� n߀��#�6�H����� �ߏ�ﴟ�>Y�\�n� ���#�6��������� �������NW�i�{�01�C�Ղ12����  ����ȏZl~ !4F���� ���įM�Nx	// .�@��S�/�/�/ ��H/��Xs/�/?(? ;��/�/[�/?�?�? ��P]?o?�?O$O7� �?�?�?�?�O�O��~ XOjO|O__2DV �O�O�_�_�O�T_f_ x_	oo._@_�_�_�_ o�o,o��Y/to�o )</�o`/�o����`�$SNPX�_ASG 2�����q�� P 0 '�%R[1]@g1.1��y?��s%�!��E�(�:�{� ^�������Տ��ʏ� ��A�$�e�H�Z��� ~���џ����؟�+� �5�a�D���h�z��� ��ů�ԯ���
�K� .�U���d�������ۿ ������5��*�k� N�uϡτ��ϨϺ��� ���1��U�8�Jߋ� nߕ��ߤ�������� ��%�Q�4�u�X�j�� ������������;� �E�q�T���x����� ������%[ >e�t���� ��!E(:{ ^������/ �/A/$/e/H/Z/�/ ~/�/�/�/�/�/�/+? ?5?a?D?�?h?z?�? �?�?�?�?O�?
OKO .OUO�OdO�O�O�O�O �O�O_�O5__*_k_ N_u_�_�_�_�_�_�_ �_o1ooUo8oJo�o�no�o�o�d�tPAR�AM �u��q �	��jP��d9p�ht���pOFT_KB_?CFG  �c�u��sOPIN_SI/M  �{vn���p�pRVQS�TP_DSBW~�r"t�HtSR }Zy � &!p�INGS EL_O5SEM���v�TOP_ON_ERR  uCy8��PTN Zu^k�A4�R��_PR�D��`V�CNT_GP 2�Zuq�!px 	 r��ɍ���׏��w�VD��RP 1�i p�y��K�]� o���������ɟ۟� ���#�5�G�Y���}� ������ůׯ���� �F�C�U�g�y����� ����ӿ��	��-� ?�Q�c�uχϙϫ��� ��������)�;�M� _�qߘߕߧ߹����� ����%�7�^�[�m� ������������ $�!�3�E�W�i�{��� ������������ /ASew��� ����+= Ovs����� ��//</9/K/]/ o/�/�/�/�/�/�/? �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O�O)�PRG_CO7UNT8v�k�GuNKBENB��FEMpC�:t}O_UPD 1}�{T  
4O r�O�O�O__!_3_ \_W_i_{_�_�_�_�_ �_�_�_o4o/oAoSo |owo�o�o�o�o�o�o +TOas �������� ,�'�9�K�t�o����� ����ɏۏ����#� L�G�Y�k��������� ܟן���$��1�C� l�g�y���������ӯ ����	��D�?�Q�c� ��������ԿϿ�� ��)�;�d�_�q�=L�_INFO 1޵E�@ �2@���������� ���8@�o6���W��´*�H@YS�DEBUGU@�@���d�If�SP_PwASSUEB?xۿLOG  ��ʠC��Qؑ�  ���A��UD1�:\��Uߦ�_MPAC�ݵE&�8�A���V� �A�SAV �!�������X����SVZ�TEM�_TIME 1"����@ 0��e�X�X�X�����$T1SVGUNYS�@VE'�E���ASK_OPTICONU@�E�A�A+��_DI��qOG�BC�2_GRP 2#�I�����@�  �C���<Ko�CFGg %z��� �����`��1�. >dO�s�� �����*N 9r]����� ��/�8/#/\/n/ ��Z+�/Z/�/�/H/�/ ?�/'??K?]�k?=� @0s?�?�?�?�?�?�? O�?OO)O_OMO�O qO�O�O�O�O�O_�O %__I_7_m_[_}__ �_�_�X� �_�_oo /o�_SoAoco�owo�o �o�o�o�o�o= +MOa���� �����9�'�]� K���o���������ɏ ���#��_;�M�k�}� �������ß�ן� �1���U�C�y�g��� ������������	� ?�-�c�Q�s������� ���Ͽ����)� _�Mσ�9��ϭ����� ��m���#�I�7�m� ߑ�_ߵߣ������� ����!�W�E�{�i� ������������� �A�/�e�S�u�w��� ����������+= O��sa���� ���9'] Kmo����� ��#//3/Y/G/}/ k/�/�/�/�/�/�/�/ ??C?��[?m?�?�? �?-?�?�?�?	O�?-O ?OQOOuOcO�O�O�O �O�O�O�O__;_)_ __M_�_q_�_�_�_�_ �_o�_%oo5o7oIo omo�oY?�o�o�o�o �o3!CiW� ������� �-�/�A�w�e����� �����я���=� +�a�O���s������� ߟ͟��o�-�K�]� o�ퟓ�����ɯ����צ��$TBCS�G_GRP 2&�ץ� � �� 
 ?�  6�H�2�l�V� ��z���ƿ��������(�d��E+�?�	 HC{���>���G�����C�  A�.�e�q�C��>ǳ33��S�/]϶�Y���=Ȑ� C\  �Bȹ��B���>�����P���B�Y�z��L�H�0�$����J�\�n�����@�Ҿ��������߀=�Z�%�7����?�3�����	V�3.00.�	cwr35��	*�����
�������� �3��4�   {�CT�v�}��J2�)�������CFG +ץe'� *������qI���� .<
�<bM�q �������( L7p[�� ����/�6/!/ Z/E/W/�/{/�/�/�/ �/.�H��/??�/L? 7?\?�?m?�?�?�?�? �? OO$O�?HO3OlO WO|O�O����Oӯ�O �O�O!__E_3_i_W_ �_{_�_�_�_�_�_o �_/oo?oAoSo�owo �o�o�o�o�o�o+ O=s�E��� Y�����9�'� ]�K�m�������u�Ǐ ɏۏ���5�G�Y�k� %���}�����ßşן ���1��U�C�y�g� ������ӯ������ 	�+�-�?�u�c����� �����Ͽ���/� A�S�����qϓϕϧ� �������%�7�I�[� ��mߣߑ߳����� �߷��3�!�W�E�{� i����������� ��A�/�e�S�u��� ������������ +aO�s�� e�����'K 9o]���� ���#//G/5/k/ }/�/�/[/�/�/�/�/ �/??C?1?g?U?�? y?�?�?�?�?�?	O�? -OOQO?OaO�OuO�O �O�O�O�O�O___ M_�e_w_�_3_�_�_ �_�_�_oo7o%o[o moo�oOo�o�o�o�o �o!3�o�oiW �{������ �/��S�A�w�e��� ����я������� =�+�M�s�a������� ��ߟ�_	���_ן ]�K���o�������ۯ ɯ���#���Y�G� }�k�����ſ׿���� ����U�C�y�g� �ϋ��ϯ�������� 	�?�-�c�Q�s�u߇� �߫��������)�� 9�_�M����/���� i������%��I�7� m�[������������� ������EWi{ 5������� �A/eS�w �����/�+/ /O/=/_/a/s/�/�/ �/�/�/�/?'?��?? Q?c??�?�?�?�?�? �?�?O�?5OGOYOkO�)O�O}O�O�O�O�N s �@S V�_R�$TBJO�P_GRP 2,��E� / ?�V	-R4S�.;\��@|�u0{SPU >���UT @��@LR	 �C�� �Vf  C����ULQLQ>�33��U�R����U�Y?~�@=�ZC��P׌�ͥR��P � B��W$o/gC���@g�dDb�^���eeao�P�&ff�e=�7L3C/kaB o�o�P��P�efb-C�p��^g`�d�o��PL�Pt<�eVoC\  �Q@�'p}�`�  A�o�L`�_wC�BrD�S�^�]�_�S~�`<PB��P0�anaa`C�;�`L�w�aQoxp��x�p:��XB$4'tMP@�PCHS��n���=�P����trd<M�gE�2pb ����X�	��1�� )�W���c�������� ����󟭟7�Q�;�PI�w���;d�Vɡ��U	V3.00�RScr35QT�*�QT�A�� �E�'E�i��FV#F"w�qF>��FZ�� Fv�RF�~�MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
�D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt���ٵ=�_t��V �R�p�V9� ]ESTP�ARtp�HFP*SH�R\�ABLE 1%/;[%�SG��Q �W�G�G�GȨ WQG�	G�
G��GȖ�QG�G�8G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ߱���w�S]�CS !ڄ�� �����������&� 8�J�\�n��������� ���� ]\�`��	� �(�:�����
��.��@�w�NUM  ��EEQ�P�	P ۰ܰw�_CFG 0��)r-P�IMEBF_TT�b��CSo�,VER�ڳ-B,R 1=1;[ 8��R��@� �@&   �������/ /)/;/M/_/q/�/�/ �/�/�/?�/?J?%? 7?M?[?m?>�@�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_l_�Y�@cY�MI_CWHAN8 c c�DBGLV��:�cX�	`ETHER_AD ?f�\`��?�_uo�oQ��	`ROUTV!�	
!�d�o�lSN�MASKQhcba255.uߣ'�9ߣY�OOLOF/S_DIb��U;i�ORQCTRL �2		�Ϸ~T �����#�5�G� Y�k�}�������ŏ׏ �����.��R�V��PE_DETAI�/h|zPGL_CONFIG 8�	����/cel�l/$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c� u�����(���ϯ�� ����;�M�_�q��� ��$�6�˿ݿ��� %ϴ�I�[�m�ϑϣ� 2����������!߰� ��W�i�{ߍߟ߱�%}F�������/�A��C�i�H�Eߞ�� ��������?��.�@� R�d�v���������� ������*<N` r������ �&8J\n� �!�����/ �4/F/X/j/|/�// �/�/�/�/�/??�/ B?T?f?x?�?�?+?�? �?�?�?OO�?>OPO�bOtO�O�O�O����User Vi�ew ��}}12�34567890 �O�O�O_#_5_=T�P,��]_���I2�I:O �_�_�_�_�_�_X_j_�B3�_GoYoko}o�o�o o�op^46o�o�1CU�ovp^5 �o�����	�h*�p^6�c�u����� �����ޏp^7R�� )�;�M�_�q�Џ��p^8�˟ݟ���%����F�L� lCamera�J ��������ӯ���E~��!�3��OM�_�`q��������y  e� �Yz���	��-�?�Q� ��uχϙ�俽���������>��e�5i�� c�u߇ߙ߽߫�d��� ���P�)�;�M�_�q� ��*�<��i������� ��)���M�_�q��� ��������������<� û��=Oas�� >����*' 9K]f�Q��� ����/�%/7/ I/�m//�/�/�/�/ n<��^/?%?7?I? [?m?/�?�?�? ?�? �?�?O!O3O�/<׹� �?O�O�O�O�O�O�? �O_!_lOE_W_i_{_�_�_FOXG9+_�_�_ oo(o:o�OKopo�o )_�o�o�o�o�o 
��	g�0�oM_q ���No����o �%�7�I�[�m�& l�n��Ə؏����  ��D�V�h������� ��ԟ柍�g�ڻ}� 2�D�V�h�z���3��� ¯ԯ���
��.�@� R���3uF�鯞���¿ Կ������.�@ϋ� d�vψϚϬϾ�e�w� ��U�
��.�@�R�d� ψߚ߬��������� ��*���w���v� �������w���� �c�<�N�`�r����� =�w��-����� *<��`r�����������  ��1CUgy��������   -/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E_W_i_�  
���(  �%( 	 y_�_�_�_ �_�_�_o	o+o-o?o@uoco�o�o�o�Z* �Q&� J\n������o ���9�(�:�L� ^�p���������܏ � ��$�6�}�Z�l� ~�ŏ����Ɵ؟��� C�U�2�D�V���z��� ����¯ԯ���
�� c�@�R�d�v������ ��п�)���*�<� N�`ϧ����ϨϺ�� ������&�8��\� n߀��Ϥ߶������� ��E�"�4�F��j�|� ����������� �e�B�T�f�x����� ��������+�, >Pb������� ���(o� ^p������ � /G$/6/H/�l/ ~/�/�/�/�//�/�/ ?U/2?D?V?h?z?�?�/�`@ �2�?�?��?�3�7�P��!�frh:\tpg�l\robots�\m20ia\c�r35ia.xml�?;OMO_OqO�O�O�O�O�O�O�O �� �O_(_:_L_^_p_�_ �_�_�_�_�_�O�_o $o6oHoZolo~o�o�o �o�o�o�_�o 2 DVhz���� ��o�
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟�ݟ� �&�8�J�\�n����� ����ȯߟٯ���"� 4�F�X�j�|��������Ŀ־�8.1 ��?@88�?�ֻ�ֿ�3�5�G� iϓ�}ϟ��ϳ����� ���5��A�k�U�w���߿��$TPGL�_OUTPUT �;�!�! ��������,� >�P�b�t����� ��������(�:�L�@^�p�������������2345678901�������� �"��BTfx� �4�����
}$L^p�� ,>��� //$/ �2/Z/l/~/�/�/:/ �/�/�/�/? ?�/�/ V?h?z?�?�?�?H?�? �?�?
OO.O�?<OdO vO�O�O�ODOVO�O�O __*_<_�OJ_r_�_ �_�_�_R_�_�_oo &o8o�_�_no�o�o�o �o�o`o�o�o"4 F�oT|����\��}�����0�B�T�e�@������� ( 	 �� Џ������<�*� L�N�`���������ޟ ̟���8�&�\�J� ��n���������ȯ���"�������*�X� j�F�����|�¿Կ�� C���ϱ�3�E�#�i� {�忇ϱ�S������� ���/ߙ�S�e�߉� ��y߿���;����� ��=�O�-�s���ߩ� ��]��������'��� �]�o���������� ��E�����5G% W}������g� ��1�Ug	 w�{��=O	/ /�?/Q///u/�/� �/�/_/�/�/�/�/)? ;?�/_?q??�?�?�? �?�?G?�?O�?OIO [O9OO�O�?�O�OiO �O�O�O!_3_�O_i_ {__�_�_�_�_�_�R��$TPOFF_�LIM >�op:���mqbN_�SV`  l��jP_MON M<6�dopop�2l�aSTRTC�HK =6�f�� bVTCOMP�AT-h�afVWV_AR >Mm�h.1d �o �oop�`ba_DEFPROG %|j�%TISCHZ�UZAUN	�j_DISPLAY`�|n"rINST_M�SK  t| ~^zINUSER�o�dtLCK�|}{QUICKMEJp�"roSCRE�p6�~�btpscdt��q��b*�_.�S�T�jiRACE_�CFG ?Mi��d`	�d
?�~u�HNL 2@|i����k r͏ߏ ���'�9�K�]�w�ITEM 2A��� �%$1234567890����  =<��П��  !���p��=��c��^��� �������.���R�� v�"�H�ί��Я��� ���*�ֿ���r�2� ������4�޿�ϰ��� &���J�\�n���@ߤ� d�v��ς������4� ��X��*��@��� ���ߨ�������T� ��x������l��� �����,�>�P����� ��FX��d����� �:�p"� �o�����F 6HZt~��N/ t/�/��// /2/�/ V/?(?:?�/F?�/�/ �/j?�??�?�?R?�? v?�?QO�?lO�?�O�O O�O*O|O_`O _�O 0_V_h_�Ot_�O__ �_8_�_
oo�_@o�_ �_�_Lodo�_�o�o4o �oXojo3�oN�or���o��s�S��B���z�  h��z ��C�:y
 P�v�]�����UD1:\������qR_GRP �1C��� 	 @Cp���$� �H�6�l�Z��|������f���˟���ڕ?�  
���<�*� `�N���r�������ޯ ̯��&��J�8�Z����	�u�����sS�CB 2D� �����(�:�L��^�pς��|V_CONFIG E����@����ϖ�OUT?PUT F�������6�H�Z� l�~ߐߢߴ������� �����#�6�H�Z�l� ~������������ ��2�D�V�h�z��� ������������
� .@Rdv��� ����)< N`r����� ��//%8/J/\/ n/�/�/�/�/�/�/�/ �/?!/4?F?X?j?|? �?�?�?�?�?�?�?O O/?BOTOfOxO�O�O �O�O�O�O�O__+O >_P_b_t_�_�_�_�_ �_�_�_oo'_:oLo ^opo�o�o�o�o�o�o �o $����!�b t������� ��(�:�-o^�p��� ������ʏ܏� �� $�6�G�Z�l�~����� ��Ɵ؟���� �2� D�U�h�z�������¯ ԯ���
��.�@�Q� d�v���������п� ����*�<�M�`�r� �ϖϨϺ�������� �&�8�J�[�n߀ߒ� �߶����������"� 4�F�W�j�|���� ����������0�B� S�f�x����������� ����,>Pa� t��������(:L/x���k}gV� K���//&/8/ J/\/n/�/�/�/W�/ �/�/�/?"?4?F?X? j?|?�?�?�?�/�?�? �?OO0OBOTOfOxO �O�O�O�?�O�O�O_ _,_>_P_b_t_�_�_ �_�O�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����o� ��� �2�D�V�h� z��������ԏ��� 
��.�@�R�d�v��� ������Ϗ����� *�<�N�`�r������� ��˟ޯ���&�8� J�\�n���������Ż��$TX_SCR�EEN 1G�g�}�ipnl/��gen.htmſ�*��<�N�`ϽPa�nel setupd�}�dϥϷ����������ω�6�H� Z�l�~ߐ�ߴ�+��� ����� �2�߻�h� z������9�g�]� 
��.�@�R�d���� �����������}� ��<N`r�� ;1��&8 �\��������QȾUALRM_MSG ?��� �Ȫ-/?/ p/c/�/�/�/�/�/�/��/??6?)?Z?%S�EV  -��6"ECFG �I��  �ȥ@�  A�1 �  B�Ȥ
  [?ϣ��?OO%O7O IO[OmOO�O�O�G�1�GRP 2J�;; 0Ȧ	 �?�O� I_BBL_N�OTE K�:T��lϢ��ѡ�0RDEF�PRO %+ (%N?u_Ѡc_�_�_ �_�_�_�_o�_o>o�)oboMo�o\INU?SER  R]�O��oI_MENHI�ST 1L�9  �( _P���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1�oCUgy�)
13/������p0��uedi�t(rTISCHZUZAUN�Q�c� u��z|o����ʏ܏�  ���$�6�H�Z�l�~� �����Ɵ؟����� ��2�D�V�h�z���� ��¯ԯ���
��h9R q��B�T�f�x����� ����ҿ����ϩ� >�P�b�tφϘ�'�9� ��������(߷�L� ^�p߂ߔߦ�5����� �� ��$����Z�l� ~����C������� � �2��/�h�z��� ������������
 .@��dv��� ��_�*< N�r����� [�//&/8/J/\/ ��/�/�/�/�/�/i/ �/?"?4?F?X?C�U� �?�?�?�?�?�?�/O O0OBOTOfO�?�O�O �O�O�O�O�O�O_,_ >_P_b_t__�_�_�_ �_�_�_�_o(o:oLo ^opo�oo�o�o�o�o �o �o$6HZl ~i?{?����� �2�D�V�h�z��� �-�ԏ���
�� ��@�R�d�v�����)� ��П��������� N�`�r�������7�̯ ޯ���&���J�\��n����������$�UI_PANED�ATA 1N����ڱ � 	�}/f�rh/cgtp/�widedev.stm���%�7�I�>Y�)priρ�@�}�ϩϻ�������� )�)��M�4� q߃�jߧߎ������߀���%�7��[�7����   }�S&�Ϙ�� ��������E����:� L�^�p���������� ������$H/ l~e������o� ݰܳ7�< N`r����-� ��//&/8/�\/ n/U/�/y/�/�/�/�/ �/?�/4?F?-?j?Q? �?�?%�?�?�?O O0O�?TO�xO�O�O �O�O�O�OKO_�O,_ _P_b_I_�_m_�_�_ �_�_�_oo�_:o�? �?po�o�o�o�o�oo �o sO$6HZl ~�o������ � �2��V�=�z��� s�����ԏGoYo� .�@�R�d�v�ɏ�� ��П������<� N�5�r�Y�������̯ ���ׯ�&��J�1� n�������ȿڿ� ���c�4ϧ�X�j�|� �Ϡϲ���+������ ��0�B�)�f�Mߊߜ� ���ߧ������� ��P�b�t������ ����S���(�:�L� ^����i��������� �� ��6Zl�S�w�'�9�}����"4FX) �}��l���� �/j'//K/2/D/ �/h/�/�/�/�/�/�/ �/#?5??Y?��C�=���$UI_POSTYPE  C��� 	 �e?�?�2QUICKMEN  �;��?�?�0REST�ORE 1OC��  �	L?��6OCC1O��maO�O�O�O�O�OuO �O__,_>_�Ob_t_ �_�_�_UO�_�_�_M_ o(o:oLo^oo�o�o �o�o�o�oo $ 6H�_Ugy�o� ����� �2�D� V�h��������ԏ ����w�)�R�d� v�����=���П��� ���*�<�N�`�r�� ������ޯ��� &�ɯJ�\�n��������G�ȿڿ�����7S�CRE�0?�=�u1sc+@�u2K�3K�4K�5*K�6K�7K�8K��2�USER-�2�D�k�sMì�3��4��5*��6��7��8���0�NDO_CFG �P�;� ��0PD�ATE ���?None�2���_INFO 1Q2C�@��10%�[� ��Iߊ�m߮��ߣ��� �������>�P�3�t����i���<-�OFF�SET T�= �ﲳ$@������1� ^�U�g���������� ������$-ZQ cu���?�
�����UFRAME � ����*�RTOL_ABRT	�(�!ENB*G�RP 1UI�1?Cz  A��~���~��������0UJ�9?MSK  M@�Z;N%8�%���/�2VCCM��YV�ͣ#RG�#Y�9Q���/����D��BH�p71C�2��3711?�C0�$MRf2_�*S��Ҵ�	���~?XC56 *�?�6����1$�5����A@3C��. ��8�?��O@OKOx1FOsO�5��51��_O�O�� B����A2�D WO�O7O_�O8_#_\_ G_�_k_}_�__�_�_��_�_"o�OFoXo�%TCC�#`mI1�i�괰��� GFSv��2aZ; �| �2345678901�o�b�����o���!5a�4BwB��`56 311:�o=L�Br5v1�1~1 �2��}/��o�a�� #�GYk}�p� ������ُ�1� C�U�6�H���5�~����ߏ���	���4�dS�ELEC)M!v1�b3�VIRTSYNC�� ���%��SIONTMOU4������F��#�bU��U��(u FR:�\H�\�A\�� �� MC���LOG��   7UD1��EX�����' B@ �����̡m��̡ / OBCL�1�H�� �  =	� 1- n6  -������[��,S�A�`=���ԗ��ˢ��TRAIN⯞b�a1l�E
0d�$j�T2cZ; (aE2ϖ�i ��;�)�_�M�g�qσ� �ϧ��������	���F�STAT d�m~2@�zߌ�*j$�i߾��_GE�#enZ;�`0�
� �02��HOMIN�� fU��UC� ~�����БC�g��X���JMPER�R 2gZ;
  ��*jl�V�7���� ����������
��2��@�q�d�v�B�_ߠR�E� hWޠ$LEXr��iZ;�a1-e���VMPHASE � 5��c&��!OcFF/�F�P2n��j�0�㜳�E1@��0ϒE1!1?Gs33�����ak�/�kxk䜣!W�m[�䦲�[����8o3;�  [i{���� /�O�?/M/_/ q/��/��//�/'/ 9/�/=?7?I?s?�/�? �/�/�?�??Om?O %O3OEO�?�?�O�?�O �O�?�O�O�O__gO \_�OE_�O�_�O�O/_ �_�_�_oQ_Fou_�_ |o�o�_�oo�o�o�o �o;oMo?qof-�o I�����7 �[P������� ��ˏ��!�3�(�:� i�[�ŏg�}�������TD_FILTE:W�n�� �ֲ:���@���+�=�O� a�s���������֯ �����0�B�T�f��x���SHIFTM�ENU 1o[�<��%��ֿ����ڿ ����I� �2��V� hώ��Ϟϰ��������3�
�	LIVE�/SNAP'�v�sfliv��E��{��ION * yUb�h�menu~߀������ߣ���p���	����E�.�S�50�s�P�@� ���AɠB8z�Bz��}��x�~�P�� ���M�Eb���<�0�֔�MO��q���z��WAITDINEND������sOK1�OUT�r��SD��TIM����o�G���#����C���b������R?ELEASE����f��TM�������_ACT[������_DATA r���%L����xR�DISb�E�$�XVR�s���$�ZABC_GRPW 1t�Q�,#��0�2���ZIP�u'�&�����[MPCF_G 1v�Q�0�/�� w�ɤ� �	�Z/  8�5�/�/H/�/l$?� �+�/�/�/?�/�/??�?r?�?  � D0�?�?�?�?�?�;����x�]hYL�IND֑y� ���� ,(  *VOgM.�SO�OwO�O�M i?�O�O^PO 1_�OU_<_N_�_�O�_ �_�__�_�_x_-oo�Qo8o�_�o�oY&#29z� ���o C�e?a?>N|�oq�����qA�$DSPHERE 2{6M��_�;o���!� io|W�i��_��,�� Ï���Ώ@��/�v� ��e�؏��p�����������ZZ�� �N