��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  9�  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81F3�K2> �! � �$SOFT�T�_IDk2TOTAoL_EQs $�0�0NO�2U SPI�_INDE]�5X�k2SCREEN_�(4_2SIGE0�_?q;�0PK_F�I� 	$TH{KYGPANE�4� � DUMMYE1dDDd!OE4LA�!R�!R�	 � $TIT�!$I��N �Dd�DPd �Dc@�D5�F6�FU7�F8�F9�G0�G��GJA�E�GbA�E�G1B�G1�G �F�G2�B� SBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��4{V�a_EDIm   � �"���PS�`(4%$�EP�1�1$OP��0�2�a�p_OKv�UST1P_C� ुd��U �PLACI4!�Q�4�( ra�COMM� ,0$D����0�`��EOWB� BIGALLOW� (K�"(2�0VARa��@�2�aI�L�0OUy�C ,Kvay��PS�`��0M_O]�����CCFS_UT~p0 "�1�3�#��ؗ`X"�}R0  =4F IMCM�`O#�S�`��upi �_��p�B}�a���M�/ h�pIMPEE_F�N��N�`��@O��r�D_��~�n�Dy�F� dC�C_�r0  T0� '��'�DI�n0�"��p�P�C$I������F�t7 X� GRP0�z�M=qNFLI�<7��0UIRE��$�g"� SWITCH^5�AX_N�PSs"�CF_LIM�� � �0EED��!��qP�t�`P�J_dVЦMODE�h�.Z`�PӺ�ELBOF� �������p� ���3���� F@B/��0�>�G�� �� WARN	M�`/��qP��n�wNST� COR-�0bFLTRh�T�RAT�PT1�� $ACC1a��N ��>r$ORI�o"6V�RT�P_S� WCHG�0I��rQT2��1�I��T��I1��� x �i#�Q��HDR�BJ; CQ�2L�3�L�4L�5L�6L�7jL�8L�9{5CO`S <F +�=�O�x�#92��LLECy�}"MULTI�b@�"N��1�!���0T��w �STY�"�R`�=l�)2`��8��*�`T  |� �&$��۱m��P�̱��UTO���E��EXT����ÁB���"G2� (䈴![0������<�b+�� "D"���ŽQ��@<煰kc '�9�#���1��ÂM�ԽP���" '�3�$ �L� E���P<��`A�$JOBn�T����l�TRIG3�% dK�������<���\h��+�Y���_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`�0Z���0��P_�P��n@ ( @F RO.���&�t�IT�c�NOM�
����S���`T)w@���Z�1P�d���RA�0��p2b"����
$T��.��MD3�T��`QU31���p(5!HGb��T1�*E�7��c�KAb�WAb�cA4#Y�NT���PDBG�D�� *(��PU�t@X��W���AX���a��eTAI^cB�UF��0!+ g� 7n�PIW��*5 P�7M�8M�9
0�6F�7SIMsQS@>KEE�3PATn�^�a" 2`#��"�L64FIX!, ���!d��D�12Bus=CCI�:FgPCH�P:BAD렀aHCEhAOGhA]HW�_�0>�0_h@�f�Ak� ��F�q\'M`#�"�:DE3�- l�p3G@��@FSOES]FgH�BSU�IBS9WC��.� ` ��MARqG쀳��FACLp�SLEWxQ�e�ӿ��MC��/�\pSM_JB�M����QYC	g�e��Y�R�0 �n��CHN-�MP�G$G� Jg�_� <#��1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�fJR���rSEG�FR�PIO� S�TRT��N��cP!V5���!41�r�Ӏ
r>İ�b�B�O�2` +�[��� ,qE`j�,q`y�Ԣ}t8��yaSIZ%����t�vT�s� �z�y,qRSINF}Oбc����k��`��`�`Lp�ĸ T`7�CRCf�ԣCC/�9��`a�ua8h�ub'�MIN��uaPDs�#�G�D�YC��C�����e�q0��� ��EV�q�F�_
�eF��N3�s�ahƔ�Xa+p,5!�#=1�!VSCA?� �A��s1�"!3 ��`F/k��_�U��g�@�]��C�� a�s���}R�4� �ߠ��N����5a�R�HwANC��$LG��lP�f1$+@NDP�t�AR5@N^��a�q���c��ME�18����}0��RAө�AZ� 𨵰�%O��FCATK��s`"�S�P.FADIJ�OJ�ʠ �ʠ���<���Ր���GI�p�BMP��d�p�Dba��AESآ@	�K�W_��BA�S�� �G�5  �M�I�T�CSXh[@@�!62�	$X�K��T9�{sC���N�`�a~P_HEIsGHs1;�WID�06�aVT ACϰ��1A�Pl�<���EXqPg���|��CU�0_MMENU��7�TIT,AE�%�)�a2��a��8 YP� a�ED�E ��PDT��REM�.��AUTH_K�EY  ������ ��b�O	���}1E�RRLH� �9 \�� �q-�OR�DB�_�ID�@l �PUN_�O��Y�$SYSP0��4g�-�I�E��EV�#��(�PXW�O�� �: $SqK7!f2!DBTd�wTRL��; �'�AC�`��ĠIND&9DJ.D��_��f1���f���PL�AF�RWAj���SD�A���!+r|��UMgMY9d�F�10d�#AX(���J�<��}1�PR� 
3�PsOS��J�= �6�$V$�q�P�L~�>���SܠK�?�����CJ�@����EkNE�@T��A��|�S_�RECOR��_BH 5 O�@o=$LA�>$~�r2�R��`�q�b`�_�Du��0RO�@�aT [�Q��b������! <}У�PAUS���d�ETURN��MeRU�  CRp��EWM�b�AGNA9L:s2$LA��!?$PX�@3$P�y A �Abx�C0 #ܠDO�`�X�k�W�v�q�GO_oAWAY��MO�a�e�����CSS_�CCSCB C q�'N��CERI�� гJ`u�QA0�p}��@�GAG� R�0�`��{`��{`OF�q�5���#MA��X��i��LL�D� �$���sU�D)E�%!`���OVR1�0W�,�OR|�'��$ESC_$`�eD�SBIOQ��l ���B�VIB&� ��c,�����f�=pScSW���f!VL���PL���ARML	O
��`����d7%3SC �bALspH�MPCh �Ch �#(h �#h 5�UU��� C�'�C�'�#�$'�d��#C\4�$�pH��O`u��!Y��!�SB� ��`k$4�C�P3W���46$VOLTF37$$`�*�^1`��$`O1*�$o��0RQY��2b4�0?DH_THE����0SЯ4�7ALPH �4�`���7�@ �0�q*b7�rR�5�88 � ×���"��%Fn�MӁVHBPF�UAFLQ"D�s�`�THR��i2dB��(���G(��PVP���P��������1�J2�B0�E�C�E�CPSu�Y@ ��Fb3���H�(V�H :U�G�
X0��FkQw�[�Na�'B���C I�NHBcFILT ���$��W�2�T1� [ ��$���H mYАAF�sDO� �Y�Rp� fg�Q�+��c5h�Q�iSh�QP�L���Wqi�QTMOU�#c�i�Q\��X�g mb��vi�h�bAi�fI�aHIG��ca	x�O��ܰ��W�"vAaN-u!��	#AV�5H!Pa8$P�ד#p�R_:�A�a��B��N0�X�MC�N���f1[1�qVE �p��Z2;&f�I�QO��u�rx�wGldDN"{G|d��aF>!��9��aM:�U�FWA�:�Ml���X�Lu�@�$!����!l�ZO����0%O�lF�s�13�DI�W�@��Q����_��!CUR3VA԰0rCR41ͰZ�C<�r�H�v���<�``��<�(�f�CH�Q R3�S���t���Xp��VS_�`�ד�Fd��ژ���9&���NSTCY_ OE L����1�tP�1��U��24�2B��NI O7������DwEVI|� F���$5�RBTxS�PIB�P���BY�X����T��HN�DG��G H tn���L��Q��C���5��Lo0 aH��閻�FBP�{tFE{�5�t��T���I�DO���uPMCS�v>�f>�t�>"HOTSW�`s���ELE��J T���e�2��25�� O� ��HA7�E��3�44�0�Ғ���A�K ݬ� MDL� 2J~PE��	A��s ��tːÈ�s�JÆG! ��rD"�ó�����\�TO��W�	��/���SLAV�L  \0INPڐ���`�%ن_CFd�M�� $��ENU��OG��b�ϑ]զPƟ0`ҕ�]�ID�MA�Sa��\�WR0�#��"]�VE�$a�SKI�STs��sk$��2u���J��������	��Q���_SV>h�EXCLUMqJ2NM!ONL��D�Y���|�PE ղI_V>�APPLYZP���HID-@Y�r�_Mz�2��VRFY�0���r�1�cIOC_�f�� 1������O̥�u�LS���R$�DUMMY3�!����S� L_TP�/Bv�"���AӞ�ّ �N ���RTy_u�� չG&r[�O D��Pw_BA�`�3&x�!F ��_5����H������ �� �P $4 KwAR�GI��� q�2O{ �_SGNZ��Q �~P/�/PIG!Ns�l�$�^ sQ�ANNUN��@�T<�U/�ߴ�LAzp]	Z�d~���EFwPI�@ Rk @�F?IT�?	$TOTA%��Pd���!�M�NIY�S+���E��A[�
DAYS\�ADx�@��	�� �EFF_AX�I?�TI��0zCO�JA �ADJ_�RTRQ��Up���<P�1D �r5̀Ll�T�p? ]P�"�p��mtpd��V �0w�G���������SK�SU� ��CTRL_CA��� W�TRAN�S�6PIDLE_�PW���!��A�V曧V_�l�V ��DIAGS���X�� /$2�_SE�#TAC���t!`�!0z*@��RR��vPA���p ; SW�!�!�  ��ol��U��oOH��P�P� ��IR�r��BcRK'#��"A_Ak� ��x 2x�9ϐZs2��%l�W�pt*�x%oRQDW�%MSx��t5AX�'�"��LI�FECAL���10��N�1{"�5Z�3�{"dp5�ZU`}�MO�TN°Y$@FL9A�cZOVC@p�5�HE	��SUPP!OQ�ݑAq� Lj (CL�1_X6�IEYRJZRJWRJ�0TH�!UC|��6�XZ_AR�p6��Y2�HCOQ���Sf6AN��w$G���ICTE�Y }`��CACHE��C9�M�PLAN���UFFIQ@@�Ф0<�1	��6
��]�MSW�EZ 8>w KEYIM�p��TM~�SwQq�wQ�#���]�OCVIEܻ �[ A�BG�L��/�}�?� 	��?��D\p�ذST��!�R� �T� ��T� �T	��PEMA�If�ҁ��_F�AUL�]�RцĆ1�U�� �TR�E�^< �$Rc�uS�% IT��BUFW}�W��9N_� SUB~d���C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p�$��_~`�e�p%yOTT(����sP��M��Ot�T�LwAX � ��XX~`9#�c_G�3
ЧYN_1�_�D���1 �2M�*��T�F��H@ ~g�`� 0p���Gb-sC_R�AIAK���r�t�RoQ8�u7h�qDSPq��rP��A�IM�c6�\����s2�U�@�A�s�M*`IP���s�!DҐ6�TH�@n�)�OyT�!6�HSDI3��ABSC���@ V`y��� �_D�/CONVI�G��H�@3�~`F�!�pd��psqSCZ"���sgMERk��qFB��Lk��pET���aeR�FU:@DUr`����x�CD,���@p;cJHR�A!��bp�ՔՔ+PSԕCJN��C��p���ғSp�cH *�LX�:cd�Rqa�|  ����W��U��U���U�	�U�OQU�7R�8BR�9R��0T�^�1k�U1x�1��1��1��U1��1��1ƪ2Ԫ�2^�k�2x�2��2���2��2��2��2*ƪ3Ԫ3^�3k�x��3���o���3��3ʹ�3ƪ4Ԣ��EX9Tk!0�d <� 7h �p�6�pO��p����Na�FDRZ$eT^`V�Gr����䂴2�REM� Fj��BO�VM��A�TR�OV�DT�`-�MX<�IN��0,�W!'INDKЗ
w�׀�p$DG~q36���P�5�!D�6�RI�V���2�BGEAR��IO�%K�¾DN �p��J�82�PB@�CZ_MCM�@�1��r@U��1�f ,⑞�a? ���P\I�!?I�E�� Q�Q�am���g� _05Pfqg RI9ej��k!UP2_ h � �cTD�p���p! a���2F��wBAC�ri T�Ph�b�`�) OG���%���p��IFI��!�pm�>��	�PT��"��FMR2��j ��Ɛ+"�� ��\��������$�B`�x%��_ԡ�ޭ_����� M������D�GCLF�%DGDMY%LDa��5�6��ߺ4�@C��Uk�~�� T�FS#p�Tl P���e�qP>�p$EX_��B�1M2��2� 3��5��G ���m Y��Ѝ�SW�eOe6DEBUG���%�GR���pU�#BK�U_�O1'� �@PO�I5�65MS��OOfswSM��E�b�Q�0�0_E n �p|p �p�TERM�yo����ORI+���p��Y�S�M_���b�q�T�A�r�UP�Rs�� -�1�2n�$�' o$SEG�,*> ELTO���$USE�pNFIAU"4�e1���#$p$UFR���0ؐ0O!�0����OT�'��TAƀU�#NST��PAT��P�"P'THJ����E�P r�PV"ART�``%B`8�abU!REL:�aSHFT��V!�!�(_SH+@M$����� ��@N8r����OsVRq��rSHI%0���UN� �aAYLO����qIl����!8�@��@ERV]��1 �?:�¦'�2��%��5�%�RCq��EA�SYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba���
5Po��0�p6OR2�MY� `GR��t2b5n� � ��UP�a�Uu Ԭ")�.��TOCO!S�1POP ��`�pC��������Oѥ`REPR3��aO�P�b�"ePR�%WU.X1���e$PWR��I�MIU�2R_	S�$VcIS��#(AUD����Dv" v��$�H���P_ADDR
��H�G�"�Q�Q�Q�БR~pDp1�w H� SZ�a��e�ex�e��SE��r���HS��MNvx ���%Ŕ��OL���p<P��-��ACROlP_!QND_C��ג�1�T� �ROUPT��B_$�VpQ�A1Q�v� �c_��i���i��hx�`�i���i��v�ACk�IOU��D�gfsu<^d�y $|�P�_D��VB`bPR�M_�b3�ATT�P_אHaz (��OBJEr��P��[$��LE�#�s>`{ � ��u��AB_x�T~�S|�@�DBGLV���KRL�YHITC�OU�BGY LO: a�TEM��e�0>�+P'�,PSS|�P��JQUERY_F;LA�b�HW��\!�a|`u@�PU�b�PIO��"�]�ӂ�/dԁ=dԁ��S�IWOLN��}����CXa$SLZ�$INPUT_g�$IP#�P��'� &��SLvpa~��!� \�W�C-�B�0���p�F_ASv���$L ��w �F1G�U�B0m!���0�HY��ڑ��?�U;OPs� `�������[�ʔ[�і"�[PP �SIP�<�іI�2�x���IP_MEMBܿ�i`� X��IP�P�b{�_N�`�����R�����bS�P��p$FOCUwSBG;��UJ�Ə� �  � o7JsOG�'�DIS[�J7�cx�J8�7�� Im!�)�7_L�AB�!�@�A��A7PHIb�Q�]�D� J7J\���� �_KEYt� {�KՀLMONa=���$XR��ɀ~��WATCH_����3���EL��}Sy�~���s� f �!V8�g� �CTR3�쓥��LG�D� ��R��I�
LG_SIZ���J�q IƖ�I�FDT�IH�_�j V�GȴI�F�%SO��� q �Ɩ���v��ƴ�ǂK�S����w�k�N����E��\���'�*�U�s5��@�L>�4�DAUZ�E�A�pՀ�Dp�f�GH��B?�BOO���� C���PITp���� ��REC��OSCRN����D_p<�b�aMARGf�`���:���T�L���S��s��W�Ԣ�Iԭ�J{GMO�MNCH�c���FN��R�Kx�PRGv�UF��p0��FWD��HL��STP��V��+������RS��H�@�몖Cr4��?B��� +�O�U�q��*�a28��2��Gh�0PO���������M8�Ģ��EX.��TUIv�I��(�4�@�t�x�J0J�~�P��J0��N�a�#ANA��O"�0�VAIA��dCLE�AR�6DCS_H�I"�/c�O�O&�SI��S��IGN_�vpq�uᛀ�T�d� DEV-�L1LA �°BUW`Ո�x0T<$U�EM��Ł����0�A�R��x0�σ\�a�@OS1�2��3�a�`� �ࠜh�AN%-���-��IDX�DP�2MRO���Գ!�ST��R�q�Y{b! �$E&C+��p.&pA&`��a� L���ȟ%Pݘ��T\Q�UE�`�Ua��_ � �@(��`�b���# �MB_PN@ �R`r��R�w�TRIqN��P��BASS��a	6IRQ6�0�{MC(�� ���CLDP�� ETRQLI��!D�O9=4�FLʡh2�Aq3zD�q7��LDq5[4q5ORG�)�2�8P �R��4/c�4=b-4�t� �rp[4*�L4q5�S�@TO0Qt�0*D>2FRCLMC@D�?��?RIAt,1ID`�D�� d1��RQQp�rpDSTB
`� 1�F�HAXD2��|�G�LEXCES?R�`�BMhPa��@�BD4���B�q`�`�F_A�J�C[�Ot�H� K��� \��d�bTf$� ��LI�q��SREQUIRE��#MO�\�a�XDESBU��,1L� M�� �p���P�c��AA,1N��
Q�q�0/�&���-cDC��B�sIN�a?�RSM��Gh� N#B��N�aa�tcPST9� w� 4��LOC��RI���EX�fA�NG��AϠ��AQ䵗�@$��9�ZMF�����f��"��p�%u#ЖVSUP�%v+1FX�@IGGo�� �rq�"��1� �#B��$���p%#by���rx���vbPDATAK�pE;����Rr��M��*� t�`+MD�qI��)�v� ��t�A�wH�`��tD�IAE��sANSW���th���uD��)p�rԣ(@$`� PCU_�V6�ʠ�Aa&�PLOr�$`�R��&�Be���B�p������0 i�MRR}2�E�  ���V�A/A d$C'ALI�@��G~��2��!V��<$R��SW0^D"��A�BC�hD_J2SqE�Q�@�q_J3M�
G�1SP�,��@	PG�n�3m�u�3p�@���JkC���2'AO�)IMk@{BCSKAP^:ܔ9�wܔJy�{BQܜ�����`�_AZ.B��?�ELx��YAOCMP�c|A)��RT�j���c1�ﰈ��@1���t����Z��SMG��pԕ� ER!���:� �INҠACk�p��⁂�
n _�������D4�/R��DIU��C�DH�@
�#a�qc$V�Fc�$x�$���`@���b���� Rc�׀�H? �$BELP�����!ACCEL����kA°IRC_R��pG0�T!��$PS�@B2L$P ���W3�ط9� ٶPATH��.�γ.�3���p�A_��_��e�-B�`C���_M=G�$DD��ٰ��$FW�@�p�����γ����DE��P�PABN�ROTSPEEu��O0��DEF>Q��$P?$USE_��J%PQPC��JY����Z-A 6qYN�@A�pL�̐�L�MOU�3NG��|�OL�y�INCU��a�¢ĻBx��ӑ�AENCS����q�B�����D�IN��I�����pzC�V�E�����23_Ux ��b�LOWL�A��:�O0��0�Di�@�B�PҠ� ��PRC�����MOS� gTMO�pp�@-GPERCH[  M�OVӤ �� ���!3�yD!e�]��6�<�� ʓA����L IʓdWɗ��:p3�.��I�TRKӥ�AY ����?Q^���m�b��`pp�CQ�� MOM��B?R�0u��D���0y�0Â��DUҐZ��S_BCKLSH_C����o�n��T������
c��CLALJ��A��/PK�CHKO0�Su�RTY� �q��M�1r�q_
#c�_UMCPr�	C���SCL�n��LMTj�_L�0X����E�� � � ���m�h���L6��PC����H� ��P�ŞCN@�"XT\����CN_��N^CL�kCSF����V6Ҁ���ϡj���nCAT�SHs���� �ָ1���֙�������f��PA���_P���_P0� e���O1u��$xJG� P{#��OG���TORQU(�p�a�~����Ry������"_W��^���@��4t�
5z�
5I;I ;Iz�F�`�!��X_8�1��VC��0�D�B�21�>	P�?�B�5�JRK�<�2�6i�D�BL_SM�Q&BM�D`_DLt�&BGR�V4
Dt�
Dz��1H�_���31�8JCOSEKr�EHLN�0hK�5 oDt�jI��jI<1�J�L�Z1�5Zc@y��1MY�qA�HQBTHWMYT�HET09�NK2a3z�/Rn�r@CB4VkCBn�CqPASfa�YR<4gQt�gQ4VSB8t��R?UGTS���Cq��a��P#���Z�C$DUu ��R� �э2�Vӑ��Q�r�f'$NE�+pIs@�$|� �$R�#QA'UPepYg7EBHBALPHEE.b�.bS�E�c�E�c��E.b�F�c�j�FR�V�rhVghd��lV�jV��kV�kV�kV�kV
�kV�iHrh�f�r�m�!�x�kH�kH�kH��kH�kH�iOclORrhO��nO�jO�kUO�kO�kO�kO�kO�FF.bTQ���E���egSPBALAN�CE��RLE�PH_'USP衅F��F|��FPFULC�`3��3��E��1�l��UTO_p �%T13T2t���2NW�� ���ǡ��5�`�擊��T�OU���� I�NSEG��R�REqV��R���DIFH�f�1���F�1�;�COB��;C��2� ��b�4LCHWA�R��;�ABW!��$MECH]Q�@k�,q��AXk�P��8IgU�i�� 
���!ܭ���ROB��CR���ͥ*�C��_�s"T � x $WEIGHh�F9�$cc�� Ih��.�IF ќ�LAG�K�8SK��K�BI�L?�OD��U��S	TŰ�P�; ���(�������
�Ы�<L��  2�`�"�/DEBU.�L&�n�=�PMMY9��qNA#δ9�$D&�ƪ�$��� Q ]�DO_�A��� <	���~��LђBX�P�N��+�_�7�L�t�OH  �/� %��T�����T�����TICYK/�C�T1��%�Ä����N��c�Ã�R� L�S���S�����P�ROMPh�E� $IR� X�~ 8���!�MAI�0��4j���_9����tt�l�R�0COD��sFU`�+�ID_" �=�����G_SU;FF<0 3�O����DO��ِ�� R��Ǔن�S����!{�������	�H)�_F�I��9��ORDfX� ����36h��X�����GR9�S��ZDTD��v��ŧ4 *�L�_NA4���K��DEF_I[�K���g� ��_���i��Ɠ�š���IS`i �萚�D���e����4��0i�Dg����D�� O��LOCKEA!uӛϭϿ���{�u�UMz�K�{ԓ�{� ��{����}��v�� ���g������^�� ��K�Փ����!w�N�P'���^���,`��W\�[R�X ��TEFĨ ����OULOMB_tu�0�VISPWITY�A�!OY�A_FRId��(�#SI���R�������3���W�W���0��0_,�EAS%��!�& "����4p�G;� �h ��7ƵCOEFF_Om���$m�/�G!%�S.�߲�CA5����u�GR�` � � �$R� �X]�TM�E�$R�s�Z�/,)�E�R�T;�:䗰� M ]�LL��S�g_SV�($~◰��@���� �"SETU��MEA��Z�x0�u������� � � �� ȰID�"���!*�D�&P���*�F�'����)3��#����"�5;`*��R�EC���!7�SKy_��� P	�?1_USER��,���4���D�0��VEL@,2�0���2�5S�I���0�MTN�CFG>}1�  ���=Oy�NORE��3�l�2�0SI���� ��\�UX-�ܑP�DE�A $K�EY_����$gJOG<EנSVIA`�WC�� 1DSWy�x��
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���z�� �@_ERR���! ��S L�-���@���s0BB$BUF�-@X1_P�AMO�R�� H	�CU �A3�z�1Q�
��3���$��FVD��27ࡐbG��� � $SI�@ G�0VO B`נ�OBJE&�!FAD�JU�#EELAYh' ���SD�WOU��p�E1PY���=0Q�T i�0�W�DI�R$ba�pےʠD#YNբHeT�@���R�^�X����OP�WORK}1�,>�SYSBU@p 1�SOP�aR�!�jUĔk�PR��2�ePA`�0�!�cu� 1OP��EUJ��a'�D�Q/IMAG�A	��`fi�IMACrIN,��bsRGOVRD=a�b�0�aP�`sʠ�� �^uz�LP�B��@��!PMC_E(,�Q��N@�M�rǱb��1Ų7�=qSL&��~0���$OVSAL\G*E��*E2y�Ȑ�_=p�w��>p�s ���s	����y�tQ=q�#}1� @�@;���MOE�RI#A��
N���X�s�f�tQ��PL�}1�,RTv�m�AT�USRBTRC_T(qR��B �����$� �Ʊ��,�~0� D��`-CSALl`�SA0���]1gqXE���%���C��J�
���cUP(4����PX���؆�q��3�w� ��PG�5� $SUB�������t�JMPWAITXO��s��LOyCFt�!D=�CVF	ь�y�⻑R`�0��CC_�CTR�Q�	�IG�NR_PLt�DB�TBm�P��z�BW�)����0U@���IG��a��Iy�TNLND��Z�R]aK� N��B�0�PE�s���r���f�SPD}1� L�	�A�`gఠ�S��U!N�{���]�R!�B�DLY�2���+�7�PH_PK�E�~�2RETRIEt�`�2�bsR���FI�BǼ ����8� �2��0DBGLV~�LOGSIZ$C��KTؑUy#u�D�7�_�_T1@�EMB�@C\1A����R��|D�FCHECKK�P1���0����@&�f(bLEc�" PA9�QT���P�C߰PN�����ARh�0����Ӯ�PO�BORMATTnaF�f1h�`��2�S��UXy`�	�
�LB��4� � rEITCH���R{ 8PL)�AL_ � $���XPB�q� C,2Dx�!��+2�J3D���� T�pPDCK�yp��oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYL�OA��m�_1t�2<t���J3AR�����դ֏�laTIA4��5��6,2MOM�CP�����������0BϐAD��������PUBk`R��;����;���2���z4�` I$PI\Ds�o�@�1yՕ�w�2�w�Z��I��I��I���p� ���n���y�e`��9S)bT�SPEED� G��(�Е��/��� Е�`/�e�>��M�<�ЕSAMP�6V0��/���ЕMO�@ 2@�A��QP���C�� n�����������LRf`�kb�ІE9h�EIN 09��7S.В9
�yPy�GAMM�%S���D$GE�T)bP�cD]��2
��IB�q�I�G$HI(0;A��LR�EXPA8)LWVM8z)���g���C5�CHKhKp]�0�I_�� h`eT��n�q���eT,���� ��$�� 1�iPI>� RCH_D�313\��30LE�1�1\��o(Y�7 �t�MSW�FL �M��SCRc�7�@�&��%n�f�;SV���PB``�'�!�B�sS_SAaV&0ct5B3NO]�C\�C2^�0�mߗ� uٍa��u���u:e;��1���8��D�P��� ������)��b9� �e�GE�3��V�d�}Ml�� � ��YL��QNQS RlbfqXG�P�RR#@dCQp� �S:AW70��B�B[�CgR:AMxP�KCL�H���W�r��(1n�g�M�!o��� �F�P@}t$W P�u�P r��P5�R <�RC�R��%�6�`���� ��qsr X��O�D�qZ�Ug�ڐ>D�[ ��OM#w� J?\?n?�?�?��9�b"�۱��]�_��� | ��X0��bf��qf�� q`�ڏgzf��Eڐ��>j�"�ܰ��FdPnB��PM�QU��� � 8L�QCsOU!5�QTHI�sHOQBpHYSY�3ES��qUE�`�"��O���  �P��@\�UN���Crf�O�� P���Vu��!����OGR)AƁcB2�O�tVu�ITe �q:pINF�O�����{�qcB�v�OI�r� (�@SLEQS��q��p�vgqS���� =4L�ENABDRZ�PTIONt�����Q���)�GCF�ЎG�$J�q^r��� R���U�g�P�����_ED����ѓ �F��PK���E'NU߇وA�UT$1܅COPY������n�00MNx���PRUT8R� �Nx�OU���$G[rf�)�qRG�ADJ���*�X_:@բ$�����P��W��P��} ��)󂐶}�EX�YCDR�|�NS.��F@r�L�GO�#�NYQ_/FREQR�W� �#�h�TsLAe#���8�ӄ �CRE� sf�IF��sNA���%a�_Ge#ST�ATUI`e#MAIL�����q t��x�����ELEM��� �/0<�FEASI?�B��n�ڢ� 1�]� � I�p���Y!q]�t#A�AB$M���E�p<�VΡY��BASR�Z��S�U8Z��0$q���?RMS_TR;�q b ���SY�	�ǡ��$����>C�Q`	� 2� _�TM ������̲�@ �A��8)ǅ�i$DOU�s]$�Nj���PR+@3�֞�rGRID�qM�B7ARS �TY@���� O�p��� Hp_"}�!����d�O�P/��� � �p�`P�OR�s��}���SReV��)����DI&0T����� #�	�#�U4!�5!�6!�7!�I8��qF�2��Ep?$VALUt��%����b��/��� !;�1�q�����(F_�AN�#�ғ�Rɀ|(���TOTAL��,S��PW�Il��REGEN�1�c�X��ks(��a���`T1R��R��_S� ��1ଃV�����⹂Z�E��p�q��Vr���7V_H��DA�S�����S_Y,1�R4�S�� AR�P2� >^�IG_SE	s��d��å_Zp��C_��~��ENHANC�a�� T ;�8������INT�.���@FPsİ_OVRsP�`p�`��Lv�҂o��7�}��Z�@�SSLG�AA�~�2 5�	��D��S�BĤ�DE�U�����T�E�P���� !�Y��
�J��$2�IL_MC�x r#_��`TQ�`��q���'�B5V�C�P_� 0ڽM�	V1�
V1��2�2�3�3
�4�4�
�!���`� � m�A�2IN~VIBP���1�U2�2�3�3�4�4�A@-�C2�p� MC_YFp+0�0L	1(1d���M50Id�%"FE� S`�R/�@�KEEP_HNA�DD!!`$^�j)C�Q���$��"	��#O�a_$A�!�0�#i�.�#REM�"�$�P�½%�!�(U}�e�$�HPWD  �`#SBMSK|)G��qU2:�P	�COLLAB� �!K5��B�� ��g��pI�TI1{9p#>D� �,�@FLAP��$�SYN �<M�`C�6���UP_DL�YAA�ErDELAh�0ᐢY�`AD�Q�4BQSKIP=E�� ���XpOfPNTv�A�0P_Xp�rG �p�RU@,G��:I+�:I B1:IG�9JT�9Ja�9J�n�9J{�9J9<��R=A=s� X����4�%1�QB� NFL#IC�s�@J�U�H�LwNO_H�0�"?�֌RITu��@_P�A�pG�Q� ���^�U��W��LV�>d�NGRLT�0_q���O�  " ��OS��T�_JvA V	�APPR_WEIGH�s�J4CH?pvTOR8��vT��LOO��]�D+�tVJ�е�ғA�Q��U�S�XOB'�'�%�� �J2P���
7�X�T�<a43DP�=`Ԡ\"<a�q\!��RsDC��L� �рER��R�`� �RV�p�jr�b�RGE��8*��cN�FLG�a�Z����SPC�s�U�M_<`^2TH2�NH��P.a 1�� m`EF11��� lQ �!#� <�p3AT� g�S�� Vr�p�tMq�Lr���HOMEwr�t2'r�-?Qcu��w3'r���P����w4'r�'�@9�K�]�o����w5'r뤏��ȏڏ����w6'r�!�3�E�W�i�{��w7'r힟��Pԟ����w8'r��@-�?�Q�c�u��uS$0
�q�p�� sF��``S0p� `P����a�`/���-�IO[�M�I֠��qPOW=E�� ��0�Zatep�� y�5��$DSB OGNAL���0Cp�m�S2323�� Ɍ~`��� / ICEQP��PEp��5PsIT����OPBx0ޣ�FLOW�@TR`vP��!U���CU�M��UXT�A��w�ERFAC�� Uf��>0˰CH��'� tQ  _��>�f�Q$����OM���A�`T�P#UP%D7 A�ct�T��U�EX@�ȟ�U EFqA: X"�1RSPT�N����T ��PPaA�0o񩩕`EXP��IOS���)ԭ�_`���%��C�WR�A���ѩD�ag֕`ԦF�RIENDsaC2U�F7P����TOOLΫ�MYH C2LE�NGTH_VTE��I��Ӆ$S�E����UFINV�_���RGI��{QITI5B��X�v��-�G2-�G1@7�w�SG�X��_��UQQD=#���AS�Äd~C�`��q�� ��$$C/�S�`�����S0�0�����VERSI� ����0�5��I𼰲�����AAVM�_Y�2 �� 0  G�5��C�O�@�.r� r�	 ����S0����������������
?Q�Y�BS���1���� < -������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO`|O�O�O�OiCC�@OXLMT&����7  ��DIN�O�A\�Dq�EXE�HPV_��ATQz
���LARMRECOV �RgLMDG *��5�OLM_IF' *��`d�O�_ �_�_�_j�_'o9oKo<]onm, 
��o db��o�o�o�o^���$� z, A  � 2D{�PPIN�FO u[ @�Vw������� �`�������*� �&�`�J���n�����DQ����
��.� @�R�d�v����������a
PPLICATf��?�P��`�Handl�ingTool �
� 
V8.3�0P/40Cpɔ_LI
883���ɕ$ME
F�0G�4�-

�398�ɘ�%�z��
7DC3x�ɜ
�Noneɘ�Vr���ɞ@�6d� Vq_A�CTIVU��C\죴�MODPye��I��HGAPONp���OUP�;1*�� i�m�����Қ_����1�*�  �@���� ����Q���Կ濸@�
����� g���5�Hʵ�l�K�HTTHKY_��/�M�SϹ��� ������%�7ߑ�[� m�ߝߣߵ������� ���!�3��W�i�{� ������������� �/���S�e�w����� ����������+ �Oas���� ���'�K ]o������ ��/#/}/G/Y/k/ �/�/�/�/�/�/�/�/ ??y?C?U?g?�?�? �?�?�?�?�?�?	OO uO?OQOcO�O�O�O�O �O�O�O�O__q_;_ M___}_�_�_�_�_�_�_kŭ�TOp��
��DO_CLEAN�9��pcNM  !{衮o�o�o�o�o���DSPDRY�Rwo��HI��m@ �or����������&�8�J���MAXݐWdak�H�h��XWd�d���PL�UGGW�Xgd��P�RC)pB�`�k�aS�Oǂ2DtSEGF0�K� �+� �o�or����������%�LAPOb�x��  �2�D�V�h�z�����య¯ԯ�+�TOT�AL����+�USE+NUO�\� e�A��k­�RGDISPWMMC.���C6�&z�@@Dr\�OMpo��:�X�_STRI�NG 1	(�
��M!�S��
��_ITEM1Ƕ  n����� �+�=�O�a�sυϗ� �ϻ���������'��9�I/O S�IGNAL���Tryout M�odeȵInp�y�Simulat{eḏOut��OVERRLp� = 100˲In cycl��̱Prog A�bor��̱u�S�tatusʳ	H�eartbeat�ƷMH Fauyl	��Aler� L�:�L�^�p����8������ Scû Saտ��-�?�Q�c�u� ���������������);M_q��WOR.�û���� ��+=Oa s�������8//'.PO���� M �6/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?H"DEVP.�0d/�?O *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�J_\_n_PALT 	��Q�o_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o�_GRIm�û9q�_ as������ ���'�9�K�]�o� ������'�R	�݁ Q����)�;�M�_� q���������˟ݟ����%�7�I�ˏPREG�^����[����� ͯ߯���'�9�K� ]�o���������ɿۿ��O��$ARG_�� D ?	����0�� � 	$O�	+[D�]D��O�e��#�SBN_CON?FIG 
0˃����}�CII_SAVE  O������#�TCEL�LSETUP �0�%  OME�_IOO�O�%M�OV_H������R�EP��J��UTOoBACK�����FRA:\�o� Q�o���'�`��o��ҟ��= �� f�o������*�!�3�`�Ԉ��f�������� ��o�{��&�8�J�\� n�������������� ����"4FXj| �������끁  ��SYS�UIF.SV V� T.TP D }M9ATE.D�\�Tfx��c�INUI�Po���c�?MESSAG������8��ODE_D����z��O�0�c�oPAUSM!!�0�? ((O3�U/ g+Q/�/u/�/�/�/�/ �/�/�/)??M?;?q?�70$: TSK  �@-�ߠf�UPD�T��d�0
&XWZD_ENB����6STA�0��5�"�XIS��UNT� 20Ž� � 	�?gOJ�VO�OzO �O�O�O�O�O�O_1_n4DMET߀2CM�P_u__�_<YSCRDCFG 1�6_�Ь�����_�_oo(o:oLo��o�Q���_�o�o �o�o�o�o]o�o> Pbt���o9ǆi�GR<@�0/�sU�P_NA�/�	�i��v_ED�1��Y� 
 �%�-BCKEDTy-�'�GET@�AU�o�9��
�-(i�H�o�f�\�ּA��  ���2 �&�ȏE�D���~� ŏ׏m����3��&� �J�\�ߟJ�����9�ǟ�4���ϯ�\�����]�o�����5 N������\�w��)�;�ѿ_��6ϊ�g� ��\�CϮ���ϝ�+��7��V�3�z�\��@z�����i����8������]���F� �ߟ�5����9~������]����Y�k�����CR�!ߖ� ��W�q���#�5���Y���p$�NO_DEL���rGE_UNU�SE��tIGAL�LOW 1���(**TE�M*}S	$SERV_GR�}V� n: REG�$�}\� NUM�
���PMUB }U�LAYNP}\�PMPAL�COYC10#6 <$\ULSU��8:!�Lr�B�OXORI�CU�R_��PMC�NV�10|L�T4DLI�0��	����BN/`/ r/�/�/�/�/�/���p�LAL_OUT ��;���qWD_ABOR=f�q;0ITR_RTN�7y�o	;0NONS�0��6 
HCCFS�_UTIL �#<�5CC_@6A ;2#; h ?�?��?O#O�]CE_O�PTIOc8|qF@RIA_Ic Rf5Y@�2�0F�Q��=2q&}�A_�LIM�2.�k ��P��]B��K*}X�P
�P�2O�QK��B�r�qF�P�Q5T1)TR�H��_:JF_PARA�MGP 1�<g^&S�_�_�_�_�V�C�  C�d��`�o!o`�`�*`�`�Cd��Ti�i:a:e>eBa�GgC��`� D� D�	�`�w?��2H=E ONFI� E?n�aG_P�1#; ���o�1CUgy�aKP7AUS�1�yC ,������ ���	�C�-�g�Q� w���������я���r�O�A�O�H�L_LECT_�B�IPV6�EN. QF�3��NDE>� �G��71234567890��sB�pTR����%
 H�/%)�������W� ��0�B���f�x���� ����ү+�����s� >�P�b���������� ο��K��(�:ϓ��^�|��B!F� |�I|�IO #��<U%e6�'�9�K߶��TR�P2$��(`9X�t�Y޼`%��x�ڥH��_MOR�3&�=��i��A� $��H�6�l�Z���~S"��'�=�r_A?�a�a�`��@K��R�dP�)F�ha�- �_�'�9�%
�k���G� ��%Z�%���`�@c.�PD�B��+���cpmidbg��	�`&:�����p��N>  ��@��b.���]ܭ@as<�^��@�sg�$��f�l�q��ud�1:��:J��DE�F *ۈ��)��c�buf.t�xt����_L�64FIX , ������l/[Y/�/}/ �/�/�/�/
?�/.?@? ?d?v?U?�?�?�?�?��?�?,/>#_E -���<2ODOVOhOXzO�O6&IM��.o�=YU>���d�
�6IMC��2/���ñdU�C��20�M��QT:Uw�Cz  B �i�Ol_W_�_{_�_��_�D��22o�DT|����� ����C�C����2
�xObi�D4cdv`�D��`/�`v`�]E��D D�` E�4�F*� E�c��FC���[F����E��fE���fFކ3FY�F�P3w��?��@�33 ;?��>L���Aw��n,a@��@e�5!و��a���`A��w�=�`<#�*
Ѫ_��ozJRSMOFST (�,bI+T1��D @3��
�c��'�a��;��b�w?���<��M�NTESTR�1O�CR@�4�4�>VC5`A�w�Ia�+a�aORI`CTPB͖U�C�`4����r��:d�*�qIj?�5��qT_�?PROG ��
��%$/ˏ�t��NUSER  k��������KEY_TBL'  ����#a��	
��� !"�#$%&'()*�+,-./��:;�<=>?@ABC��GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?�����������LCK�
����S�TAT/��s_AU�TO_DO ��	�c�INDT_ENBP���Rpqn�`�sT2����STOr`쓯�XC�� 26��) 8
SONY XC-56��"b����@��F(� А�H�R50w���>�P�7<b�t�Aff����ֿ� Ŀ����C� U�0�yϋ�fϯ��Ϝ���������-ߜ�TR�L��LETEͦ ���T_SCRE�EN ���kcs���U�MMENU 17�� <ܹ���w� ��������K�"� 4��X�j������ ������5���k�B� T�z������������� ��.g>P� t������ Q(:�^p� ���/��;// $/J/�/Z/l/�/�/�/ �/�/�/�/7?? ?m? D?V?�?z?�?�?�?�? �?!O�?
OWO.O@OfO��OvO�O�O(y��RE�G 8�y�����`�M�ߎ�_MAN�UAL�k�DBC�O��RIGY�9�DBG_ERRL��9�ۉq��_�_��_ ^QNUML�I�pϡ�pd
�
�^QPXWORK 1:���_5oGoYo�ko}oӍDBTB_NN� ;������ADB_A�WAYfS�qGC�P 
�=�p�f_A!L�pR��bbRY�[�t
�WX_�P 1<{y�n�,�%oc�Pl��h_M��ISO���k@L��sONTImMX��
���v�y
��2sMOTN�END�1tREC�ORD 1B��� ���sG�O� ]�K��{�b�������� V�Ǐ�]����6�H� Z���������#�؟ ������2���V�ş z��������ԯC��� g��.�@�R���v�� ��	���п���c�� ��#ϫ�`�rτϖ�� ��)ϳ�M���&�8� ��\�G�Uߒ�߶��߀��I������4��  �p7�n���ߤ��� ������"���F�1� ��|��������[��� ��i���BTf����bTOLERE�NC�dB�'r�`L���^PCSS_CCSCB 3C>y�`IP�t}�~� <�_`r�K������/�{� �5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O��O_�~�LL� D���&qET�c�ao C[C��P�ZP^r_ A� p� �sp��QGPt[	 A�p�Q�_�[A? �_�[oU�pc�P�pSB�V �c�(a�PWoio{h+
�o�h�o�oY���[	r�hLU��NQ]�7�n�2G#�2ܘ߈�c��aD�@VB��|�G����+��K� �otGhXGrcso����e�B   =���2�a>�tYB�� �pQC�p�q�aA"�H�S �Q-��q���ud�v������AfP ` 0����D^P��p@5�a
_�XTHQH����a aW>� �a9P��b�e:�L�^� h�Hc�́PQ�RFQ �PU�z�֟�o\^� �-�?��c�u���zCz�ů�b2x�Щ�RD��m��m�%����S̡0� �]�0�.��@���EQ�p��F�X�ѿUҁ�п�VSȺNST�CY 1E��]�ڿ��K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߒ���DEVICE ;1F5� MZ�� �a��	� ��?�6�c���	{䰟���_HNDGD G5��VP���R�LS 2H�ݠ��/�A�S�e��w����� ZPARA�M I�FgHe~�RBT 2K�܋8р<��WPpCU�C��,`¢P�Z��z�����C*  �2�jMTLU,`"nPB, s� �M� }�gT�g��
#B��!�bcy� [2Dchz�����/��/gT#�I%D��C�` �b!�R��A��A�,��Bd��A5��P��_C4kP�!�2�C��$Ɓ�]�f�fA�À��B�� �| ���/�/�T (��54a5�} %/7/d?/M?_?q? �?�?�?�?�?O�?O O%O7OIO�OmOO�O �O�O�O�O�O�OJ_!_ 3_�_�_3�_�_�_�_ �_o�_(ooLo^oЁ =?k_IoS_�o�o�o�o �o�o�o#5G �k}����� ��H��1�~�U�g� y�ƏAo�Տ���2� D�/�h�S���go���� ԟ����ϟ���R� )�;���_�q������� ���ݯ�<��%�7� I�[�m��������� }�&��J�5�n�Yϒ� �Ϗ��ϣ�ѿ���� ��F��/�Aߎ�e�w� �ߛ߭���������B� �+�x�O�a���� ��������,���%�b� M���q����������� ����L#5� Yk}��� � �61CUg �������� 	//h/���/w/�/�/ �/�/�/
?�/.?@? I/[/1/_?q?�?�?�? �?�?�?�?OO%OrO IO[O�OO�O�O�O�O �O&_�O_\_3_E_W_ �_?�_�_�_�_�_"o oFo1ojoE?s_�_�o m_�o�o�o�o�o0 f=Oa��� �������b� 9�K���o���Ώ��[o ��(��L�7�I����m������$DCS�S_SLAVE �L���ё���_4D�  љ��CFoG Mѕ��������FR�A:\ĐL-�%0�4d.CSV�� � }�� ���A Vi�CHq�z����p��|�����  ������Ρޯ̩ˡҐ-矩*����_CR�C_OUT N�������_FS�I ?њ ����k�}����� ��ſ׿ �����H� C�U�gϐϋϝϯ��� ������ ��-�?�h� c�u߇߽߰߫����� ����@�;�M�_�� ������������� �%�7�`�[�m���� ������������8 3EW�{��� ���/X Sew����� ��/0/+/=/O/x/ s/�/�/�/�/�/�/? ??'?P?K?]?o?�? �?�?�?�?�?�?�?(O #O5OGOpOkO}O�O�O �O�O�O _�O__H_ C_U_g_�_�_�_�_�_ �_�_�_ oo-o?oho couo�o�o�o�o�o�o �o@;M_� �������� �%�7�`�[�m���� ����Ǐ������8� 3�E�W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿� ��'�P�K�]�oϘ� �ϥϷ���������(� #�5�G�p�k�}ߏ߸� ������ �����H� C�U�g������� ������ ��-�?�h� c�u������������� ��@;M_� ������� %7`[m� ������/8/ 3/E/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO�sO�O�O�O�O�C�$�DCS_C_FS�O ?�����A P �O�O_?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo ~o�o�o�o�o�o�o�o 72DVz� ������
�� .�W�R�d�v������� ������/�*�<� N�w�r���������̟ ޟ���&�O�J�\� n���������߯گ� ��'�"�4�F�o�j�|� ������Ŀֿ�������G�B�T��OC_RPI�N_jϳ��� �ς��O����1�Z�U��NSL��@&�h߱� ��������"��/�A� j�e�w������� ������B�=�O�a� ���������������� '9b]o� ������� :5GY�}�� ����///1/ Z/U/g/y/�/�/�/�/ �/�/�/	?2?-???Q? z?u?��ߤ߆?�?�? �?OO@O;OMO_O�O �O�O�O�O�O�O�O_ _%_7_`_[_m__�_ �_�_�_�_�_�_o8o 3oEoWo�o{o�o�o�o �o�o�o/X Sew����� ���0�+�=�O�x� s���������͏ߏ� ��'�P�K�]�o������ �PRE_CH�K P۫�A ~��,8�2x��� 	 8�9�K���+�q���a� ������ݯ�ͯ�%� �I�[�9����o��� ǿ��׿���)�3�E� �i�{�YϟϱϏ��� ��������-�S�1� c߉�g�y߿��߯��� �!�+�=���a�s�Q� ����������� ���K�]�;�����q� ������������#5 �Ak{�� ����CU 3y�i���� ��/-/G/c/u/ S/�/�/�/�/�/�/? ?�/;?M?+?q?�?a? �?�?�?�?�?�?�?%O ?/Q/[OmOO�O�O�O �O�O�O�O_�O3_E_ #_U_{_Y_�_�_�_�_ �_�_�_o/ooSoeo GO�o�o=o�o�o�o�o �o=-s� c������� '��K�]�woi���5� ��ɏ��������5� G�%�k�}�[������� ן�ǟ����C�U� o�A�����{���ӯ�� ��	��-�?��c�u� S�������Ͽ῿�� ���'�M�+�=σϕ� w�����m������%� 7��[�m�K�}ߣ߁� ���߷����!���E� W�5�{��ϱ���e� ������	�/��?�e� C�U������������� ��=O-s� ���]���� '9]oM�� �����/�5/ G/%/k/}/[/�/�/� �/�/�/�/?1??U? g?E?�?�?{?�?�?�? �?	O�?O?OOOOuO SOeO�O�O�/�O�O�O _)__M___=_�_�_ s_�_�_�_�_o�_�_ 7oIo'omoo]o�o�o �O�o�o�o!�o1 W5g�k}�� ����/�A��e� w�U�������я��o ����	�O�a�?��� ��u���͟����� '�9��]�o�M����� ����ۯ��ǯ�#�ů G�Y�7�}���m���ſ �����ٿ�1��A� g�E�wϝ�{ύ����� ��	�߽�?�Q�/�u� ��e߽߫ߛ������� �)���_�q�O�� ������������ 7�I���Y��]����� ����������!3 WiG��}�� ��%�A�1 w�g����� �/+/	/O/a/?/�/ �/u/�/�/�/�/? �/9?K?�/o?�?_?�? �?�?�?�?�?O#OO GOYO7OiO�OmO�O�O �O�O�O_�O1_C_%? g_y__�_�_�_�_�_ �_�_o�_+oQo/oAo �o�owo�o�o�o�o �o);U__q� �������%� �I�[�9����o��� Ǐ�����ۏ!�3�M ?�i��Y�������՟ �ş����A�S�1� w���g�����������ӯ�+�=��$DC�S_SGN Q�K�c��7m� �14-JAN�-19 08:3O8   O�l� ����� N.D�Ѥ���������h��x,rWf*σ��^M��  O�V�ERSION �[�V3.5�.13�EFLO�GIC 1RK���  	���P�?�P�N�!��PROG_ENB  ��6Ù�o�ULSE  T����!�_ACCL{IM���������WRSTJN�T��c��K�EM�Ox̘��� ���INIT S.�G�Z����OPT_SL �?	,��
 	�R575��Y�7�4^�6_�7_�50
��1��2_�@ȭ��><�TO  Hݷ�t��V�DEX���dc����PAT�H A[�A\��g�y��HCP_�CLNTID ?<��6� @ȸ�����IAG_GR�P 2XK�? ,`��� � �9�$�]�H������123456�7890����S�� |�������!�� ��H���;� dC�S���6� ����.�R v�f��H� �//�</N/�"/ p/�/t/�/�/V/h/�/ ?&??J?\?�/l?B? �?�?�?�?�?v?O�? 4OFO$OjO|OOE� �Oy��O�O_�O2_��@_T_y_d_�_,
�B^ 4�_�_~_`Oo �O&oLo^oI��Tjo�o .o�o�o�o�o �O' �_K6H�l�� �����#��G� 2�k�V���B]���Ǐ ُ�������(��L� ^�p�;������������ٟ���CT_C�ONFIG Y���Ӛ�e�gU���STBF_TTS��
��b����Û�u�O�MAU���|��MSW_CuF6�Z��  伿OCVIEW��[ɭ������-� ?�Q�c�u�G�	����� ¿Կ������.�@� R�d�v�ϚϬϾ��� ����ߕ�*�<�N�`� r߄�ߨߺ������� ��&�8�J�\�n�� ��!����������� ��4�F�X�j�|����KRC£\�e��!*� B^������C2�g{�SBL_FA?ULT ]��ި>�GPMSKk���*�TDIAG �^:�աI���UD1: 6789012345�G�BSP�-?Q cu��������//)/;/M/� �
@q��/$��TRECP��

 ��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOi/{/�xO�/UMP_OP�TIONk���AT�R¢l��	�EPM�Ej��OY_TEM�P  È�33B�J�P�AP�D�UNI��m�Q��Y�N_BRK _�ɩ�EMGDI_�STA"U�aQSUN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 I�#X��,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;���m��څ �!�� ��~�ߢ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$
T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����裆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7����; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  D�B���ȕ?\�?&}�B�?�1�3�ٸ*9�N SMTT#t�[)��X}�C�f�HoOSTCd1ux�o��� 	zHMzKzOx��O�Ie�O�O	__-_ ;Z�O^_p_�_�_�O�_�KP	anonymous�_�_�_oo1o yO�O�Ozo�_�O M_�o�o�o�o?_. @Rd�o�_�_�� ���;oMo_oqos `��o��������̏ ����&�8�[��� ��������ȟ�!�3� �G�4�{�X�j�|��� Տ��į֯����� e�B�T�f�x���џ� ���	��=��,�>� P�bϩ��ϘϪϼ��� �'�9��(�:�L�^� ����ɿw��������  ��$�6���Z�l�~� ��ߴ����������  �g�yߋߝ�z����� ����������?�. @Rd������� ���;�M�_�q�s `������� �//&/I7/�n/��/�/�/�/#O\AEN�T 1v
; P�!J/?  � �/3?"?W??{?>?�? b?�?�?�?�?�?O�? AOOeO(O�OLO^O�O �O�O�O_�O+_�O _ a_$_�_H_�_l_�_�_ �_o�_'o�_Koooo 2o{oVo�o�o�o�o�o �o5�oY.��R�v��zQUICC0���3���t14��"����t2���`�r�ӏ!ROUTERԏ��#�!PCJOG$����!192.�168.0.10���sCAMPRT,t�P�!d�1m�����RT폟�����$NAME !�*?!ROBO����S_CFG 1u��) ��Auto-sta�rtedFTP&��=?/֯s ����0�B��f�x� ��������S����� �,���������ϼ� ޯ���������ʿ'� 9�K�]�oߒ�ߥ߷� ��������(: ~�k�Ϗ������� ������1�C�f��� y������������,� >�R�?��cu� �`�����( �$M_q���� �� /H%/7/ I/[/m/4�/�/�/�/ �/�~/?!?3?E?W? i?����?�/�?/ �?OO/O�/�?eOwO �O�O�?�ORO�O�O_ _+_r?�?�?�?�O|_ �?�_�_�_�_o�O'o 9oKo]ooo�_o�o�o �o�o�o�oF_X_j_ ~ok�_����� �o���1�TU���y���������U�)�_?ERR w3�я��PDUSIZ � g�^�p����>�WRD ?�r�Cq�  ?guestb�Q��c�u�������"�SC�DMNGRP 2�xr�����Cqg�\�b�K� �	P01.00� 8(q   e�5p�5pz�5p�B  �{ ����H����L��L��L�����O8�����l������a4� x��Ȥ�Zx��8���\����)�`�;�������d�.�@�R��ɛ_GROUېy*�����	ӑ����QUPD  d?u����İTYg�����TTP_AUTH 1z��� <!iPeOndan��-�l����!KARE�L:*-�6�H�K�C]�m��U�VI�SION SET ���ϴ�g�G�U����� �R�0��H�Bߏ�f��x��ߜ߮���CTRL {����g��
g�FFF9�E3��AtFRS�:DEFAULT�;�FANUC� Web Server;�)���9�K� �ܭ���������߄�WR_CONFI�G |ߛ �;��IDL_CP�U_PCZ�g�B��Dpy� BH_�M�INj�)�}�GNR_IO��g���a��NPT_SIM_�D_�����STA�L_SCRN�� ����TPMODN�TOL������RT�Y��y���� �EN�O���Ѳ]�OLN/K 1}��M���������eM�ASTE��ɾeSLAVE ~��|c�O_CFG�ٱBUO�O@C�YCLEn>T�_?ASG 1ߗ+�
 ����/ /+/=/O/a/s/�/�/p�/�/��NUM���
@IPCH��^RTRY_CNZ���@��������� @kI��+E�z?E�a�P_�MEMBERS �2�ߙ� $���2���ݰ7�?�9a��SDT_ISOL�C  ����$�J23_DSM�+�3JOBPRO�CN��JOG��1�+�d8��?��+�O�/?
�LQ�O__/_@�OS_e_w_�_`�O� Hm@��E#?&BPO�SREQO��KANJI_���a[�?MON ����b�yN_goyo�o�o�oH�Y�`3�<� ��e�_ִ��_L���"?�`EYLOGGI�NLE��������$LANGUA�GE ��<�T� {q�LGa2��	�b���g�xP��W  ��g��'��b���>��MC:\RSCH�\00\<�XpN_DISP �+�G�J��O�O߃LOClp�Dz���As�OGBOOK ������󑧱����X�����Ϗ�����a�*��	 p�����!�m��!����=p_BUFF 1-�p��2F幟����՟D� Co�llaborativǖ���F�=�O� a�s�������֯ͯ߯����B�9�K���D�CS �z� =���'�f��?ɿۿ����H@{�IO 1�� ~?9ü��9�I�[�mρϑϣ� �����������!�3� E�Y�i�{ߍߡ߱���h�����E��TMNd�_B�T�f�x��� ������������,� >�P�b�t�������L�N�SEVD0��TYPN1�$6���QRS"0&��><2FL 1�"�J0��������GTP:pO}F�NGNAM1D��mr�tUPS�G�I"5�aO5�_L�OADN@G %��%DF_MO�TN�y�� MAXUALRM�'���(���_PR"4F0�d��1�B_PNP�� V 2�C	�MDR0771�ߕ�BL"806=3%�@ �_#?�hߒ|/�C��z��6��/���/Po@P �2��+ �ɖ	�T 	t  ��/�%W?B?{?� k?�?g?�?�?�?O�? *OONO`OCO�OoO�O �O�O�O�O_�O&_8_ _\_G_�_�_u_�_�_ �_�_�_o�_4ooXo joMo�oyo�o�o�o�o �o�o0B%fQ �u������ ��>�)�b�M����� {��������Տ�� :�%�^�p�S��������D_LDXDI�SApB�MEM�O_APjE ?=C
 �,� (�:�L�^�p�������ISC 1�C ����4�����૟4��X���C_M?STR ���w��SCD 1��� L�ƿH��տ���2� �/�h�Sό�wϰϛ� �Ͽ���
���.��R� =�v�aߚ߅ߗ��߻� ������<�'�L�r� ]���������� ����8�#�\�G���k� ��������������" F1jUg�� �����B -fQ�u����h�MKCFG 񓆽�/�#LTAR�M_��7"�0�0N/V$� MEgTPUᐒ3�����ND� ADCOLxp%� {.CMNT�/s �%� �����.E#>!�/4�%PO�SCF�'�.PR�PM�/9ST� 1���� 4@��<#�
1�5�?�7 {?�?�?�?�?�?�?)O OO_OAOSO�OwO�O��O�O�O_�A�!SI�NG_CHK  ��/$MODAQ�,#����.;UDE�V 	��	M�C:o\HSIZE�ᝢ��;UTASK� %��%$12�3456789 ��_�U9WTRIG +1���l3%%��9o���"ocoFo5#�VYP�QNe��:SEM_�INF 1�3'� `)�AT&FV0E0�po�m)�aE0V�1&A3&B1&�D2&S0&C1�S0=�m)ATZ�o;"tH?g�a[o�xA��z���� �o>��o '��K������ ��я:�L�3�p�#� 5���Y�k�}������ $�[�H���~�9��� ��Ưد��������ӟ �V�	�z�������c� Կ����
��.��� d��)�;��Ͼ�q��� ����˿<���`�G� �ߖ�IϺ�m�ϑϣ� ���8�J��n�!ߒ��M�������h_NIwTOR� G ?�[�   	EX�EC1�/�25�3�5�45�55��P7�7*5�85�9�0�� ��4��@��L��X� ��d��p��|�������2��2��2���2��2��2��2���2��223ʡ�3��3@�;QR_�GRP_SV 1��k (��7U��Q_D��^�PL�_NAME !�3%,�!De�fault Pe�rsonalit�y (from �FD) �RR2�� 1�L6(�L?�,0	l d������ ��//(/:/L/^/ p/�/�/�/�/�/�/�/ZX2u?0?B?T?f?@x?�?�?�?�?\R<? �?�?O O2ODOVOhO�zO�O�O�OZZ`\R�?�N
�O_\TP�O:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHo_)_~o�o�o�o �o�o�o�o 2D Vhz�[omo�� ��
��.�@�R�d��v���������Џ�� Ef  Fb�� F7���Q��!��d�?� Q�6�t�������pş���� ݘ ����"�@�F�d����ܐ"𩯹�ݐA�#  ϩU[�$n��B�E ��� � @D7�  �?�� ��?�@��A@�;f���FH� ;�	l>,�	 |��j�ys�d�>���� ��ܐK(��K�d$2K ��J�7w�KYJ˷�ϜJ�	�ܿ��ܐ@I���_�f�@�z���f�γ�N��}����	Xl��������S��ĽÔ��X������5���  �����A?oi#��;��A��� o���l� �π��-���ܛG�G�ܒ���@n�@a �  �  ���ܟ*�͵	'�� � H�I� �  �Р�n�:�Èl�È�=��̈́��@�ߚЕ����/������̷NP� � ',���-�@�
�@���?�=�@A���B� � Cj�a�Be�Czi��@#�B�~��������bbdʷB Р��P����̠�����ADz՟�n�3�� C�i�@�R�R�Yщ���  �@� �  ��?�faf������n� ɠ #U�y9G
(���I�(�@uP~�����t�t���>����;��Cd;��.<�߈<�g�<F+<L��������,�d�,�̠?ff�f?��?&&��@���@x��@��N�@���@T�H�ِ�!-� ȹ�|��
`��� ����//</'/�`/r/]/�/��eF ���/�/�/�/m?���/J?�(E��G��#�� FY�T?�? P?�?�?�?�?�?O�? /OO?OeOPD�O�I QOG�?�O1?�OmO_0_B_T_������A_�_	_�_�_�_ o
��A��An0 bФ/o� C�_Uo�_�Op�Ƀ؃o�o�o�o���mW�����oC�E� q�H�d���؜a@q��e�F�B���WB]�NB2��(A��@��u\?�D������������b�0�|�uR����
x~��ؽ��B�u*C��$��)`�$ ����GC#����rAU�����1�eG�D�I��mH�� I�:�I�6[Fߍ��C�I���J�:\IT��H
~QF��y��p�*J��/ I8Y�I���KFjʻC e�o��s�����Џ�� �ߏ�*��N�9�r� ]������������۟ ���8�#�\�G����� }�����گů���"� ��X�C�|�g����� Ŀ�������	�B� -�f�Qϊ�uχ��ϫ� �������,��P�b� M߆�qߪߕ��߹��� ����(��L�7�p�[��������s(����3:���9�$���3���d�,�4��@�R�wa�����l�~�wa����e����wa4 �{������((L:ueP�P~�A�O������	����G 2W}h���� ��/���O�O7/m/[(d=�s/U/�/�/ �/�/�/?�/1??U?�C?y?�=  2 �Ef9gFb��77��9fB)aa)`C9A`�&`w`@-o�?O@O(O:OLO]M{c�?@�?�O�O�O�O9c?�0T�A7h$w`w`�!w`xn
  �O9_K_]_o_�_�_�_ �_�_�_�_�_o#ozz�Q ��h��G����$MR_CA�BLE 2�hO �a�T� @@�0�Ae��a�a��a��`��0�`C<�`�aO8�t/o�l��o�f�#��0�<�0�DO��h?���o�h8  ���Cu�07�d4
H.�d�`y`By`9C�p�bHE�^p��dҠ`��0�q�p�b0�����c -���H� �2���V��� ��������'�"���LD���CH�Do<� \���������������*,�** �\cOM �ii�����r��%�% 234567O8901i�{� f�H����������1�����
��`��not sent� 5���;��TESTFECS�ALGR  eg�`��1d.�š
:�� �DCbS�Q�c��u��� 9UD1�:\mainte�nances.xsml��ֿ  Z��DEFAU�LT�mi4\bGRPw 2�M�  =���7�E  �%F�orce�sor� check  �����z��p����h5-��ϻ���������%!1st c�leaning �of cont.� v�ilatiCon��}�Rߗ+��@[�ߔߦ߸����mech�cal,`������0��h5k�@�R�d�v������(�rolle _Ƶ����/����(�:�L��Ba�sic quarterly��������,����������F�M��:(�"GpBP(�X_h5��@�����#C���M"��{Pb�t���Sup�pq�grease���?/&/�8/J/\/��C+ ge���. batn�y`/��/h5	/�/�/��/? ?_�ѷenB'�v��/�/��/����?�?�?�?�?�GX=?O(�Dp"CrB1O��0�/`OrO�O�O`�O�t$��Lf��C!-(��A�O:�OO$_�6_H_Z_l_�t*cgabl�O(���S!<(��Q�_:�
_�_ �_oo0oo)(Ӂ/�_�_���_�o�o�o�o��o�O@haul1�l�2r x(�<qC:��op�������Repla�W�fUȼ2�:�.�_4�F�X�j�|�(�$ %���ߟ����#���
� �.�@���d���ŏ׏ ����П����U�*� y�����r��������� 	�q��?�߯c�8�J� \�n���ϯ�����ڿ )����"�4�Fϕ�j� ��˿����������� �[�0�ϑ�fߵϊ� �߮�����!���E�W� ,�{�P�b�t����� ������A��(�:� L�^���������� ���� $s�H�� ����q����� 9]o�Vhz ���U�#�G /./@/R/d/��/�/ ��//�/�/??*? y/N?�/�/�?�/�?�? �?�?�???Oc?u?JO �?nO�O�O�O�O+Jkb	 H�O�O__6M 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<ND@� �bA?�  @!Q _����Fw�� �H;* �** @A>F �pRT�f�x�:�������ҏ��eO^C7� Տ#�5�G�	�k�}��� ُ���c�����W� �C�U�g���ß)��� ��ӯ���	��-�w� ����9�������m�Ͽ���=�O�E!Q��$MR_HIST� 2�>EN�� �
 \
B$ 23�45678901P^�f�#��]�9O ���φϸ�O�)�;� ���q߃ߕ�L�^߬� ���ߦ����7�I� � m�$���Z���~��� ���!���E�W��{��2�����h�����:�S�KCFMAP  ]>EQ��r�5�!P����ON�REL  .��3���EXCFENB8
��Q�FNCXJJOG_OVLIM8dN�\� ��KEY8�=�_PAN7�\���RUN�����SFSPDT�YPxC��SIG�N8JT1MOT��G��_CE_�GRP 1�>EV��@���� �/Ⱥ��/�/ U//y/0/n/�/f/�/ �/�/	?�/???�/c? ?\?�?P?�?�?�?�?��?O)OOMO,���Q?Z_EDIT5 �)TCOM_CF/G 1���[�O�O�O 
�ASI �y3�
__B+[_O_��>O��_bHT_ARC_�U.Ń	T_MN�_MODE5���	UAP_CPL��_gNOCHEC�K ?�� �� o.o@oRodo vo�o�o�o�o�o�o�o�*!NO_WAIT_L4~GiNT�A���EUw�T_ERRs2���3��ƱJ���b��>_)��|MO�sű�}x:Ov���8�?����� |l��rPARAM�r����lTh��p9I5�5�G� = �� d�v�~�X�������������֟�0��e���b�t�����SUM_RSPACE������Aѯۤ�$OD�RDSP�S7cO�FFSET_CAqRt@�_�DIS���PEN_FIL�E:�7�AF�PT?ION_IO���q�M_PRG %��%$*����M�WORK �y=f ��춍�D�� �����	 ������gT���RG_DSBOL  ��C�{�u��RIENTT5O7 �C� �A �UT_SIM_Dy����V�LCT ���}{B �٭��_PEqX�P=��RAT�W� dc��UP� ���`���`e�w�]ߛߩ��$��2r�L6(L�?���	l d������&�8�J� \�n��������� �����"�4�F�X���2�߈����������� ��*�<w�T fx������p�J`[�ˣG���Tz��P g������/ "/4/F/X/j/|/�/�/ �/���/�/??0? B?T?f?x?�?�?�?�? �?�?�?�/�/,O>OPO bOtO�O�O�O�O�O�O �O__(_:_��Oe�C�y_�]2ӆ��_ �^�_�_�W^]^]��/ooSog�Hgroho zo�o�o�o�o�oF`��#|`�A�  �9y����OK�1�k�����}<�EA��nq @D� � �q����nq?��Cᾄs�q1� ;��	l��	 |��Q�s�r�q>��u �sF`H<z�H~�H3k�7GL�zHpG�99l7�k_�B�T�F`C4��k�HJ���t��-�Ae��}�k�����s�?��  �ሏ�����EeBVT����dZ=�����ڏ ���q-�PFk�y�{FbU�= �n@6�  ���z�Fo��Be	'� � ���I� �  ��:p܋=���8ڟ웆�@�� �B�,���B���g�rAgN����  '|�X��g��B��p��BӀC׏����@ � #�Bu�&����� �b/bd�B:p2����>�m�6p�Z�=Dz?o}�܏������׿@������Ǒ��� f�?  � �M���=*�?�ff�_8�J�ܿ 3pϑ�ñ�8= �ϵʖq.·�(= ��P���'��s�t�L�>��/�;�Cd�;��.<߈�<�g�<F+�<L ��^oiΚrd�@��r6p?fff?��?&�п�@���@x��@�N��@���@T����Z���ћtމ�u �߈w	�x��ti�>�)� b�M��q������� ������:�%�^��������W���S�E� � G�=F�� Fk���������1 U@yd��� ���q��	��{� A��h�����"a��ird��A{/@w/J/5/n/vA��aA���":t�/ C^/��/Z/ ލ?��`�/�/1??���W�����g��pE� ~1�?04�0
1�1�@IӀ��Bµ�WB]�NB2��(A��@�u�\?����������b�0�|�u�R����
�>��ؽ��B�u*C��$�)�`�? ����GC#����rAU�����1�eG���I��mH�� I:��I�6[F�﫹C4OI���J�:\IT��H
~QF�y��Ol@�*J��/ I8Y�I��KFjʻC�� -?�O�O__>_)_b_ M_�_�_�_�_�_�_�_ o�_(oo%o^oIo�o mo�o�o�o�o�o �o $H3lW�{ �������2� �V�h�S���w����� ԏ�������.��R� =�v�a�������П�� ��ߟ��<�'�`�K� ]���������ޯɯ�@�&�8�#�\��3(J�ϳ�3:a������J�3��c4��������������ǲ��ڿ�n�����e��n�4 �{2�2�r�`ϖτϺϔ���%PR�P���! �h�!�K�6�o�Z�����u�|ߵߠ� ���������3��W� B�{�f�4���������d�A����!��1� 3�E�{�i��������������  2 E�f�7Fb�7�b�6B�!�!� C9� 	�� n�@�/`r� �����#x�� +=�3?, V*�8v�n�n��un��.
 D �����//%/ 7/I/[/m//�/�:�� ��ֻ�G����$PARAM_MENU ?2���  �DEFPU�LSE�+	WAITTMOUT�+�RCV? �SHELL_WR�K.$CUR_S�TYL� 4<OsPTJJ?PTB_?�Y2C/?R_DECSN 0�Ű<�?�?�? �?�?OO?O:OLO^O��O�O�O�O�O�!SS�REL_ID  �.����EUSE�_PROG %��*%�O0_�CCCR�0�B��#CW_HO�ST !�*!HT�_=ZT��O_�Sh_�zQ�S�_<[_TI�ME
2�FXU� GDEBUG�@�+�C�GINP_FLM3SKo5iTRDo5gWPGAb` %l��tkCHCo4hTYPE�,� �O�O�o #0Bkfx� �������� C�>�P�b��������� ӏΏ�����(�:��c�^�p�����7eWO�RD ?	�+
 �	RSc`n��PNS��C4�J9Ov1��TE�P�COL�է�2��g�LP 3��n���OjTRACECToL 1�2��! ��Ғ����q�DT Q�2��Ǡ��D � ��ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ����Я0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~�T�� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�3��$PGTRACELEN  �1�  ����0��6_UP �����A�@�1  @�1_C�FG �ET�3�1
@�<D<D�VOaG�0uO$BDEF�SPD �/L��1�0��0H_C�ONFIG �\E�3 �0�05d�D��2 �1�A�PpDsA�A�0�AI�N'@TRL �d/MOA8pEQPE�E;��G�A<D\�AILID(C�/M�	bTGRP 1þ�I l�1B  �����1�A�33FC� �F8� E�� @eN	�A�AsA�Y�Y��A�@� 	 pvO�Fg�_ ´8cokB;`baBo,o>o�xobo�o�1>о�?B/�o�o~�o� =%<���
C@yd� �"������  Dz@�I�@A0� q� �������ˏ��� ڏ���7�"�4�m�X�Б�|���Ú)ґ
�V7.10bet�a1HF @�{���Aq��Qn  �?� ��BܠP�p �C���&�B�EQAA���Q�P�Q�� ß [�m����<CA��0 �b�A��̯ޯ�GeQ�KNOW_M  �lE7FbTSV ĽJ�BoC_�b� t�������������1��]aSM�SŽK ����	NE����ĿK���ODbb��A�RP�����0�Ŗ� @bQMR�S��T�iN����d���V]ST�Q1� 1�K
 4 MU�i��c�kFK�]�o� �ߓߥ߷�������2� �#�h�G�Y��}�� �����
������,��27�I��1�<t�H��P3^�p������,�4��������,�5 (:,�6Wi{�,�7�����,�8�!3,�M�AD�6 ER�O�VLD  K�D�xO.�PARNU�M  �/�T�_SCH� E
�9'!G)�3Y%UPD�/%�E�/P�_CM�P_��0@�0'�7E�$ER_CHK��%5H�&�/�+RS8���bQ_MO�+?�=5_'?O�_RES_G6��:�I�o�? �?�?�?O�?O7O*O [ONOOrO�O�O�{4]��<�?�Oz5���O __|3 #_B_G_|3 V b_�_�_|3� �_�_ �_|3� �_�_o|3O�o>oCo|2V 1��:�k1!�@c?��=2THR_INR�c0i!�o5d�fMA�SS�o Z�gMN��o�cMON_QU?EUE �:�"�Tj0��t4N� U1qNv�+DpENDFqd?`yEXEo`u� �BEnpPAsOPT�IOMwm;DpPROGRAM %$z�%Cp}o(/BrTA�SK_I��~OCFG �$/�^K�DATA��T���j12,ź�̏ ޏ�����&�8�J�\��n��������ȟ{�IWNFO�͘��3t ��!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w�����Θ� 4�FJ�a K�_N��T��˶ECNBg ڽw1��2���GN�2�ڻ �P(O�=��=�]ϸ�@���v� �u�uɡdƷ�_EDIT ��T�����G�WERF�L�x�c)�RGAD�J Ҷ�A�  $�?j00��a�Dq�ձӆ5�?��ʨ�<u�j0涁%e������FӨ�2Y�R��	H;pl�G��b_�>�pAodɻt$�*�/� **:�j0�$�@�5Y�T���^��q��:�~�L��\� n���������� �����4�F�t�j�|� ������������b LBT�x�� ��:��$, �Pb���/� ���/~/(/:/h/ ^/p/�/�/�/�/�/�/ V? ??@?6?H?�?l? ~?�?�?�?.O�?�?O O O�ODOVO�OzO�O _�O�O�O�O�Or__ ._\_R_d_�_�_�_�_�_�_�f	g�io�pWo �o{d�o�~o�ozo�B�PREF S�Rږp�p
�?IORITY�w[�}��MPDSP�q���pwUT6����OoDUCT3������OG��_T�G��8��ʯrTOE�NT 1׶� �(!AF_IN�E�p,�7�!t�cp7�_�!u�dN���!ic�mv��ޯrXYK��v����q)� ,�����p��&�	� �R�9�v�]�o����� П������*��N�`�*�sK��9}�ߢ�\��Ư ,�/6�H�������خ�At�?,  �Hp���P�b�t����u�w�HANCE �R��:�wd��连�2s��9Ks��POR_T_NUM�s�p����_CAR�TREP{p�Ω�SoKSTA�w dʷLGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_a_seiban�o \��olߒ�}߶ߡ��� ������"���X�C� |�g���������� ���	�B�-�f�Q��� u������������� ,<bM�q� ������(|L�VERSIyp��w} di�sabledWS�AVE ߾z	�2600H76%8S?�!ؿ����/ 	5(�r)og+^/y�e{/�/�/��/�/�*�,/? ��p���_�p 1��Ћ� ������Wh?z?�W*pURGE��B�p}vgu6,�WF�0DO�vƲ©vW%��4(�C�WR�UP_DELAY� �\κ5R_HOT %Nf�q׿�GO�5R_NORM�AL&H�r6O�OZGS�EMIjO�O�O(qQ/SKIPF3��W3x=_98_J_\_] �_�_{_�_�_�_�_�_ �_	o/oAoSoowoeo �o�o�o�o�o�o�o +=aOq�� ������'���7�]�K�������)E�7$RA{���K/��zĀÁ_PARA�M�A3��K @�.�@`�61�2C�<���B�C��6$�BÀBTIF��4`�RCVTMO�Uu�c��ÀD�CRF3��I ��+Q-�H�D�3D�?ޅ�2̪>_އ��?S��:k_-_��yS;�Cd;���.<߈<��g�<F+<L����Ѱ��d�u� L�������ϯ�����)�;�M�_���RD�IO_TYPE � M=U�k�EFP�OS1 1�\�
 x4/����� +�$/<��$υ�pϩ� D���h��ό��'��� ���o�
ߓ�.ߤ�R� ��������5���Y� ��i��*�<�v���r� ��������U�@�y� ���8���\������������?��c����2 1�KԿX��T�x��3 1����nY�>S4 1�'9�K�/�'/�S5 1���/�/��/�/:/S6 1� Q/c/u/�/-??Q?�/S7 1��/�/
?�D?�?�?�?d?S8 1�{?�?�?�?WOBO�{O�?SMASK �1L��O�D�GX�NO���F&�^��M�OTEZ�Ż��Q_�ǁ�%]pA݂��P?L_RANG!Q]��_QOWER ��ŵ�P1VSM_D�RYPRG %�ź%"O�_�UTAR�T �^�ZUME_PRO�_�_4o���_EXEC_E�NB  J�e�GSPD`O`WhՅjbgTDBro�jRM�o��hINGVERS�ION Ź�#o�)I_AIR7PURhP �O(.�MMT_�@T�P#_�ÀOBOT_I/SOLC�NTV@Az'qhuNAME�l���o�JOB_OR�D_NUM ?��X#qH7�68  j1Zc�@�r
�rV��s��r�?��r?�r�pÀP?C_TIMEu�a��xÀS232>R1��� LT�EACH PEN�DANw�:GX��!O Main�tenance /Consj2�����"��No UseB�׏������p1�C�y�V�NPO�P\@�YQ�cS�oCH_L`�%^� �	ő��!U�D1:럒�R�@VGAIL�q@�Ӏ�J��QSPACE1 ;2�ż ��YR s�i�@Ct�YRԀ'{~��8�?�� ˯����"���7�2� c�u�����G���߯ѿ 򿵿�(��u�AC� c�u�����Ͻ�߿�� �ϵ��(��=�_�q� �ϕ�C߹������߱� �$��9�[�m�ߑ� ��Q������߭��� � ��	�W�i�{���M� ������5���. S�e�w�����I���� ���*?a s��E���� �/&//;/]o� �����/2/�/? "?�/7?Y/k/}/�/�/ O?�/�/�?�?�?O0O�OKA��*SY�PpM*�8.30�261 yB5/2�1/2018 gA �WPfG|�H��_TX`� !$�COMME��$USAp �$ENABLE=DԀ$INN`QpgIOR�B�@RY�E?_SIGN_�`�A�P�AIT�C�BWR�K�BD<�_TYP<�CRINDXS�@�W�@%VFRI{�_�GRPԀ$UF�RAM�rSRTOO}L\VMYHOL�A�$LENGTH�_VTEBTIRS�T�T  $S�ECLP�XUFIN�V_POS�@�$MARGI�A�$WAIT�`�ZX�2�\�VG2�GG1��AI�@�S�Q	g�`_�WR�BNO_USE�_DI�BuQ_RE�Q�BC�C]S$CUR_TCQP�R"a�^f �GP_ST�ATUS�A @� �A3`�BLk�HE$zc1�h�P@���@}_�FX �@�E_MLT_CTf�CH_�J�`CO�@�OL�E�CGQQ$�W�@w�b#tDE�ADLOCKuD�ELAY_CNT��a3qGt�a$wf _2 R1[�1$X<�2[2�{3[3$Zwy�q%Y�y�q`%V�@�c�@�b$V�`�RV�UV3oh>b�@ � �d�0ar'MSKJ�LgWaZ��C`NRK�PS_RATE�0$���S
`�Q�TAC��PRDH���e�S*��a4�At�0�DG�A 0�P��flp bquS2�ppI�#`
`�P �
�S\`  }�A�R_ENBQ� �$RUN?NER_AXI�<`�ALPL�Q�RU�TH�ICQ$FLI�P7��DTFERE�N��R�IF_CH�SU�IW��%V)�G!1����$PřA�Q�P�ݖ_JF�PR�_P�	�RV_D�ATA�A  {$�ETIM����$VALU$��	�OP_  � �A  2� �SC*��	� �$ITPa_!�SQ]PNPOU}��o�TOTL�o�DS}P��JOGLIb�N�PE_PKpc�Of�ji��PX]PTAS��$KEPT_M#IR��¤"`M�b�APq�aE�@�y�`q�g@١c�q�PG��BRK6�x���L�I��  ?�SJ�q��P�ADEz�ܠBS{OCz�MOTNv�DUMMY16Ӂ�$SV�`DE_�OP��SFSPDO_OVR
���@�LD����OR��T-P8�LE��F����6��OV��SF��F����bF�d�ƣ&c)��fQc�LCHDLY>��RECOV���`���W�PM��gŢ�R�O������_F�?�� @v�S �NVE�R�@�`OFS�PC,�CSWDٱc�ձ��X�B����TRG�š��`E_FDO��MOB_CM}���B���BLQ�¢	�Q�̄V�za�BUP�g��G
��AM���@`K�̊�e�_M!�d�AMxf�Q��T$CA����DF���HBKXd�v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�d�9�1A��9�3�A��ATIO�0��͠��US����WaAB��R+c�`tá`xDؾA��_AUXw�?SUBCPUP���S�`����3Եжc���3�FLA�B�HW_Cwp"�Ns&�]s�Aa��$UNI�TS�M�F�ATT�RIz�Z�CYC=L�CNECA����FLTR_2_F�I��TARTUP`Jp����A��LP�������_SCT*cF�_F�F_P���b�FqS��+�K�CHA/Q���*�d�RSD���Q����Q���_T�H�PROr���հE#MPJ���G�T�� �Q�DI��@y�RAILAC4/�bMX�LOf�xS��ځ���拁���+PR#�S`app��C� 	��F�UNC���RIN�`QQP� ԱRA)]R ��AƠ���AWAR֓��BLZaWrAkg�ng�DAQ�B�rkL�D�र&q�M�K���TI���j���$�@RIA_S�W��AF��Pñ�#��%%�p9r1��MsOIQ���DF_~P�(�PD"LM-�F�A�PHRDY�DORG�H; _QP�>s%MULSE~Pz�T��*�� J��Jײ���FAN_AL�MLVG��!WRN�%HARDP��Uc�O�� K2$SHADOW]�kp�a02���� STOf�+�_,^�w�AU{`R��eP_SBR�z5����:F�� �3MPINF?�\�4��3gREGV/1DG�b+cVm �C�CFL(��?�DAiP��ҌZ`�� �����Z�	� �P(Q$�A�$Z�Q V�@�[�
o� ��EG��o���kAAR���㌵�2�axG��AXEROB��RED���W�QD�_�Mh�S�YA��AF��FS�GW�RI�P~F&�STRP����E�˰EH�)�$�D�a\2kPB6P��t=V��Dv�OTO�19)���ARYL�tR0�v�3���FI&�ͣ?$LINKb!\�J�Q�_3S���E���QXYZ2�Z5N�VOFF���R�RJ�XxPB��d0s�G�cFI�03g��������_J ��'�ɲ�S&qR0LTV[6���aTBja�"�b�C���DU�F7.�TUR� X��eĂQ�2XP�ЊgFL��E���x@�`�U9Z8����� 1	)�K��Mw��F9��劂����ORQj��G;W3���#�Ґd ���uz����1�tOVE�q_�M��ё?C�uEC �uKB�v'0�x-�wH� �t���& `��qڠ �B�ё�u�q�wh�EC�h����ER��K	B�EP����AT�K�6e9e�W����AXs�'��v�/� �R ����!�� � �P��`��`�3p�Yp�1�p�� ��  �� (�� 8�� H��  X�� h�� x�� ����ޙ�DEBU�$�%3�I��·RAB����ٱ�sV��� 
d�J、��@� ��������Q���a�� �a��3q��Yq+$�`%"\<�cLAB0b�u�'�GRO���b<��B_s��"Tҳ *`�0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθ0uݸ��PNT0��?�SERVE �Z@� $`EAV�!�PO����nP�!�P@�$!Y@ � $>�TRQ"�b
=��BG�K�%"�2\��� _ � l��5�D6ER)RVb(�I��V0`;�N��TOQ:�7�L�@P
�R��e G�%�Q��� <�50F� ,h�`�z�>�RA�? 2 d!�����S�  M��p0xU ����OCuG��  ��CO�UNT6Q��FZN�_CFGF� 4#��6��TG4�_�=������Î�VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@H�EL�0��� 5b`B_BASN��RSR�6�C�SH����1�Ǌ�2���3��4��5��6ʭ�7��8��}�ROaO����P�PNLEAƭcAB)ë ��AC-Ku�INO�T��(B�$UR0� =�_P�U��!0��OU+�P�d�8j��� V��T�PFWD_KAR���� ��RE(ĉ P��P�>QUE�:RAO�p�`r0P1I� �x�j�P�f��6�QSCEM��0��� A��7STYL�SO j�DIX�&�����S!�_TMCMANR�Q��PENDIt�$KEYSWIT�CH���kHE��`BEATM83PE{@LE��>]���U��F��SpD_O_HOM# O�6@�EF�pPRaB(�A#PY�C� O�!���OV_M|b<0 �IOCM�dFQ��h�HKYA �D�Q�7��UF2��M����p�cFORC��3WAR�"�OM>|@  @S�#�o0U)SP�@1�2*&3&4E���TЕO��L���8U�NLOv�D4K$E}DU1  �SY��HDDNF� ~M�BLOB  p��SNPX_AS�� 0@�0�о81$SIZ�1�$VA{���MUL�TIP-��# A�� � $ ��� /4`�BS��0�yC���&FRIFB�O�S���3� NF�ODBUP߰�%�@3;9(�)"��Z@ mx��SI��TEs\�r�cSGL�1T�R�p&�Н3B��@�0S'TMTq�3Pg@V�BW�p�4SHOWܾ5@�SV��_Gv�� 3p$PCJ�XPИ���FB�PH�SP AW�EP@V�D�0WC� ���A00��PB XG@ XG XG$ XG5VIU6VI7VI8VI9VIAVIBVI�XG�YF��0XGFVH��XbI1�oI1|I1�I1�I1��I1�I1�I1�I1��I1�I1�I1�I1�Y1Y2UI2bI2*oI2|I2�I2�I�`��X�I2p�X�I2�I2��I2�I2�I2Y2PY�p�hbI3oI3|IU3�I3�I3�I3�IU3�I3�I3�I3�IU3�I3�I3Y3YU4�i4bI4oI4|IU4�I4�I4�I4�IU4�I4�I4�I4�IU4�I4�I4Y4YU5�i5bI5oI5|IU5�I5�I5�I5�IU5�I5�I5�I5�IU5�I5�I5Y5YU6�i6bI6oI6|IU6�I6�I6�I6�IU6�I6�I6�I6�IU6�I6�I6Y6YU7�i7bI7oI7|IU7�I7�I7�I7�IU7�I7�I7�I7�IU7�I7�I7Y7T��VP� UD�y"ՠ��
<A62���t�R��CM)D� ��M5�Rv�]��Q_h�R���e�8���<�YSL���  � �%\2�׀+4�'��W�BVALU��b��'���=FH�ID_L����HI��I���LE1_��㴦�$0C��SAC�! h ��VE_BLC�K��1%�D_CPU5ɧ 5ɛ ������C�� ��R "? � PWj��l#0��LA�1SB���ì���RUN_FLG�Ś����ĳ ����������H����z���TBC2��_# � @ B���e �S�8=�FTDC����V���3d�Q�THF������R�L�ESERV!E9��F��3�2��E��Н�X -$��LEN9��F���f�RA��W"G�W_�5�b�1��д2�MIO-�T%S60U�Ik��0�ܱF����[�DE<k�21LACEi0��CCS#0�� _MA�� j��z��TCV����z�T�������@.Bi�'A�z�'AJh�#EM5���J��@@i�)V�z���2Q �0�&@o�h��JK��V�K9��{���щ�J�0����JJ��JJ��AAL����������4��5�ӕ N1�������.�LD�_d�1* �CF�"�% `�GROUP���1�AN4�C�#~m REQUIR�ҎEBU�#��6�$Tk�2$���z�я #�& \�A�PPR� C� 0�
�$OPEN�CLOS�St��	i�
��&' �M�fЩ���W"-_MG߱7CB@�A����BBRK@NOL�D@�0RTMO_�5ӆp1J��P ��������������6��1�@ �)!�#�(� �����'��+#PATH''@!6#@!��<#� � '��1S�CA���6INF��UCJ�[1� C0@UM�(Y ��#�"������*���*��� PA�YLOA~J2L�ؠR_AN^�3L���91�)1AR_�F2LSHg2B4L�O4�!F7�#T7�#ACRL_�%�0�'��$��H��.�$H�A�2FLEX�:�J!�) P�2��D߽߫���0��* :����z�FG]D�����z���%�F1 ]A�E�G4�F�X�j�|����BE�������� ����(��X�T*�A� ���@�XI�[�m�\At�	T$g�QX<�=��2T X���emX�������� ����������+	9��2>+ �-�K0]o|�٠AT�F��4�ELFPѪs�Jڕ *� JEmCTR�!�ATN�vzHAND_VB.�q�1��$, $8`�F2Av���SW�u	#-� $$M*0.�]W�l g��PZ����A��� 1����:AK��]AkAz��LN�]UDkDzPZ G���C�ST_K�lK�N}DY��� A���� 0��<7]A<7W1�'��d�@g`�P���@����"
"J"�. M�2D%"p�H�<�~�ASYMj%0�	� j&-��-W1�/_�{8� �$���� �/�/�/�/ 3J<��:9�/�89�D_VI��v����V_UCNI�ӛ��cD1J�� ��╴�W<��n5Ŵ� w=4��9��?�?<�ucI�4�3�Oq%�H����/�j��0�D)IzuO���Oqk�N>0 �`��I��A��#���@ģ���@����IPl� 1 �� /�ME.Q�p��9�ơT}�PT@�;pG �+ Gt� ����'��T�0� $DUMMY}1��$PS_�@�RF�@  G b�n'FLA@ YP(c�|��$GLB_TP�ŗ���9 P�q��2 X� z!�ST9�� SBR�M M21_V�T�$SV_ER*0O��p����CL����A�GPO��f�GL~�E�W>�3 4H �+$YrZrW@�x��A1+�A���"j� �U.&�4 8`NZ�"��$GI�p}$�&� -� �Y�>�5� LH {��}$Fz�E��NEAR(P�N�CF��%PTAN9C�B	!JOG�@�� 6.@$JO�INTwa?pd�MS�ET>�7  x�E��HQtpS{r��up>�_8� �pU.Q�?�� LOCK_�FOV06���BGL�V�sGLt�TES�T_XM� 3�EM�P�����_�c$U&@%�w`24� �Y��5��2�d��3���CE- ���� $�KAR�QM��TP�DRA)�����VE�Cn@��IU��6���HEf�TOOL��C2V�DRE I�S3ER6��@ASCH� 7?Ox L�Q�29Z�H I��  @$RAI�L_BOXEwa��ROBO��?�~�HOWWAR�1x�_�zROLMj� �:qw�jq� �@ �O_Fkp! �d�l>�9�� �R
 O8B: �@�Y	""�OU�;��º�3ơ�r�q_�$PIP��N&`H��l�@��#@CORDEDd�p >f�fp�O�� < D ��OB⁴sd����Kӕ���qSYS�ADR��f���TCHt� = M,8`ENo��1Ak�_{�-$Cq_�f�V�WVA��> ��  &��PRE�V_RT�$E�DITr&VSHW�Rkq�֑ &R:��v�D��JA�$�a$HEAD�6�� ��z#KE:�E�C�PSPD�&JMP��L~��0R*P��Q?��1%&I��S�r�C�pNE; �q�wT'ICK�C��M�13��3HN��@ @p� 1Gu�!_GPp6���0STY'"xL�O��:�2l2?�A �t 
m G3%%$�R!{�=��S�`!�$��w`���ճ���Pˠp6SQU��E�Ҟu�TERC�0��{TSUtB �����hw&`gw�Q)�pO����@IZ��{��^�PR�kюB1�XPU���E_DO���, XS�K~�A�XI�@���UR �pGS�r� ^0�&��pY_) �ET�BPm��o��0Fo��0A|���Rԍ��a�;�SR�Cl>@P��b_�yUr��Y ��yU��yS��yS���U Ї�U���U���U�]���Ul[��Y�bXk�]C�m�����YRSC��� D h�D1S~0��Q�SP���eATހ���A]0,2~N�ADDRES<=B} SHIF{s��_2CH���I\��=q�TVsrI��AE"���a�Ce�
���
;�VW�A��F 	\��q��0l|\A@�rC�_B"R{zp����q�TXSCRE�E�Gv��1TICNA���t{�c�8�A�b?�H T1�� �B�����I��A��BE�y RRO�������� B���1UE4I# �g�!p�S���RSM]0�GUNEaX(@~Ƴ�j�S_S�ӆ��Á։񇣣�ACxY�0� 2H�pUE;�J�����@WGMT��Lֱ�Az��O	�BBL_| 9W8���K ��0s�5OM��LE/r��� TO!�s�RIG�H��BRD
�%qC�KGR8л�TEX��@����WIDTH@�� �B[�|�<���I_��Hi� L 8K���_�!=r���R:�_��Yґ�R�O6q�Mg0璴�U��h�Rm��L�UMh��FpERV�w �P���`�Nz��&�GEUR��iFP)�)� LP��(RE%@�a)ק�a�P!��f �5�6�7�8Ǣ#B�É@����tP�fW�S@�M�USR&�O <����U�Qs��FOC)��PRI�;Qm� :���TRI}P�m�UN��
��Pv��0��f%�p�'���@�0 Q�\���AG �0T� ��a>q�OS�%�R Po���8�R/�A� H�L4����U¡��SU�g��¢5��OSFF���T�}�=O�� 1R���:��S�GUN��}6�B_SUB?Ҝ��,�SRTN�`TU0g2��mCOR| D�'RAUrPE�TZ�#'��VCC��	3V �AC36MFB�1�%d�PG �Ws (#��ASTEM�a����0PE��:T3G�X �\ �ڏMOVEz�A��A�N�� ���M���LIM_X��2��2� �7�,�����ı�
�BVF�`E�+�~��024Y��IB�7��
�5S��_Rp� 2�^�� WİGp�+@��}СP��3�ZGx ���3����A�ݠCZ�D#RID����Vy08��90� De�MY_UBYd���6��@��!��X��P_Sh��3��L�KBM,�$+0DEY(#E�X`�����UM_M�U� X����ȀUSн� ���G0`PACI���а@��:��`:,�:����RE/��3qL�+��:[^��TARG��P�r���R<�\ d�`��A��$�	��ARF��SW2 ��-���@Oz�%qA7p�yREEU�U�01�,�+HK�2]g0�0qP� N� �EAM0G�WOR���MR�CV3�^ ���O*�0M�C�s	���|�REF_��� x(�+T� ����������3_RC H4(a�P�І�hrj��NA��$��0�_ ���2����L@��n�@@OU~7w6����Z��a2[��RE�p�@;0\�c�a'2]K�@SUL��]���C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��Q5(I�]7q�}�Tg`4D�`�0.`0�AP_�HUC�5SA��CMPz�F�6�5�5�0_�aR��a�1I\!yX�9XQVGFS��_ad ��M��0p�UF_x��B� �ʼ,RO��Q��'��6��UR�3GR�`.��3IDp���)�D`�;��A��~�IN��H{D���V@AJ���S͓UWmi=�0����TYLO*�5��b����bt� +�cPA� �cCACH�vR�U@vQ��Y��p�#CF�-I0sFR�XT���VNn+$HO����P !A3�XBf�(1 ����$�`VPy� ^b_'SZ313he6K3he12J�eh chG�ch�WA�UMP�j��IkMG9uPAD�i�iIMRE�$�b_SIZ�$P����0 ���ASYNBUF��VRTD)u5tq~ΓOLE_2DJ�(Qu5R��C��U��vPyQuECCUl�VEMV �U�r�WV�IRC�aIuVTP G���rv1s��5qMP#LAqa��v����0�cz � CKL�AS�	�Q�"��dC  �ѧ%ӑӠ@}�ؾ�~ �GE�Ue A|�0!�rSr�T�# 0! �r�iI��ml�vK�BG��VE�Z�PK= �v�Q�&��_HO�0��f �� >֦3�@Sp�SgLOW>�RO��ACCE���!� 9��VR�#���p:���A1D�����PAV�j��� D����M_B8"���^�JMPG ���g:�#E$SSC@��F�vPq��hݲ�vQS�`qVN��L;EXc�i T`�s�r���Q�FLD �DEsFI�3�0p2���:��VP2�V�j� �A��V|�4[`MV_PIs���t���A�@��F	I��|�Z��Ȥ����`�A���A��~�GAߥ�1 LOO��1 JC�B���Xc��^`�#P�LANE��R��1F@�c�����pr�M� [`�噴��S����f� ���Af��R�Aw�״t9U��pRKE��d�VANC�A���� k���ϲ�BwR_AA� l���2� ��p�#��m h���O K�$����2��kЍ0OU&A�"eA�
p�pSK�T�M@FVIEM 2l� ��P=���n �<<��dK�UMM�YK1P��`D6�ȡ�CU��#A�U��o $��T�IT�$PR�����OP���V�SHIF�r�p`J�Qsԙ�fOxE[$� _R�`U�# ����s��q������ G�"G�޵'�T�$��SCO{D7�CNT Q i�l�>a�-�a�;� a�H�a�V���1�+�2u1��D���� w � SMO�U�q��a�JQ���%��a_�R[�r�n׍*@LIQ�AA/`��XVR��s�n�T�L���ZABC��t�t�c�
L�Z�IP��u���LV�bcLn"���MPkCFx�v:�$��� ���DMY_L�N�������@y�w �Ђ(a�u� MCM��@CbcCART_��DPN� $J71D��=N�Gg0Sg0�BUXW|� ��UXEUL|ByX���	|��  �Z��x 	���m��YH�Db  y �80���0EIGH��3n�?(� H����$z ���|������$B� Kd'��_X��L3�RVS�F`���OVC�2' �$|�>P&��
q����5D�TR�@ �V��1�SPHX��!{� ,� *<�$�R�B2 2 ����C!�?  �L�V+�@b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/?�/�/V(7%3@/R/d/ v/�/6?�/�/�?�?�? O4OOION;4]?o? �?�?�?SO�?�?�O_@�O0_Q_8_f_N;5zO �O�O�O�Op_�O_o�8o�_MonoUo�oN;6 �_�_�_�_�_�oo%o 4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8�����Ǐ =�_�n���R���ş���ڟN;G �S џ�
���� ��W�i�{������� ï�.�������A��dW�<�N�|��� ����Ŀֿ�ޯ�� �0�B�_�R�d�꿤� �������������� *�L�^��rτ�
��� ���������&�8߸J�l�~� `ҟ @�з����ߩ��-����&�,�� �9�{�����a����� ����������A 'Y������ ���a#1��
��N;_MOD�E  ��S ���[�Y� B���
/\/*	|/�/�R4CWORK_A�D�
<wdT1R  ���� �/�� _INTVAL��+$��R_OPoTION6 ��q@V_DATA_GRP 27���D��P�/~?�/ �?�9��?�?�?�?O O;O)OKOMO_O�O�O �O�O�O�O_�O_7_ %_[_I__m_�_�_�_ �_�_�_�_!ooEo3o ioWoyo�o�o�o�o�o �o�o/eS �w������ �+��O�=�s�a��� ����͏���ߏ���9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_TI�M����ΑR ���Ƙ��5�;#U!AP"�1!��� �? E�W�i�{�����.�ï�կ�����'(�~�T"2F���d�R�I�Y��2�o+@�a얿����)�u��� �k0ϴ��_ ��  T� � �2��D�)�T D�� Q�zόϞϰ������� ��
��.�@�R�d�v���ߚ�/V凷������߽��R��;�o �W�p���
�t��D�iz$� �0 � �T"1!���� ������������ �*�<�N�`�r����� ����������& 8J\n���� ����"4FX ��࿁��� ����/`4�=/ O/a/s/�/�/�/�/�/�/�!!/ �0޲k�ݵ u�0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ ok$o6oHoZolo ~o�o�o�o�o1/�o�o  2DVhz�/ 5?������� �&�8�J�\�n����� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?�`Q�c�u��� ��� `Ò�ϯ����)� ;�M�_�q���������˿ݿ� ����3�. ���&2,���	123456�78v�h!B�!��2�Ch���0�ϵ������� ���!�3�9ѻ�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�h� K߰���������
�� .�@�R�d�v������� �������*< N`r����� ��&��J\ n������� �/"/4/F/X/j/|/ ;�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�/�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_�?L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o=_�o�o�o�o�o�o  2DVhz� ����h�������u�o.�@�R����Cz  B�� �  ���2&�� � _�
��_�  	�_�2�`Տ����_�p��	����ďi�{��� ����ß՟����� /�A�S�e�w������� ��N������+�=� O�a�s���������Ϳ ߿���'�9�K�_�������<v�_���$SCR_GRP� 1
� ��� t �ޗ� ��	 ���� �������������_�������)�a�����&�DE� DW�8���l�&�G�C�R-35iA 9�01234567�890��M-2�0��8��CR335 ��:�
����"����������:�@��Ӧ�G���&������	��]�o������:���H���>���������� �&���ݯ:��j�����g������B�Bt����������A�����  @�`��@9� ( ?�=���Ht�P
��F@ F�`z�y�� ���� �$ H��Gs^p��B��7��/ �0//-/f/Q/�/u/ �/�/�/8���P�� 7%?����"?W?-2?6�Q]? Hh�1�?t�ȭ7�� �����?-4A, �&HE@�<�@G�B�-1 3OZOlO-:HAp�H�O�O|O P�B�(�B�O�O_��EL�_DEFAULT�  �����`SHOT�STR#]A7RMI�POWERFL � i�/UYTWF�DO$V /URR�VENT 1�����NU L!�DUM_EIP�_-8�j!AF�_INE#P�_-4!'FT�_->�_;o9!��`o �*o�o�!RPC_MAIN�ojh�vo�o�c'VIS�oii��oo!TPpPU��Ydk!
PM�ON_PROXYl�VeZ�2r��]�f��!RDMO_SRV��Yg��O�!R��k��Xh,>���!
�`M��\�i���!RLSgYNC�-98֏>3�!ROS�_-<��4"��!
CE>4pMTCOM���V�kn�˟!	��CO�NS̟�Wl���!}��WASRC���Vm�c�!��USBd��XnR���No ӯ�������!��E���i�0���WRVI�CE_KL ?%��[ (%SVCPRG1��-:Ƶ2ܿ�˰3�	�˰4,�1�˰5T�Y�˰6|ρ�˰7�ϩ�˰H�����9����ȴ f�!�˱οI�˱��q� ˱ϙ�˱F���˱n� ��˱���˱��9�˱ ��a�˱߉��7߱� �_�������� )����Q����y�� '���O����w��� ������˰ ��İd�뱭�� ��=(as ^������/ �/9/$/]/H/�/l/ �/�/�/�/�/�/�/#? ?G?2?k?V?}?�?�? �?�?�?�?O�?1OCO .OgORO�OvO�O�O�O��O�O	_�O-_��_D�EV �Y��MC:5Xd�}GTGRP 2SV�K ��bx 	_� 
 ,�P5_ �_�R�_�_�_�_�_�_ 3ooWo>o{o�oto�o �o�o�o�o�o/A �_e����� ���� �=�$�6� s�Z���~���͏��� H�'�ޏK�2�o��� h�����ɟ۟��� #�5��Y�@�}�d�v� ��
�ׯ�Я���1� �*�g�N���r����� ���̿	���?�&� c�u�̯��PϽ��϶� �����)��M�4�q� X�jߧߎ��߲���� ��%�|��[���f� ������������� 3��W�i�P���t��� ������>�A (eL^���� ��� =O6 sZ�� ��� /�'//K/]/D/�/ h/�/�/�/�/�/�/�/ #?5??Y?�N?�?F? �?�?�?�?�?O�?1O CO*OgONO�O�O�O�O��O�O�O�O_kT �"V		_R_=_v_a_�_�_�_�[%��_�_�S���a�Qeo )goIo7omo[o�o�i �_�oi�o�o�o %'9o�o��o_ ������!�w �n��G�����ŏ�� �׏�O�4�s���g� ��w����������'� �K�՟?�-�c�Q�s� ���������#���� �;�)�_�M�o���ׯ �������ݿ��7� %�[ϝ��ϔ�K�m�G� ���������3�u�Z� ��#ߍ�{ߝߟ߱��� ���M�2�q���e�S� ��w������%�
� I���=�+�a�O���s� �������!��� 9']K������ q�m��5# Y���I��� ��/�1/sX/� !/�/y/�/�/�/�/�/ 	?K/0?o/�/c?Q?�? u?�?�?�??�?O�? �?�?)O_OMO�OqO�O �?�OO�O_�O__ %_[_I__�O�_�Oo_ �_�_�_�_oo!oWo �_~o�_Go�o�o�o�o �o�o	_o�oV�o/ �w�����7 �[�O��_���s� ����͏��3���'� �K�9�[���o���� ̟������#��G� 5�W�}������m�ׯ ů�����C���j� |�3�U�/���ӿ���� ��]�Bρ��u�c� �χϙ��Ͻ���5�� Y���M�;�q�_߁߃� �������1߻�%�� I�7�m�[�}������� 	������!��E�3� i������Y���U��� ����A��h�� 1������� [@	sa� �����3/W �K/9/o/]/�/�/�/ ��/�/�/�/�/?G? 5?k?Y?�?�/�?�/? �?�?�?�?OCO1OgO �?�O�?WO�O�O�O�O �O�O	_?_�Of_�O/_ �_�_�_�_�_�_�_G_ m_>o}_oqo_o�o�o �o�o�ooCo�o7 �oGm[���o ����3�!�C� i�W�������}�� Տ���/��?�e��� ��ˏU������џ� ��+�m�R�d��=�� ������߯ͯ�E�*� i��]�K�m�o����� ��ۿ��A�˿5�#� Y�G�i�k�}ϳ����� ϣ����1��U�C� e߻��ϲ��ϋ����� 	���-��Q��x�� A��=��������� )�k�P������q��� ��������C�(g� ��[Im��� � ?�3!W E{i����� ���///S/A/w/ ��/�g/�/�/�/�/ �/+??O?�/v?�/?? �?�?�?�?�?�?�?'O i?NO�?O�OoO�O�O �O�O�O/OUO&_eO�O Y_G_}_k_�_�_�__ �_+_�_o�_/oUoCo yogo�o�_�oo�o�o �o	+Q?u�o ��oe����� �'�M��t��=��� ��ˏ���ݏ�U�:� L��%���m�����ǟ ���-��Q�۟E�3� U�W�i�����ï�� )�����A�/�Q�S� e���ݯ¿������ ��=�+�Mϣ�ɿ�� ٿs��ϻ������� 9�{�`ߟ�)ߓ�%ߣ� �߷������S�8�w� �k�Y��}����� ��+��O���C�1�g� U���y��������'� ��	?-cQ� ����w�s� ;)_���O �����//7/ y^/�'/�//�/�/ �/�/�/?Q/6?u/�/ i?W?�?{?�?�?�?? =?OM?�?AO/OeOSO �OwO�O�?�OO�O_ �O_=_+_a_O_�_�O �_�Ou_�_�_o�_o 9o'o]o�_�o�_Mo�o �o�o�o�o�o5wo \�o%�}��� ��="�4���� U���y�����ӏ��� 9�Ï-��=�?�Q��� u����ҟ����� )��9�;�M���ş�� �s�ݯ˯��%�� 5���������[����� ٿǿ���!�c�Hχ� �{�ϋϱϟ����� ��;� �_���S�A�w� e߇߭ߛ������7� ��+��O�=�s�a�� �����������'� �K�9�o������_� ��[�������#G ��n��7���� ���aF� yg������ 9/]�Q/?/u/c/ �/�/�/�%/�/5/�/ )??M?;?q?_?�?�/ �?�/�?�?�?�?%OO IO7OmO�?�O�?]O�O �O�O�O�O!__E_�O l_�O5_�_�_�_�_�_ �_�_o__Do�_owo eo�o�o�o�o�o%o
 �o�o�o=sa�����o�!+q�$�SERV_MAI�L  +u!��~�OUTPUT��$�@�RV� 2�v  $�� (�q�}��SA�VE7�	�TOP1�0 2W� d 'ݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ�u���YP���FZN_�CFG �u�$�~����G�RP 2�D� ,B   A[�~+qD;� B\���  B4~��RB21��HELL��u��j�k��2�����%RSR�������
�C�.� g�Rߋ�v߈��߬������	���-�?�Q��/  �_�%Q��P��_���,p��L���ޖ�g�2,p�d����HK 1�� ��E�@� R�d������������� ����*<e`�r���OMM ������FTOV�_ENB�_���H�OW_REG_U�I�	�IMIOFWDL� �^�)/WAIT���$�V1�^�NTI�M���VA��_)_UNIT�����LCTR�YB��MB�_HDDN 2W� 2�:%0  �pQ/�qL/^/�/�/�/��/�/�/�/�"!ON�_ALIAS ?5e�	f�he�A? S?e?w?�:/?�?�?�? �?�?OO&O8OJO�? nO�O�O�O�OaO�O�O �O_"_�OF_X_j_|_ '_�_�_�_�_�_�_o o0oBoTo�_xo�o�o �o�oko�o�o, �oPbt�1�� �����(�:�L� ^�	���������ʏu� � ��$�Ϗ5�Z�l� ~���;���Ɵ؟��� �� �2�D�V�h���� ����¯ԯ���
�� .�ٯR�d�v�����E� ��п���ϱ�*�<� N�`�r�ϖϨϺ��� w�����&�8���\� n߀ߒߤ�O������� ����4�F�X�j�|� '����������� �0�B���f�x����� ��Y��������� >Pbt��� ���(:L �p����c� � //$/�H/Z/l/ ~/)/�/�/�/�/�/�/�? ?2?D?V?]3�$�SMON_DEF�PRO ����1 �*SYSTE�M*0m6REC�ALL ?}9 ( �}]?�?�?�?OO)O �?NO`O rO�O�O�O;O�O�O�O __&_�OJ_\_n_�_ �_�_7_�_�_�_�_o "o�_FoXojo|o�o�o 3o�o�o�o�o�o BTfx��/� ������>�P� b�t�������=�Ώ�� ���(���L�^�p� ������9�ʟܟ� � �$���H�Z�l�~��� ��5�Ưد���� � ��D�V�h�z�����1� ¿Կ���
�ϯ�@� R�d�vψϚ�-Ͼ��� ������*߽�N�`� r߄ߖߨ�;������� ��&��J�\�n�� ���7���������� "���F�X�j�|����� 3����������� BTfx��/� ����>P�bt���}5c�opy frs:�orderfil�.dat vir�t:\temp\�=>147.87�.149.40:8008�//)/w }-�*.d����~/�/�/5
x�yzrate 61 J/\/n/�/?#?6�'�/� �/�/�?ȓ?�?�8��mpback�/q?OO�)O }/�2mdbG *�?�?�?�O�O�O6�3x�4:\HO�@�ZO[1tO__)_ }4�Ea�O�OpE�O�_ �_�_�?�?WOrOoo 'o:O�_^O�_�o�o�o �OK_]_�O�o#6_��o�ol_}���v��$SNPX_AS�G 2�����q� P� 0 '%�R[1]@1.1,��y?��s%�!� �E�(�:�{�^����� ��Տ��ʏ���A� $�e�H�Z���~���џ ����؟�+��5�a� D���h�z�����ů� ԯ���
�K�.�U��� d�������ۿ���� ��5��*�k�N�uϡ� ���ϨϺ������1� �U�8�Jߋ�nߕ��� �����������%�Q� 4�u�X�j������ �������;��E�q� T���x��������� ��%[>e� t������! E(:{^�� ����/�/A/ $/e/H/Z/�/~/�/�/ �/�/�/�/+??5?a? D?�?h?z?�?�?�?�? �?O�?
OKO.OUO�O dO�O�O�O�O�O�O_ �O5__*_k_N_u_�_ �_�_�_�_�_�_o1o oUo8oJo�ono�o�o��d�tPARAM ��u�q W�	��jP�d9p��ht��pOF�T_KB_CFG�  �c�u�sOP�IN_SIM  �{vn��p��pRVQSTP_DSBW~r"t��HtSR Zy� � &��r��vTOP_ON_?ERR  uCy~8�PTN Zu�k�A4�RING_PRMB�� �`VCNT_�GP 2Zuq�!px 	r��ɍ����׏��wVD��ROP 1�i p� y��K�]�o������� ��ɟ۟����#�5� G�Y���}�������ů ׯ�����F�C�U� g�y���������ӿ� �	��-�?�Q�c�u� �ϙϫ���������� �)�;�M�_�qߘߕ� �߹���������%� 7�^�[�m����� ��������$�!�3�E� W�i�{����������� ����/ASe w������� +=Ovs� ������// </9/K/]/o/�/�/�/ �/�/�/?�/?#?5? G?Y?k?}?�?�?�?�?��?�?�?OO)�PRG_COUNT8v��k�GuKBENBĀ�FEMpC:t}O_U�PD 1�{T  
4Or�O�O�O __!_3_\_W_i_{_ �_�_�_�_�_�_�_o 4o/oAoSo|owo�o�o �o�o�o�o+ TOas���� ����,�'�9�K� t�o���������ɏۏ ����#�L�G�Y�k� ��������ܟן��� $��1�C�l�g�y��� ������ӯ����	�� D�?�Q�c��������� ԿϿ����)�;��d�_�q�=L_INF�O 1�E-�@ �2@���π������ ��D�<LY?SDEBUGU@�@����d�If�SP_�PASSUEB?~x�LOG  �ƕ�C��Qؑ� � ��A��UD�1:\��Uߦ�_M�PC�ݵE&�8�A���V� �A�SAV !��>�����X����SVZ�TE�M_TIME 1u"���@ 0[A�X��������$T1?SVGUNS�@VE�'�E��ASK_OPTIONU@�E�A�A+�_DI���qOG�BC2_GRP 2#�I���~��@�  C����<Ko�CFG %�z��� =���`��1�.>dO �s������ �*N9r]� ������/� 8/#/\/n/��Z+�/Z/ �/�/H/�/?�/'?? K?]�k?=�@0s?�?�? �?�?�?�?O�?OO )O_OMO�OqO�O�O�O �O�O_�O%__I_7_ m_[_}__�_�_�X�  �_�_oo/o�_SoAo co�owo�o�o�o�o�o �o=+MOa �������� �9�'�]�K���o��� ������ɏ���#��_ ;�M�k�}�������� ß�ן��1���U� C�y�g����������� ����	�?�-�c�Q� s����������Ͽ� ���)�_�Mσ�9� �ϭ�������m��� #�I�7�m�ߑ�_ߵ� ������������!� W�E�{�i������ ��������A�/�e� S�u�w����������� ��+=O��sa ������� 9']Kmo� ������#// 3/Y/G/}/k/�/�/�/ �/�/�/�/??C?�� [?m?�?�?�?-?�?�? �?	O�?-O?OQOOuO cO�O�O�O�O�O�O�O __;_)___M_�_q_ �_�_�_�_�_o�_%o o5o7oIoomo�oY? �o�o�o�o�o3! CiW���� �����-�/�A� w�e����������я ���=�+�a�O��� s�������ߟ͟��o �-�K�]�o�ퟓ������ɯ���צ��$�TBCSG_GR�P 2&ץ��  �� 
 ?�  6� H�2�l�V���z���ƿ��������(�_d�E+�?��	 HC���>Ǚ��G����C��  A�.�e�q�C;��>ǳ33��SƑ/]϶�Y��=Ȑ� ?C\  Bȹ��{B���>����,P���B�Y�z��L�H�0�$����J�\�n�����@�Ҿ�� �������=�Z�%�7���?3������	V3.00~.�	cr35��	*����
��������� 3��4��   {�CT��v�}��J2�)�������CFG [+ץ'� *�������I��.<
�<b M�q����� ��(L7p[ ������/ �6/!/Z/E/W/�/{/ �/�/�/�/.�H��/? ?�/L?7?\?�?m?�? �?�?�?�? OO$O�? HO3OlOWO|O�O��� �Oӯ�O�O�O!__E_ 3_i_W_�_{_�_�_�_ �_�_o�_/oo?oAo So�owo�o�o�o�o�o �o+O=s� E���Y���� �9�'�]�K�m����� ��u�Ǐɏۏ���5� G�Y�k�%���}����� ßşן���1��U� C�y�g�������ӯ�� ����	�+�-�?�u� c����������Ͽ� ��/�A�S�����q� �ϕϧ��������%� 7�I�[���mߣߑ� �������߷��3�!� W�E�{�i����� ��������A�/�e� S�u������������� ��+aO� s��e����� 'K9o]� ������#// G/5/k/}/�/�/[/�/ �/�/�/�/??C?1? g?U?�?y?�?�?�?�? �?	O�?-OOQO?OaO �OuO�O�O�O�O�O�O ___M_�e_w_�_ 3_�_�_�_�_�_oo 7o%o[omoo�oOo�o �o�o�o�o!3�o �oiW�{��� ����/��S�A� w�e�������я���� ���=�+�M�s�a� ��������ߟ�_	� ��_ן]�K���o��� ����ۯɯ���#�� �Y�G�}�k�����ſ ׿��������U� C�y�gϝϋ��ϯ��� �����	�?�-�c�Q� s�u߇߽߫������ ��)��9�_�M���� /����i������%� �I�7�m�[������� ������������E Wi{5���� ����A/e S�w����� /�+//O/=/_/a/ s/�/�/�/�/�/�/? '?��??Q?c??�?�? �?�?�?�?�?O�?5O GOYOkO)O�O}O�O�O��O�N  �@S� V_R�$T�BJOP_GRP� 2,�E�  ?�Vi	-R4S.;\��@�|u0{SPU �>��UT� @�@LR	 ��C� �Vf  �C���ULQLQ>�33�U�R�����U�Y?�@=�Z�C��P��ͥR�>�P  B��W$o�/gC��@g�d�Db�^����eeao�P&ff�e=��7LC/kaB� o�o�P��P�ef�b-C�p��^�g`�d�o�PL�Pt<�eVC\  �Q�@�'p�`�  �A�oL`�_wC�BrD�S�^��]�_�S�`<P�B��P�anaa`C�;�`L�w�aQo�xp�x�p:���XB$'tMP@�PCAHS��n���=�P𥅡�trd<M�g E�2pb����X�	� �1��)�W���c�� ����������󟭟�7�Q�;�I�w���;d��Vɡ�U	V3�.00RScr35QT*�QT�A��� E�'�E�i�FV#�F"wqF>���FZ� Fv�R�F�~MF����F���F��=�F���F�ъ�F��3F����F�{G
�GdG��G#
�D���E'
EMK�E���E����E�ۘE����E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F���vF�u�<#�_
<t���ٵ�=�_��V� �R�p�V9� ]E_STPARtp�H�FP*SHR\�ABL/E 1/;[%�S�G�� �W�G�BG�G� WQG�	G�E
G�GȖ�QG��G�G�ܱv�RD	I~�EQ�ϧϹ�������W�O_�q�{ߍߐ�߱���w�S]�CS  !ڄ���������� ��&�8�J�\�n��� ���������� ]\�`� ��	��(�:������
��.�@�w�NUoM  �EEQ�P	P ۰ܰw�_CFG 0���)r-PIMEBF_TTb��CSo�,GVERڳ-B,�R 11;[ 8I��R�@� �@&  ����� ��//)/;/M/_/ q/�/�/�/�/�/?�/ ?J?%?7?M?[?m?> �@�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_l�_�Y@cY�M�I_CHAN8 �c cDBGLVĂ�:cX�	`ET�HERAD ?*f�\`��?�_�uo�oQ�	`ROUT6V!	
!�d�o~�lSNMASKQh|cba255.u�ߣ'9ߣY�OOLOFS_DIb���U;iORQCT�RL 2		�Ϸ~T����� #�5�G�Y�k�}����� ��ŏ׏�����.���R�V�PE_DE�TAI/h|zPGL�_CONFIG �8�	���/�cell/$CID$/grp1V�@̟ޟ����Ӏ�o ?�Q�c�u�����(��� ϯ������;�M� _�q�����$�6�˿ݿ ���%ϴ�I�[�m� ϑϣ�2��������� �!߰���W�i�{ߍ��߱�%}F�������/�A�C�i�H� Eߞ����������?� �.�@�R�d�v���� ������������* <N`r��� ����&8J \n��!��� ��/�4/F/X/j/ |/�//�/�/�/�/�/ ??�/B?T?f?x?�? �?+?�?�?�?�?OO �?>OPObOtO�O�O�O����User� View ��}�}1234567890�O�O�O_#_`5_=T�P��]_���I2�I:O�_�_�_�_�_�_X_j_�B3�_GoYo�ko}o�o�o o�op^4 6o�o1CU�ovp^5�o���� �	�h*�p^6�c� u����������ޏp^7R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!�3� �OM�_�q��������y  e��Yz���	�� -�?�Q���uχϙ�俀����������>�� e�5i��c�u߇ߙ߫� ��d������P�)�;� M�_�q��*�<��i� ��������)���M� _�q������������ ����<�û��=Oa s��>����* '9K]f� Q�������/ �%/7/I/�m//�/ �/�/�/n<��^/? %?7?I?[?m?/�?�? �? ?�?�?�?O!O3O �/<׹��?O�O�O�O �O�O�?�O_!_lOE_�W_i_{_�_�_FOXG9 +_�_�_oo(o:o�O Kopo�o)_�o�o�o�oP�o ��	g�0�o M_q���No� ���o�%�7�I�[� m�&l�n��Ə؏ ���� ��D�V�h� ��������ԟ柍� g�ڻ}�2�D�V�h�z� ��3���¯ԯ���
� �.�@�R���3uF�� ����¿Կ������ .�@ϋ�d�vψϚϬ� ��e�w���U�
��.� @�R�d�ψߚ߬��� ��������*���w� ��v������� w�����c�<�N�`� r�����=�w��-��� ��*<��`r ����������  ��1C Ugy�����<��    -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_��  
��(  }�%( 	 y_ �_�_�_�_�_�_o	o +o-o?ouoco�o�o�o:�Z* �Q &�J\n�� ����o���9� (�:�L�^�p������ ���܏� ��$�6� }�Z�l�~�ŏ����Ɵ ؟���C�U�2�D�V� ��z�������¯ԯ� ��
��c�@�R�d�v� ����᯾�п�)�� �*�<�N�`ϧ����� �Ϻ��������&� 8��\�n߀��Ϥ߶� ��������E�"�4�F� ��j�|������� �����e�B�T�f� x�������������+� ,>Pb��� ������� (o�^p��� ���� /G$/6/ H/�l/~/�/�/�/�/ /�/�/?U/2?D?V?�h?z?�?�/�`@  �2�?�?�?�3�7�P���!frh:\�tpgl\rob�ots\m20i�a\cr35ia.xml�?;OMO_O qO�O�O�O�O�O�O�O ���O_(_:_L_ ^_p_�_�_�_�_�_�_ �O�_o$o6oHoZolo ~o�o�o�o�o�o�_�o  2DVhz� �����o�
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ �ݟ��&�8�J�\� n���������ȯߟٯ ���"�4�F�X�j�|�@������Ŀ־�8.1� �?@88�?�ֻ�ֿ� 3�5�G�iϓ�}ϟ��� ���������5��A��k�U�wߡ߿��$T�PGL_OUTP�UT ;�!�!/ ������ ��,�>�P�b�t�� ������������ (�:�L�^�p�������������2345678901������ ���"��BT fx��4�����
}$L^ p��,>���  //$/�2/Z/l/~/ �/�/:/�/�/�/�/?  ?�/�/V?h?z?�?�? �?H?�?�?�?
OO.O �?<OdOvO�O�O�ODO VO�O�O__*_<_�O J_r_�_�_�_�_R_�_ �_oo&o8o�_�_no �o�o�o�o�o`o�o�o "4F�oT|� ���\��}���@��0�B�T�e�@�������� ( 	 ��Џ����� �<�*�L�N�`����� ����ޟ̟���8� &�\�J���n�������@��ȯ���"������ �*�X�j�F�����|� ¿Կ��C���ϱ�3� E�#�i�{�忇ϱ�S� ���������/ߙ�S� e�߉ߛ�y߿���;� ������=�O�-�s� ���ߩ��]������� �'����]�o���� ��������E����� 5G%W}����� �g���1� Ug	w�{�� =O	//�?/Q/// u/�/��/�/_/�/�/ �/�/)?;?�/_?q?? �?�?�?�?�?G?�?O �?OIO[O9OO�O�? �O�OiO�O�O�O!_3_ �O_i_{__�_�_�_��_�_�R�$TPOFF_LIM >�|op:��mq�bN_SV`  �l�jP_MOoN <6�d�opop2l�aST�RTCHK =�6�f� bVTCOMPAT-h�af�VWVAR >rMm�h1d �o� �oop`ba_�DEFPROG �%|j%	Pd_DISPLAY`�|n"rINST_M�SK  t| ~^zINUSER�o�dtLCK�|}{QU?ICKMEN�dtoSCRE�p6�~�btpscdt��q��b*�_.�S�T�jiRACE_�CFG ?Mi��d`	�d
?�~u�HNL 2@|i����k r͏ߏ ���'�9�K�]�w�ITEM 2A��� �%$1234567890����  =<��П��  !���p��=��c��^��� �������.���R�� v�"�H�ί��Я��� ���*�ֿ���r�2� ������4�޿�ϰ��� &���J�\�n���@ߤ� d�v��ς������4� ��X��*��@��� ���ߨ�������T� ��x������l��� �����,�>�P����� ��FX��d����� �:�p"� �o�����F 6HZt~��N/ t/�/��// /2/�/ V/?(?:?�/F?�/�/ �/j?�??�?�?R?�? v?�?QO�?lO�?�O�O O�O*O|O_`O _�O 0_V_h_�Ot_�O__ �_8_�_
oo�_@o�_ �_�_Lodo�_�o�o4o �oXojo3�oN�or���o��s�S��B���z�  h��z ��C�:y
 P�v�]�����UD1:\������qR_GRP �1C��� 	 @Cp���$� �H�6�l�Z��|������f���˟���ڕ?�  
���<�*� `�N���r�������ޯ ̯��&��J�8�Z����	�u�����sS�CB 2D� �����(�:�L��^�pς��|V_CONFIG E����@����ϖ�OUT?PUT F�������6�H�Z� l�~ߐߢߴ������� �����#�6�H�Z�l� ~������������ ��2�D�V�h�z��� ������������
� .@Rdv��� ����)< N`r����� ��//%8/J/\/ n/�/�/�/�/�/�/�/ �/?!/4?F?X?j?|? �?�?�?�?�?�?�?O O/?BOTOfOxO�O�O �O�O�O�O�O__+O >_P_b_t_�_�_�_�_ �_�_�_oo'_:oLo ^opo�o�o�o�o�o�o �o $����!�b t������� ��(�:�-o^�p��� ������ʏ܏� �� $�6�G�Z�l�~����� ��Ɵ؟���� �2� D�U�h�z�������¯ ԯ���
��.�@�Q� d�v���������п� ����*�<�M�`�r� �ϖϨϺ�������� �&�8�J�[�n߀ߒ� �߶����������"� 4�F�W�j�|���� ����������0�B� S�f�x����������� ����,>Pa� t��������(:L/x���k}gV� K���//&/8/ J/\/n/�/�/�/W�/ �/�/�/?"?4?F?X? j?|?�?�?�?�/�?�? �?OO0OBOTOfOxO �O�O�O�?�O�O�O_ _,_>_P_b_t_�_�_ �_�O�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����o� ��� �2�D�V�h� z��������ԏ��� 
��.�@�R�d�v��� ������Ϗ����� *�<�N�`�r������� ��˟ޯ���&�8� J�\�n���������Ż��$TX_SCR�EEN 1G�g�}�ipnl/��gen.htmſ�*��<�N�`ϽPa�nel setupd�}�dϥϷ����������ω�6�H� Z�l�~ߐ�ߴ�+��� ����� �2�߻�h� z������9�g�]� 
��.�@�R�d���� �����������}� ��<N`r�� ;1��&8 �\��������QȾUALRM_MSG ?��� �Ȫ-/?/ p/c/�/�/�/�/�/�/��/??6?)?Z?%S�EV  -��6"ECFG �I��  �ȥ@�  A�1 �  B�Ȥ
  [?ϣ��?OO%O7O IO[OmOO�O�O�G�1�GRP 2J�;; 0Ȧ	 �?�O� I_BBL_N�OTE K�:T��lϢ��ѡ�0RDEF�PRO %+ (%N?u_Ѡc_�_�_ �_�_�_�_o�_o>o�)oboMo�o\INU?SER  R]�O��oI_MENHI�ST 1L�9  �(�0 ���)/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,1133�,1�oDVhz~�s� }9361 �����r�$�6� H�Z�l�~������Ə ؏����� �2�D�V� h�z�	�����ԟ� ��
���.�@�R�d�v� �������Я���� �9Rq��B�T�f�x� ��������ҿ���� ϩ�>�P�b�tφϘ� '�9���������(� ��L�^�p߂ߔߦ�5� ������ ��$���� Z�l�~����C��� ����� �2��/�h� z��������������� 
.@��dv� ����_� *<N�r��� ��[�//&/8/ J/\/��/�/�/�/�/ �/i/�/?"?4?F?X? C�U��?�?�?�?�?�? �/OO0OBOTOfO�? �O�O�O�O�O�O�O�O _,_>_P_b_t__�_ �_�_�_�_�_�_o(o :oLo^opo�oo�o�o �o�o�o �o$6H Zl~i?{?��� ���2�D�V�h� z����-�ԏ��� 
����@�R�d�v��� ��)���П����� ����N�`�r������� 7�̯ޯ���&����J�\�n�����������$UI_PAN�EDATA 1N����ڱ  	�}������!�3�E�W� ) Y�}�7�뿨Ϻ����� ���i�&��J�\�C� ��gߤߋ������������"�4��X�7�� �q}�ϕ��� ������B����%�I� [�m������
����� ������!E,i {b������l�ܳ7�<N` r����-��� //&/8/�\/n/U/ �/y/�/�/�/�/�/? �/4?F?-?j?Q?�?�? %�?�?�?OO0O �?TO�xO�O�O�O�O �O�OKO_�O,__P_ b_I_�_m_�_�_�_�_ �_oo�_:o�?�?po �o�o�o�o�oo�o  sO$6HZl~�o ������� � 2��V�=�z���s��� ��ԏGoYo�.�@� R�d�v�ɏ����П ������<�N�5� r�Y�������̯��� ׯ�&��J�1�n��� ����ȿڿ���� c�4ϧ�X�j�|ώϠ� ����+��������0� B�)�f�Mߊߜ߃��� ����������P� b�t���������� S���(�:�L�^��� ��i�����������  ��6ZlS�0w�'�9�}��� "4FX)�} ��l�����/ j'//K/2/D/�/h/ �/�/�/�/�/�/�/#?�5??Y?��C�=��$�UI_POSTY�PE  C�� 	 e?��?�2QUICKM_EN  �;�?��?�0RESTOR�E 1OC�  �L?B��6OCC1O��maO �O�O�O�O�OuO�O_ _,_>_�Ob_t_�_�_ �_UO�_�_�_M_o(o :oLo^oo�o�o�o�o �o�oo $6H �_Ugy�o��� ��� �2�D�V�h� �������ԏ�� ��w�)�R�d�v��� ��=���П������ *�<�N�`�r����� ���ޯ���&�ɯ J�\�n�������G�ȿ�ڿ�����7SCR�E�0?�=�u1sc+@u2�K�3K�4K�5K�6�K�7K�8K��2US#ER-�2�D�T,�M�SksUô�4��5�ĕ6��7��8���0N�DO_CFG �P�;� ��0PDA�TE ����None�2��_INFO 1QC�@��10%�[��� Iߊ�m߮��ߣ����� �����>�P�3�t���i���<-�OFFS_ET T�=�� ��$@������1�^� U�g������������ ����$-ZQcu���?�
�����UFRAME  �����*�RTO?L_ABRT	(��!ENB*GR�P 1UI�1Cz  A��~��@~���������0UJ�9MSK  M@�;-N%8�%��/��2VCCM��V��ͣ#RG�#Y�9����/����D�BeH�p71C����3711?�C0�$MRf2_�*S��괰	���~XC56 *�?�6�Y��1$�5����A@3C��. 	��8�?��OO KOx1FOsO�5�51ⴰ_O�O�� B����A2�DWO �O7O_�O8_#_\_G_ �_k_}_�__�_�_�_��_"o�OFoXo�%TCC�#`mI1�i���u��� GFS�»2aZ; �| 2�345678901�o�b�����o@��!5a�4BwB�`�56 311:�o=L�Br5v1�1~1�2 ��}/��o�a��# �GYk}�p�� �����ُ�1�C� U�6�H���5�~���ߏ����	���4�dSEGLEC)M!v1b3��VIRTSYN�C�� ���%�SIONTMOU�������F��#b�U��U�(�u FR:\�H�\�A\�� ��� MC��L�OG��   U�D1��EX����'� B@ �����̡m��̡R�OBCL�1�H�� �  =	 �1- n6 � -������[�,xS�A�`=��͗���ˢ��TRA�IN⯞b�a1l�
�0d�$j�T2cZ; (aE2ϖ�i�� ;�)�_�M�g�qσϕ� ���������	��F�STAT dmB~2@�zߌ�*j$i�\���_GE�#eZ;7�`0�
� 0}2��HOMIN� �fU��U�� ~�����БC�g��X���JMPERR� 2gZ;
   ��*jl�V�7������ ��������
��2�@��q�d�v�B�_ߠREr� hWޠ$LEX�ԹiZ;�a1-e��V�MPHASE  �5��c&��!OF�F/�F�P2n�jJ�0�㜳E1�@��0ϒE1!1?s#33�����ak/�@kxk䜣!W�m[�䦲�[����o3;� [ i{���� /�O�?/M/_/q/ ��/��//�/'/9/ �/=?7?I?s?�/�?�/ �/�?�??Om?O%O 3OEO�?�?�O�?�O�O �?�O�O�O__gO\_ �OE_�O�_�O�O/_�_ �_�_oQ_Fou_�_|o �o�_�oo�o�o�o�o ;oMo?qof-�oI �����7� [P��������� ˏ��!�3�(�:�i��[�ŏg�}������TD_FILTEW��n�� �ֲ:���@���+�=�O�a� s���������֯� ����0�B�T�f�x����SHIFTME�NU 1o[�<��%��ֿ����ڿ� ���I� �2��V�h� ���Ϟϰ�������3��
�	LIVE/�SNAP'�vs�fliv��E�����ION * U<b�h�menu~߃������ߣ���p����	����E�.ォ50�s�P�@� �Z�AɠB8z�z�!�}��x�~�P��� ���MERb���<�0���kMO��q���z��WAITDINE�ND������O9K1�OUT���SD��TIM����o�G���#����C���b������RELEASE������TM�������_�ACT[�����_DATA r�%L����xRD�ISb�E�$X�VR�s���$Z�ABC_GRP �1t�Q�,#�r0�2���ZIP�u'�&����[�MPCF_G 1	v�Q�0�/� �w�ɤ� 	|�Z/  85�`�/�/H/�/l$?��+ �/�/�/?�/�/???|r?�?  �D0 �?�?�?�?�?�;����x�]hYLI�ND֑y� ���� ,(  * VOgM.�SO�OwO�O�M i?�O�O^PO1_ �OU_<_N_�_�O�_�_ �__�_�_x_-ooQo�8o�_�o�oY&#2z� ���oC� e?a?>N|�oq��햋qA�$DSPH�ERE 2{6M� �_�;o���!�io |W�i��_��,��Ï ���Ώ@��/�v��� e�؏��p�����������ZZ�� � N