��   u��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����UI_CON�FIG_T  �� A$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�62�ODE�
3�CFOCA �4VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�;�  &USTOM~0 t $} RT_SPID�r,DC4D*PAG� �?^DEVIC�EPISCREuE�F��IGN�@$/FLAG�@C��1  h 	$P�WD_ACCES� E �8��C��!�%)$LABE�� $Tz jа@�3�B�	CUS�RVI 1  < `�B*�B��A7PRI�m� t1�RPTRIP�"m��$$CLA�@ O���sQ��R��RhP\ SI�qW�  �5�QIRTs1q_�P'�2 L3hL3!�pR	� ,��$?����R�P�S�S��Q@o�P� � o��
 ���)/SOFTP�.@/GEN�1?c�urrent=m�enupage,?1133,18o�o��o�o��Mo_o,13�88vo/A �'�o�n9�o�����ocmc480`|�%�7�I� �zQ a�s���������͏\� ���'�9�K�ڏo� ��������ɟX���� �#�5�G�Y��}��� ����ůׯf������1�C�U��� TPTX��y��|��o� s �o����$/soft�part/gen�link?hel�p=/md/tpia.dgd����"��4��r&ɿۻpwd 꿁ϓϥϷ������ ���#�5���Y�k�}� �ߡ߳�B�T�������1�C����zQ2'f	oC ($�ߕ����������i zQ�Q�c�Sj�n������
)��Q(a)��*����� c ��P����@�"�n�����P#`  �V������S�B 1�XR �\ }%`�REG VED��� whol�emod.htm�4	singlE�doub\t�riptbrows�@�!�� ��/AS|��/Adev.EsJl�o�1�	t���w�G/ Y/k/5/�/�/�/�/�/ ?� �P?*?<? N?`?r?�?�?�?�?�6 �@?�?�?�? O2ODO E	�/�/wO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_� �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-??z� ������
�� O@�R�!�3�����QO cOI�ݏ��*�%� 7�I�r�m�������� ǟٟ�����_/�)� W�i�{�������ïկ �����/�A�S�e� w�����iֿ���� �0�B�T�f�x�s��� ��}Ϗ����ϭ����� >�9�K�]߆߁ߓߥ� ����������#�5� ^�Y�k�9������� ��������1�C�U� g�y������������� ��ſ2DVhz� �������
� �@R	���� �����/*/%/ 7/I/r/m//�/�/�/ �/���/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSO! �O�O�O�O�O�O�O_ _0_+T_f_5_G_�_��_�Z�$UI_T�OPMENU 1��P�QR� 
d�QfA)�*defaul�tqOZM*le�vel0 *\K	G o� So�_�Qocbtpio[2�3]�(tpst[1�heo�ouo3oEo��-
h58e01�.gif�(	m�enu5&ypHq1!3&zGr%zEt4M{4�a������� ��eB�C�U�g�y������,�prim�=Hqpage,1422,1��ݏ� ��%�0�I�[�m��葟��2���class,5�����h�)�4���130�@f�x�������5���53ʏ���� �2�
5���8ٯm���� ����4�ٿ����!�3�^I�P�Q�_k�m�]��a[ϕ�ϝftyx�m�o�amf[0�o���	��c[164�g.�59�h�a���k�Ax2uK}��azm Ww%{�ߩsK�]�6�H� Z�l�~�ɿ������� ����� �2�D�V�h�z�	���2�������� ��	��ʟ?Qcu �(T�������Ѥ1$�N`r�����ainedic����/�/�confi�g=single}&��wintpĀ  /`/r/�/�/E�W��/<{���gl[47��o�w�?���!8��� 6�i.?h?>82ڀ??`�?�?z\rLz\r4s&x�? OVx`�6O ��O�O�O�O�O�O� �O_#_5_G_Y_k_�O��_�_�_�_�_�_,$;^4$doub?%o���13ؠ&dual6i38#�,4�_Pobo�_9o,n'o9ato �o�o�o}_,>P bt����� ������o4�F�X�j� |������ď֏���=J�/,�wω¯���YOw���s�͔�������u��l�V�ȟ.��?�RO<��߬ߚ�6��u7��� �����/� A���e�w��������� N������+�=�O�
."$13�ϛϭ� ����ܿ����+�=� O���s߅ߗߩ߻��� ��"���'�9�K�]�����6d��������,$۬74��/�A�S�e�C����?��	TPTX[209�,���2�(��������1I8��
��
��0P2���1_�1�Y�tv������0�
�1�
ïqC�:4$treevi�ewA#.f3�m381,26=o�� �l����//+/ �O/a/s/�/�/�/�_B�5$oq�?)? ;?F/_?q?�?�?�?�? H?�?�?OO%O7O�/$�/�1�/r2V��O��O�O �6XO�edit2azO�O_._ @_�?���OSL_�_ �_�_~��_�_G�o} o�CoUogoyo�o�o �o�o/o�o�o	- ?Qduӥ��� �����?2�D�V� h�z������ԏ� ��
����@�R�d�v� ����)���П���� ���<�N�`�r����� %���̯ޯ���&� ��J�\�n�������3� ȿڿ����"��_�_ X�o|��o��ϱ��� �������ߋ�)�S� e�x߉ߛ߭߿��ߓ ��,�>�P�b�t￿ ������������ (�:�L�^�p������ �������� ��$6 HZl~��� ���� 2DV hz����� �
/�./@/R/d/v/ �/7�IϾ/m��/I��� ??)?;?M?`?q?�? �/�?�?�?�?�?OO %O7O��nO�O�O�O�O �O�O%/�O_"_4_F_ X_�O|_�_�_�_�_�_ e_�_oo0oBoTofo �_�o�o�o�o�o�oso ,>Pb�o� �������� (�:�L�^�p������ ��ʏ܏/�/$��/ H��?MOk�}������� ş؟�W����1�C� U�h�y�����_Oԯ� ��
��.�y�@�d�v� ��������M����� �*�<�˿`�rτϖ� �Ϻ�I�������&� 8�J���n߀ߒߤ߶� ��W������"�4�F� ��X�|�������� e�����0�B�T����*defau�lta�2�*level8����������{� tpsOt[1]��y�tpio[23��u�������	menu7.�gif�
�13��	�5�
��
�4�u6�
ʯ?Qc u������� //�;/M/_/q/�/��/�/6"prim�=�page,74,1�/�/�/??�+?6"�&class,130?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO�~O�O�O�O�/�"18 �/�O__'_9_DON26@_u_�_�_�_�_���$UI_USE�RVIEW 1���R 
���_>��_
o�m(oQocouo�o �o<o�o�o�o�o�o );M_qo~� �����%�� I�[�m������F�Ǐ ُ������.�@� ��{�������ßf�� ����/�ҟS�e�w������F�*zoo}m��ZOOM�� W�I��$�6�H�Z��� ~�������ƿi������ �2�DϦ�max�resH�MAXRES߯E�㿬Ͼ� �����ϗ��*�<�N� `�߄ߖߨߺ���w� ������o�%�J�\�n� ���5���������� ��"�4�F�X�j��w� ����������� ��BTfx��? ������' =�t����_ ��//(/�L/^/ p/�/�/?�/�/�/7/ �/?$?6?H?Z?�/~? �?�?�?�?i?�?�?O  O2O�/?OUOcO�?�O �O�O�O�O�O
__._ @_R_d__�_�_�_�_ �_sQ