��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ��5/IRTU�AL-9LOO�R G��DD?8�?�������k,  1 <DwH82 �����D����/��Z�Z]/o/�/S/�/�/�-_ �/�/�/�;�$MNU>A�P"�� 8��=���?{��<��i��t-ｇ�D	?x
 ?t�t>2qn>|�l��F�Ͽ9�����0����+?��&�����S��R��ǿ����Ѯ���w<S���ʢ��Č��C�-�b{5��3�?���;�[�?���7J�j:>��e:>�@�0�����ãAz�D���#�
�{5��x?��o;'��7ue_��'�&�0��0��<�i8��/�ȭOĘ���^��{5?}��z�B�>�d���O0f�>>���@��>��?yB�B��hį%"�=%&C*/fO���_O�O�O�O�O�O�E��?��A��H
T�߉������1���<H)���ʠ Č� �C���%7NUM�  ��>� �"5TOOL/?4 
E3�O�_�O�_��_  ¢����ZDCF��_��_e?�+���?�YC�;��_o�=e�1#B�1�CG��)o;o�V����zC���aoso�o�_�o��o�o�o/l������33C�@:RW1fTIVyWZ