��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �� �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$�VERSI3 ����!COUPLED�� $!PP_�� CES0s!_81�s!  K2> �!� � $SOF�T�T_IDk2TOTAL_EQs 3$�0�0NO�2U �SPI_INDE�]�5Xk2SCRE�EN_(4_2SI�GE0_?q;�0P�K_FI� 	�$THKYGPA�NE�4 � DU/MMY1dDDd!ROE4LA!R�!R��	 � $TI=T�!$I��N ��Dd�Dd �Dc@�D5��F6�F7�F8�F9�G0�G�GJA�E�GbA�E�G1�G1�G �F��G2�B�1SBN_�CF>"
 8F CNV_J� ; �"�!�_CMNT�$�FLAGS]�C�HEC�8 � EL�LSETUP �� $HO30I�O�0� %�SMA�CRO�RREPR�X� D+�0��R{��T� UTOBAC�KU�0 }�)DEVIC�CTI*0�� �0�#��`B�S$INT�ERVALO#IS�P_UNI�O`_�DO>f7uiFR_F�0AIN�1��x�1c�C_WAkd�a�jOFF_O0N.�DEL�hL� ?a8A�a1b?9a�`FC?��P�1E��#�sATB�d��MyO� �cE D �[M�c��^qRE�V�BILrw�1X�I� QrR  �� OD�P�q�$NO^PM�!!�q�r/"�w@� �u�q�r�0D`S� p E R�D_E�pCq$F�SSBn&$CHK�BD_SE^eAG� G�"$SLOCT_��2=�� V�d¾%��3�0a_E�DIm   �S �"��PS�`�(4%$EP�1�1'$OP�0�2�a�p�_OK�UST1P_C� ��d��U �P/LACI4!�Q�x4�( raCOMM� ,0$D����0�`���EOWBJ0BIGA�LLOW� (�K�"(2�0VAR�a��@�2B n�L�0OUy� ,Kvay�r�PS�`�0M_O]�����CCFS'_UT~p0 "�1 �3�#�ؗ`X"�}R�0  4F IMC	M�`O#S�`��up�i �_�p�BA&�1���M/ h��pIMPEE_F �N��N���@O��Fr�D_�~�n�Dy�)F�� ��_�r0  T� '��'��DI�n0"��p:�P�$I��t����F�t X� �GRP0��M=qN�FLI�7��0UI�RE��$g"� SW�ITCH5�AX_�N�PSs"CF_L�IM� � �0EED��!��PqP�t�`PJ_dVЦMODEh�.Z`�P|Ӻ�ELBOF�  ������p� ���3���� FB/��0t�>�G� �� �WARNM�`/�p�qP��n�NST� �COR-0bFL{TRh�TRAT�P�T1�� $ACC�1a��N ��r$OcRI�o"V�RT�Ps_S��0CHG�0I��rT2��1�I��T�m���� x i#�Q�.�HDRBJ; C�Q�2L�3L�4L�5�L�6L�7L� N�9�s!6�CO`S <F +�=�O��#92�ЯLLECy�"MULTI�b�"N��1�!���0T�� �STY�"�R`�=bl�)2`��  '�`T  |� �&$��۱m��P�̱�UT�O���E��EXT�����ÁB���"2Q� (䈴![0�������<Ұ�+�� "D"���ŽQ��<煰kc��'�9�#���1���ÂM�ԽP��" q'�3�$ L� �E���P<��`A�$�JOBn�T���q�TwRIG3�% dK� ������<���\��+�zY��J0CO_M���& t�pFL�ܐBNG AgTBA� ���M��
�!�@�p� �q��0�P[`X��O�'[����0tna*���"J��_)R���CDJ��I*dJk�D�%C�`�0Z���0��P_�P��n@ ( @F RO.���&�t�IT�c�N�OM�
����S*��P`T)w@���bZ�P�d���RA�0଱2b"����
$T\����MD3�T�䢣`U31���p(5!H,Gb�T1�*E�7�c�KAb�WAb�cA4#�YNT���PDB�GD�� *(��P�Ut@X��W���AqX��a��eTAI^c�BUF��0!+� � 7n�PIVW�*5 P�7M�8�M�9
0�6F�7SI�MQS@>KEE�3PATn�^�a" 2�`#�"�L64FIX!, ���!d��bD�2Bus=CCI��:FPCH�P:BAD �aHCEhAOGhA]HW�_�0>�0_h@�f�A k���F�q\'M`#�"t�DE3�- l�p�3G��@FSOES]F gHBSU�IBS9WC���. ` ��MA�RG쀳��FAC<Lp�SLEWx`Qe�ӿ��MC��/�\pSM_JBM����QYC	g�exp��Д0 ā��CHN-�MP�#$G� Jg�_� #���1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�f�JR���rSEGF�R�PIO� ST�RT��N��cPV5���!41�r��
r�>İ�b�B�O�2` +�[���,q E`�,q`y�Ԣ}t���yaSIZ%���t��vT�s� �z�y,qRSINF}Oбc��@�k��`��`�`L��8� T`7�CRCf�ԣCC/�9��`a�uah�ub�MIN��uaD�s�#�G�D�YC��C �����e�q0��� �SEV�q�F�_�eF��N3�s�ah��X�a+p,5!�#1��!VSCA?� A䕖s1�"!3 � �`F/k��_�U��g��]@��C�� a�s���R�4� ����N�����5a�R�HANC��$LG��P�f1�$+@NDP�t�AR5@N^��a�q���c��ME�18���}0��3RAө�AZ �t���%O��FCTKѐ�s`"�S�PFADIJ�OJ�ʠ�ʠ����<���Ր��G8I�p�BMP�d�p8�Dba��AES�@	�vK�W_��BAS��| �G�5  M�=I�T�CSX[@@��!62�	$X�R��T9�{sC��N�`��~P_HEIGH�s1;�WID�0�V�T ACϰ�1Ap�Pl�<���EXPg�܈�|��CU�0MM�ENU��7�TI-T,AE�%)�ap2��a��8 P� �a�ED�E.`��P;DT��REM.���AUTH_KEY#  ������ �b��O	�.a}1ERRLH� �9 \� �q-�sOR�DB�_ID�@<l �PUN_O��Y�$SYS0��4g�j-�I�E�EV�#���_P(�PXWO��� �: $SK�7!f2%�Td�TRLn��; �'AC�`ܱ�ĠIND9DJ$.D��_��f1��f����PL�A�RWA�j���SD�A��!�+r|��UMMY9d�F�10d�&���J��<��}1PR� �
3�POS��J�=� �$V)$�q�PL~�>���S�ܠK�?����CJ�@\����ENE�@T���A���S_�REC�OR��BH z5 O�@=$LA�>$~�r2�R��`�q�U�`�_Du��0RO�@V�T[�Q�U��������! }У�PAU�S���dETURN,��MRU�  ;CRp�EWM�b�A�GNAL:s2$L�A�!?$P�X�@$P�y A �Ax�C0 #ܠDO�`X�k�W�v�q�GO_AWAY��MO�ae���]�C�SS_CCSCB� C �'N��CERI����J`u�QA�0�}��@�GAG� R�0| ��0{`��{`OF�q��5��#MA��Xf��&шLL�?D� �$���s�U�D)E%!`���O�VR10W�,�OR�|�'�$ESC_|$`�eDSBIOQ���l ��B�VIB&� �c,�����f�=pSSW���f!�VL��PL���AORMLO
�| �����d7%SC �bA1LspH�MPCh @�Ch �#h �#h 5�UU���C�'�C�'�#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$4�C��P3Wұ46$V7OLT37$$`�*�^1��$`O1*��$o��0RQY���2b4�0DH_TH�E����0SЯ4�7ALPH�4�`���7�@Q �0�qb7�rR�5�88� ×���"(��Fn�MӁ!VHBPFUAFLQ"Dt�s,��THR��@i2dB�����G(��P�VP�����������1��J2�B�E�C�E�CPSu�Y@��Fb3��� w`(V�H:U�G�
X0��FkQw�[�Na�'B���C INHBcFILT���$��W �2�T1�[ ��$h���H YАAF�sDO��Y�Rp� fg �Q�+�c5h�Q�iSh�QPL���Wqi�QTMOU�#c�i�Q \��X�gmb��vi�h�biAi�fI�aHIG��ca	xO��ܰ��W�"vAN-u!��	#�AV�H!Pa8�$P�ד#p�R_:�A(�a��B�N0�X�MCN���f1[1�qVE�p��Z2;&f��I�QO�u�rx�wGldDN{G|d��a!F>!�9��aM:�U�'FWA�:�Ml��� X�Lu��$!����!l��ZO����0%O�lF��s�13�DI�W� @��Q���_��!�CURVA԰0rC	R41ͰZ�C<�r�H� v���<�`U�<�(�f�CH�QR3�S���t0���Xp�VS_�`�$ד�F��ژ������NSTCY_ E L�����1�t�1��U��2*4�2B�NI O7������DEVI|� �F��$5�RB]TxSPIB�P�F��BYX����T�ކHNDG��G �H tn���L���Q�C���5��Lo0 H��閻�3FBP�{tFE{�5��t��T��I�DO<���uPMCS�v>��f>�t�"HOTS�W�`s�MMA�E;LE��J T���e �2��25�� O� ���HA7�E��344�0J����A�K �� MDL� 2J~PE��	A��s��tːÈ�s�JÆG!�rD"�ó�����\�T�O��W�	��/��S�LAV�L  �0INPڐ���`%��_CFd�Mw� $��ENU��OG��b�ϑ]զP�0�`ҕ�]�IDMaA�Sa��\�WR�#���"]�VE�$a�SKI�STs��sk$��	2u���J�������p	��Q���_SVh�EXCLUMqJ2M!'ONL��D�Y��|r�PE ղI_V��APPLYZP��HcID-@Y�r�_M�2=��VRFY�0��xr�1�cIOC_f�D�� 1������O���u�LS���R$D_UMMY3�!��z�S� L_TP/B�v�"���AӞ�ّ �N ���RT_$u��� ?G&r[��O D��P_BA��`�3x�!$F ��_5���H��CP�A�P�� P y$�KwARGI���� q�2O  �
��SGNZ�Q q�~P/�/PIGNs�l�$�^ sQ>ANNUN�@�T`<�U/�ߴ�LAzp�]	Z�d~,?E�FwPI�@ R �@�F?IT�	$TOTA%��d����!�M�NIY�S+���E�yA[�
DAYS\ԃADx�@��	� ��EFF_AXIb?�TI��0zCOJ�A �ADJ_RWTRQ��Up��H<P�1D �r5̀Ll�T�p? ]P�"p���mtpd��V 0@w�G���������SK�SU� ��C�TRL_CA�� �W�TRANS��6PIDLE_PAW���!��A�V���V_�l�V ��DIAGS���X� /$2�_SE�#TAC���t!�!00z*@��RR��vP�A���p ; SW��!�!�  ��ol�U���oOH��PP̱ ��IR�r��BR1K'#��"A_Ak��� x 2x�9ϐZs2���%l�W�pt*�x%R7QDW�%MSx�t5�AX�'�"��LIF�ECAL���10��N�1{"�5Z�3{"�dp5�ZU`}�MOT�N°Y$@FLA��cZOVC@p�5H�E	��SUPPOQ�ݑAq� Lj (C��1_X6�IEYRJZRJWRJ�0TH�!UC��>6�XZ_AR�p�Y2�HCOQ��S�f6AN��w$�IC�TE�Y `��CACHE�C9��M�PLAN��UFFIQ@�Ф0<Ѩ1	��6
��M�SW�EZ 8�K�EYIM�p��TM~�SwQq�wQ#���}�OCVIE� ��[ A�BGL���/�}�?����D�?��D\p�ذST��!�R� �T� �T�� �T	��PEMAI�f�ҁ��_FAKUL�]�Rц�1��U�� --�D�TRE�^<' $Rc�uS�% ;IT��BUFW}��W��N_� SUB~d��C|��Sb�q�bSAV�e�bu �B��� �gX�^P�d�u+p��$�_~`�e�p%yO�TT����sP��M0��OtT�LwAX � b��X~`9#�c_G�3N��YN_1�_�QD��1 �2M�U��T�F��H�@ g�`� p0p��Gb-sC_R�A�IK���r�t�RpoQ�u7h�qDSPq�2�rP��A�IM�c6�\����s2�U�@�A�sM*`IP���s�!D��6�TH�@n�)��OT�!6�HSDI3�ABSC���@ �Vy��� �_D^�CONVI�GÐ��@3�~`F�!�pd0��psqSCZ"����sMERk��qFB���k��pET���a6eRFU:@DUr`����x�CD,���@p�;cHR�A!��b`p�ՔՔ+PSԕ�C���C��p��ғSp�cH *�LX�:cd�Rqa� | ����W��U��U�@�U�	�U�OQU�7R��8R�9R��0T�^�1�k�1x�1��1��1���1��1��1ƪ2RԪ2^�k�2x�2��U2��2��2��2��U2ƪ3Ԫ3^�3k�Bx�3���o���3���3��3ƪ4Ԣ�EsXTk!0�d <�  7h�p�6�pO��p�����UPFDRZ$eT^`V�Gr����\䂴2REM� Fj�N�BOVM��A�oTROV�DT�`6-�MX<�IN��0�,�W!INDKЗ
xw�׀�p$DG~q 36��P�5�!D�6��RIV���2�BGE[AR�IO�%K���DN�p��J�82�P|B@�CZ_MCM�@ȴ1��@U��1�f y,②a? ��r�PI�!?I�E��Q�^�am���g�� _0Pfqg RI�9ej�k!UP2_ gh � �cTD�p ���! a����bwBAC�ri T�Ph�b�`�) OG���%���p��IFI��!�pm�>��	�PT|�"F��FMR2��j ��Ɛ+" ����\��������$�(B`x%��_ԡ�ޭ_���� M�������DGCLF�%DG�DY%LDa��5(�6�ߺ4���M���S�k��� T�sFS#p�Tl P���e�qP�p$EX_���1M2��2j� 3�5��G ����m ��Ѝ�SW��eOe6DEBUG����%GR���pUn�#BKU_�O1'�7 �@PO�I�5�5MS��OYOfswSM��E�c��@�0�0_E n� �pp �p�TE�RM�o��O�ORI+�p�GSM_���b�q�kTA�r�UP�R�s� -�1�2�n$�' o$SEyG,*> ELTO���$USE�pNFIAU"4�e1���>#$p$UFR���0`ؐO!�0����OT�'��TAƀU�#NST�PAT��P�"OPTHJ����E�P8 rF�V"ART�``%pB`�abU!REL:�aSHFT��V!�!.�(_SH+@M$���"� ��@N8r�����OVRq��rSHI�%0��UN� �aAY#LO����qIl���p�!�@��@ERV]� �1�?:�¦'�2��0%��5�%�RCq��E�ASYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba���
5Po��0�p6OeR�MY� `GR��t2b5n� � ��8��a�Uu Ԭ")�]��TOCO!S�1POP ��`�pC��������Oѥ`R%EPR3��aO�P�b�"ePR�%WU.X|1��e$PWR��3IMIU�2R_	S�$�VIS��#(AUDp��%�av" v���$H���P_AD+DR��H�G�"�Q��Q�QБR~pDp1�w H� SZ�a��e`�ex�e��SE���r���HS��MN~vx �0��%Ŕ��OL���p�<P��-��ACROxlP_!QND_C���ג�1�T �ROUP$T��B_�VpQ�A1Q�v��c_��i���i ��hx��i���i��v�ACk�IOU��D`�gfsu^d�yh�qa_D��VB`boPRM_�b�Q�TTP_אHaz{ (��OBJEr�l�P��$��LE�#��s`{ � \��u�AB_x�T~��S�@�DBGL�V��KRL�YHIoTCOU�BGY �LO a�TEM���e�>�+P'�,PSS�|�P�JQUERY�_FLA�b�HW(��\!a|`u@�3PU�b�PIO��"��]�ӂ/dԁ=dԁ�� _�IOLN��}�����CXa$SL�Z�$INPUTM_g�$IP#�P��L'���SLvpa~���!�\�W�C-�B$�I�O�pF_ASv��$L ��w �F1"G�U�B0m!��`���0HY��ڑ��(UOPs� ` ������[�ʔ[�і"�[PP�SIP�<�іI��2���P_MEMBܿ�i`� X��IP�P�b{�_N�`�����R�����bS�P��p$FOCU�SBG;� �UJ�Ƃ �  � o7�JOG�'�DISf[�J7�cx�J8��7� Im!�)�7_LAB�!�@�A��oAPHIb�Q�:]�D� J7J\���޷ _KEYt� ��KՀLMONza���$XR���ɀ��WATCH_0��3���EL��}S1y~���s� f �!qV�g� �CTR3�򲓥\aLG�D� ��R��I�
LG_SIZ���J�q I�,��I�FDT�IH�_� jV�GȴI�F�%SO� ��q �Ɩ���v��ƴ���K�S����w�kA��LN�����E��\���'�*�UȢs5��@L>�4�DAUZ�EA�pՀ�Dp��f�GH�B�ᢐBO}O��� C����PIT���� ��R{EC��SCRN��ⵖD_p�b�aMARGf�`��:���T�$L���S�s��W�Ԣ��Iԭ�JGMO�MN3CH�c��FN��R��Kx�PRGv�UF���p0��FWD��H]L��STP��V��+���Є�RS��H�@�몖Cr4��?B��� +�O�U�q��*�a2�8����Gh�0P!O��������M8�Ģv��EX��TUIv�	I��(�4�@� t�x�J0J�~�P���J0��N�a�#ANA8��O"�0VAIA��d�CLEAR�6DCS_HI"�/c�5O�O�SI��9S��IGN_�vp�q�uᛀT�d� DE�V-�LLA���B�UW`��x0T6<$U�EM��Ł�����"Qa���x0�σ�a�@OS1*�2�3�"a�`� �ࠜh�AN%�-���-�IDX�DP��2MRO��Գ!�S�T��Rq�Y{b! _�$E&C+��p.&A&&���`� L��ȟ%Pݘ��T\Q�UE�`�Ua��?_ � �@(���`�b���# �MBG_PN@ R`r��R�w�TRIN��P���BASS�a	6IR�Q6��@MC(��� ��CLDP|�� ETRQLI��0!D�O9=4FLʡh2��Aq3zD�q7��LqDq5[4q5ORG� )�2�8P�R��4/cp�4=b-4�t� �rpP[4*�L4q5S�@TO0�Qt�0*D2FRCLMC@D�?�?RIAtasMID`�D� d1���RQQprpDS3TB
`� �FᆻHAXD2���G�LE�XCES?R�ёBMhPa�͠�BD4VԨq`�`�F_A@�J�C[�O�H� K��G� \���bTf$� 橁LI�q�SREQoUIRE�#MO�\��a�XDEBU��_�P�ML� M䵔 �p���P�c�AAE�AN��
Q�q�/Ҙ&���-cDC��B�I9N�a?�RSM�Gh�� N#B��N�iPS}T9� � 4��7LOC�RI���;EX�fANG��A^�AODAQ䵗�@c$��9�ZMF�� ���f��"��%u#�ΖVSUP�%+1FX�@IGGo�� �rq�"��1��#B��$���p%#by��rx��x�vbPDATAKB�pE;���Ρ��M��n*� t�`MD�qI��)�v� �t�A�wqH�`��tDIAE��sANSW��th���uD��)�bԣ(@n$`� PCU_�aV6�ʠ�d�PLOr�"$`�R���B���B�p������ARR2>�E�  ��V��A/A d$CA�LI�@��G~�2p��!V��<$R��SW0^D"��AB�C�hD_J2SE��Q�@�q_J3M�
�G�1SP�,��@P�G�n�3m�u�3p�@B��JkC���2'AO)�IMk@{BCSKP ^:ܔ9�wܔJy�{B�Qܜ�����`_cAZ.B��?�EL<��YAOCMP�c|A�)��RT�j���11�ﰈ��@1�����:��Z��SMG��p�ԕ� ER!��}�� �INҠACk�p����b�n _�������D��/R��DIU��CD�H�@
�#a�q$�V�Fc�$x��$���`@���b���̂�E�H �$�BELP����!ACCEL���kA°�IRC_R�pG0��T!�$PS�@B2L�����W3��ط9� ٶPAT!H��.�γ.�3���p�A_��_�e�-B�`�C���_MG��$DD��ٰ��$FW�@�p����γ�����DE��PPAB�N�ROTSPE�Eu��O0��D�EF>Q����$U�SE_��JPQPCD��JY����-A �!YN�@A�L�̐�nL�MOU�NG���|�OL�y�INC U��a�¢ĻB��ӑ�AENCS���q�B��X���D�IN�IY�0���pzC�VE�����23_U ��b�/LOWL���:�O0��0�Di�B�PҠȠ ��PRC����MOS� gTMOpp�@-GPERCH  M�OVӤ �����! 3�yD!e�]�6�<�� ʓAY���LIʓdW�ɗ��:p3�.�I�TRKӥ�AY����?Q ^�Y�m�b��`p�CQ�� MOM�B?R�0u��D���y�0Â擰DUҐZ�S_BCKLSH_CY� ��o�n��TӀ���x
c��CLALJ���A��/PKCHKtO0�Su�RTY� B�q��M�1�q_
#Nc�_UMCP�	C�΂�SCL���LMTj�_L�0X����E�� �� ����m�h���6��P	C����H� �P�Ş�CN@�"XT����C�N_��N^C�kCS	F����V6����ϡpjY��nCAT�SHs�����ָ1����֙���������PAL���_P���_P0�� e���O1u�$xJaG� P{#�OG�>��TORQU(�p� a�~����Ry������"_W��^�����4t��
5z�
5I;I ;Iz�F�`�!��_8�1���VC��0�D�B�21��>	P�?�B�5JRK��<�2�6i�DBL_�SM�Q&BMD`_D9Lt�&BGRV4
D0t�
Dz��1H_���31�8JCOSEKr�EHLN�0hK�5oDt�jI���jI<1�J�LZ1�5Zc@y��1MYqA�HQB�THWMYTHET=09�NK23z�/Rln�r@CB4VCBn�CqPASfaYR<4gQt�gQ4VSBt��R?U'GTS���Cq��a���P#���Z�C$DUu ��R䂥э2�V�ӑ��Q�r�f$NE��+pIs@�|� �$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b�FP�c�j�FR�VrhVghTd��lV�jV�kV�kUV�kV�kV�kV�iHrh�f�r�m!�x�kUH�kH�kH�kH�kUH�iOclOrhO���nO�jO�kO�kO��kO�kO�kO�FF�.bTQ���E��egSPBALANCE���RLE�PH_'US�P衅F��F��FPFULC�3��3��E��1�l�UTOy_p �%T1T2t���2NW�����ǡ@��5�`�擳�T��OU���� INSE9G��R�REV��R����DIFH��1�l��F�1�;�OB��;C��2� �b�4?LCHWAR��;��ABW!��$ME�CH]Q�@k�q��AXk�P��IgU�i��� 
���!����ROB��CRY�ͥ�!*�C��_s"T �� x $W�EIGHh�9�$�cc�� Ih�.�IF� ќ�LAGK�8S�K��K�BIL?�O1D��U��STŰ�P�; �����������
�Ы�L�� � 2�`�"�DEB�U.�L&�n��PM'MY9��NA#δ�9�$D&���$���� Q �D�O_�A��� <@	���~��L�BX�P�N��+�_7�L�t��OH  �� E%��T���ѼT��<���TICK/�C��T1��%������N��c�Ã�R L�S���S�����PROM�Ph�E� $IR� X�~ ���!҇MAI�0��j���_�9����t�l�Rn�0COD��FU`�+�ID_" =����~�G_SUFF<0G 3�O����DO��ِ��R��Ǔـ��S����!{�������	�H)�_FI���9��ORDX� ����36��X������GR9�S��Z�DTD��v�ŧ�4 *�L_N�A4���K��DEF_I[�K���g��_����i��Ɠ�š���IS`i �萚����e����4�0i��Dg����D� O|��LOCKEA!�uӛϭϿ���{�u�UMz�K�{ԓ�{ԡ�{� ���}��v�Ա�� g������^���K‒Փ����!w�N�P@'���^���,`�W\��[R�x� �T�EFĨ �O?ULOMB_u��0�VISPIT�Y�A�!OY�A_�FRId��(�SI���R������)3���W�W��0��0_,�EAS %��!�& "����4p�G;� h ���7ƵCOEFF_Om���m�/��G!%�S.�߲CA�5����u�GR` � � $R�4�� �X]�TME�$`R�s�Z�/,)�ER�qT;�:䗰�  ]��LL��S�_S�V�($~�����@���� "SwETU��MEA���Z�x0�u������ g� � �� ȰID�"���!*��&P���*�F�'�� ��)3��#���"��5;`*��REC����!{ MSK_���� P	�1_USER��,��4p���D�0��VEL,2 �0���2�5S�I��0w�MTN�CFG}1��  ���Oy�NORE��3��26�0SI���� ���\�UX-�ܑPD�E�A $KE�Y_����$J3OG<EנSVIA�0WC�� 1DSWy���
��CMULT�G�I�@@C��2� �4 �#t�+�z�X�YZ��쑡���z� ޜ@_ERR��� ��S L�-���@��|s0BB$BUF-@qX17ࡐMOR�7� H	�CU�A3��z�1Q�
��3���'$��FV��2�TbG�� � �$SI�@ G�0V�O B`נOBJE<&�!FADJU�#E�ELAY' ���SD�WOU�мE1PY���=0QT i�0�W�DIR$ba�8pےʠDYN�HeT�@��R�^�X�����OPWORK�}1�,�SYSsBU@p 1SOP�aHR�!�jU�k�PR��2�ePA�0�!�cu�V 1OP��UJ��a�'�D�QIMAGb�A	��`i�IMAC�rIN,�bsRGOVRD=a�b�0�aP�`sʠ� �^u�z�LP�B�@��!P�MC_E,�Q��N"@�M�rǱ��1Ų{ �=qSL&�~0���$OVSL\G*E�D��*E2y�Ȑ�_=p �w��>p�s���s	�����y�7�=q�#}1�� @�@;���OE�R	I#A��
N��X�s�Ff��| ��PL}1�,RTv�m�ATU}SRBTRC_T(qR��B �����$ �pƱ��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���U1P(4����PX��؆��q��3�w� �P�G�5� $SUB������t�JMPWAITO�,�s��LOyCFt�!D=�CVF	ь�y����R`�0��CC_C�TR�Q�	�IGN�R_PLt�DBTeBm�P��z�BW)�d���0U@���IG�az��Iy�TNLN��"Z�R]aK� N��B�0�PE�s���r��f�wSPD}1� L	��A�`gఠ�S��UN��{���]�R!�BD�LY�2���tP��H�_PK�E��2RE�TRIEt��2�b�z���FI�B� ����8� 2���0DBGLV�L�OGSIZ$C�K%TؑUy#u�D7�_��_T1@�EM�@C\1A����R��D�F�CHECKK�R�)P�0����@&�(b�LEc�" PA9�T(���P�C߰PN�����ARh�0������PO�BORMATTnaF�f1h���02�S��UXy`	���LB��4� { rEITCH�B�7�9PL)�AL_ � $��XP)B�q� C,2D�!���+2�J3D��� =T�pPDCKyp��|oC� _ALPH�Æ�BEWQo����T���I�wp � ��b@PAYLOA,��m�_1t�2t���J3AR��؀դּ��laTIA4��5:��6,2MOMCP�Ӡ���������0BϐA�D��������PUBk`R��;���;����tQ��z4�` I$PI\Ds�oӓ1y�P��w�2�w�Z��I��I��I���p����n���y�e`�9S)b�T�SPEED� G ��(�Е��/���Е� `/�e�>��M��ЕSAMP�6V��/����ЕMO�@ 2@ �A��QP���C��n��� ��������LRf`kb��0�E9h�EIN09 ��7S.В9
yP�y�GAMM%S|���D$GET)b�P�cD]��2
�I�B�q�I�G$HID(0;A��LREXPbA8)LW VM8z)��g�:��C5�CHKKp]�0�I_��h`eT ��n�q��eT,�|��� �$�ȯ 1�iPI� RCH_D�313\��30LE�1�1\�o(Y��7 �t�MSWFL� �M��SCRc�7��@�&��%n�f�SV���PB``�'�!|�B�sS_SAV&0Xct5B3NO]�C\� C2^�0�mߗ�uٍa ��u���u:e;��1����8��D�P������� ��)��b9��e�@GE�3��V���Ml��� � �YL(��QNQSRlb fqXG�P�RR#dCQ�p� �S:AW70�B �B[�CgR:AMxP�K�CL�H���W�r�(1�n�g�M�!o�� �8F�P@}t$WP�u �P r��P5�R<�R C�R��%�6�`��� (��qsr X��OD�q�Z�Ug�ڐ>D� ��OM#w�J?\?�n?�?�?��9�b"�L:]�_��� |��X 0��bf��qf��q`���gzf��Eڐ�0�EcJ�"����FdPB���PM�QU�� �� 8L�QCO�U!5�QTHI�H�OQBpHYSY�ES��qUE�`�"�]O���  �P�@L\�UN���Cf�9O�� P��Vu���!����OGRA�ƁcB2�O�tVuI�Te �q:pINFOB�����{�qcB��s��r� (�@SLE�QS��q��p�vgqS����� 4L�E�NABDRZ�PTIONt�����Q���)��GCF��G�$�J�q^r�� R����U�g��OS_sED����� �F�R�PK��E'sNU߇وAUT$1܅COPY�����n�00MN����PRUT8R �Nvx�OU��$G[r|f�2�RGADJ����*�X_:@բ$P�����P��W��P��`} ��)�}�EX��YCDR�RGN�S.��F@r�LGO��#�NYQ_FREQR�W� �#�h�TsLAe#����ӄ ��CRE� s�I�F��sNA��%�a�_Ge#STAT�UI`e#MAIL �����q t��������ELEM�� ��/0<�FEASI ?�B��n�ڢ�vA�]� � I�p��Y!0q]�t#A�ABM����E�p<�VΡY�BA!S��Z��S�UZ���0$q���RMS_TR;�qb �� �SY�	�ǡ��$���>C��Q`	� 2� _�TM���� ��̲�@ �A��)ǅ�Ni$DOU�s]$Nj����PR+@3���rG�RID�qM�BAR�S �TY@��OTIO�p��� Hp_}��!����d�O�P/��� � �p�`PO�R�s��}���SRV���)����DI&0T������ #�	�#�4�!�5!�6!�7!�8���aF�2��Ep$VALUt��%���=b��/��� ;�.1�q�����(_�#AN�#�ғ�Rɀ(�>��TOTAL��S��PW�Il��R�EGEN�1�cX���ks(��a���`TR��R��_S� ��1����V�����⹂Z�E���p�q��Vr���V_H��DA�S����GS_Y,1�R4�S� {AR�P2� ^�IG_SE	s����2å_Zp��C_�ƂѿENHANC�a_� T ;�������INT�.��@yFPsİ_OVRsP�`p�`��Lv��o���7�}��Z�@�SL)G�AA�~�25��	��D��S�BĤD�E�U�����TE|�P���� !Y���
�J��$2�IL�_MC�x r#_��`T�Q�`��q���'�BV�C�P_� 0�mM�	V1�
V1�U2�2�3�3�4�4�
�!���� �� m�A�2IN~V�IBP���1�2��2�3�3�4�4�A@-�C2����p� MC_F,p+0�0L	11d���M50Id�%"Eã S`�R/�@K�EEP_HNADED!!`$^�j)C�Q����$��"	��#O �a_$A�!�0�#i��#REM�"�$��¨�%�!�(U}�e�$HPWD  `#_SBMSK|)G�q�U2:�P	�COLLAB� �!K5�B��� ��g��pIT�I1{9p#>D� ,��@FLAP��$SSYN �<M�`C6����UP_DLYzAA�ErDELA�04ᐢY�`AD�Q� �QSKIP=E�� ���XpOfPN1Tv�A�0P_Xp�r G�p�RU@,G��:I+� :IB1:IG�9JT�9JaР9Jn�9J{�9J9<��{RA=s� X����4�%1�QB� NFGLIC�s�@J�U�<H�LwNO_H�0�"�?��RITu��@_�PA�pG�Q� )��^�U��W��LV|�d�NGRLT�0 _q��O�  " ��OS���T_JvA V	�AP�PR_WEIGH��sJ4CH?pvTOqR��vT��LOO�Ј]�+�tVJ�е�ғA0�Q�U�S�XOB'�'�?� �J2P���7�X�T�<a43 DP=`Ԡ\"<a�q\!��RDC��L� ��рR��R�`� �R�V��jr�b�RGEp��*��cN�FLG�a8�Z���SPC�s��UM_<`^2TH�2NH��P.a 1�� m`EF11��� lQ �!#� <�p3AT� g�S� �Vr�p�tMq�Lr����HOMEwr +Rt2'r�-?@Qcu��t3'r�������4'r�'�9�K�]�o����5'r뤏��ȏPڏ����6'r�!�@3�E�W�i�{��7'r힟��ԟ����8'r��-�?�Q�c��u��S$0�q�p �� sF��`�1�"`P�����`/���-�IO[M�I֠��q�POWE�� ���0Za�0p�� ��5��$DSB� GNAL���0C�pm�S2323�� �~`��� / I3CEQP��PEp���5PIT����OPB�x0��FLOW�@T�RvP��!U���CU:�M��UXT�A��>w�ERFAC�� mU��ȳCH��'� tQ  _��>�f�Q$����OM���A�`T�P#UP%D7 A�ct�T��U�EX@�ȟ�U EFqA: X"�1RSPT�N����T ��PPaA�0o񩩕`EXP��IOS���)ԭ�_`���%��C�WR�A���ѩD�ag֕`ԦF�RIENDsaC2U�F7P����TOOLΫ�MYH C2LE�NGTH_VTE��I��Ӆ$S�E����UFINV�_���RGI��{QITI5B��X�v��-�G2-�G1@7�w�SG�X��_��UQQD=#���AS�Äd~C�`��q�� ��$$C/�S�`������S0S0 }��VERSI� ������5���I��������AA�VM_Y�2 �� 0  �5��C�O��@�r� r�	  ����S0����������������
0?QY�BS����1��� <-����� �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO�XOjO|O�O�O�OiC=C�@XLMT&�����  ��DINp�O�A�Dq�EXE�HiPV_��ATQ�z
��LARMRECOV ��RgLMDG �*�5�OLM_�IF *��`d �O�_�_�_�_j�_'o�9oKo]onm, 
 ��odb��o�o�o�o�^��$� z, A�   2D{�PPINFO u[ �Vw��������`������ �*��&�`�J���n�����DQ����
� �.�@�R�d�v����������a
PPLIC�AT��?�P���`Han�dlingToo�l 
� 
V8.30P/40Cp�ɔ_LI
88�3��ɕ$ME�
F0G�4�-

398�ɘ��%�z�
7D�C3�ɜ
�Non�eɘVr���ɞ@/6d� Vq?_ACTIVU�r�C죴�MODP����C�I��HGAP�ON���OU�P�1*��  i�m����Қ_�����1*�  �@��������Q����Կ�@�
������ ���5��Hʵl�K�HTTHKY_��/�M�S� ����������%�7� ��[�m�ߝߣߵ��� �������!�3��W� i�{���������� ����/���S�e�w� �������������� +�Oas�� �����' �K]o���� ����/#/}/G/ Y/k/�/�/�/�/�/�/ �/�/??y?C?U?g? �?�?�?�?�?�?�?�? 	OOuO?OQOcO�O�O �O�O�O�O�O�O__ q_;_M___}_�_�_�_`�_�_�_kŭ�TOp���
�DO_CLE�AN9��pcNM  !{衮o�o�o��o�o��DSPDgRYRwo��HI��m@�or���� �����&�8�J���MAXݐWdak�H�h�XWd�d���PLUGGW�Xgd���PRC)pB�`"�kaS�Oǂ2^DtSEGF0�K�  �+��o�or�������8���%�LAPOb� x�� �2�D�V�h�z��������¯ԯ�+�T�OTAL����+�U�SENUO�\� �e�A�k­�RGDI_SPMMC.����C6�z�@@Dr\�O�Mpo�:�X�_STRING 1	(��
�M!�S��
��_ITE;M1Ƕ  n�� ����+�=�O�a�s� �ϗϩϻ����������'�9�I/O SIGNAL���Tryout� ModeȵI�npy�Simul�ateḏOu�t��OVER�RLp = 100�˲In cyc�l�̱Prog� Abor��̱~u�Statusʳ�	Heartbe�atƷMH F�aul	��Aler�L�:�L�^�p�����������  ScûSaտ��-�?�Q� c�u������������� ��);M_q��WOR.�û�� ����+= Oas��������//'.PO ����M �6/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�?�?H"DEVP.�0d/ �?O*O<ONO`OrO�O �O�O�O�O�O�O__�&_8_J_\_n_PALT	��Q�o_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o�_GRIm�û9q �_as���� �����'�9�K��]�o�������'�R 	�݁Q����)�;� M�_�q���������˟ ݟ���%�7�I�ˏPREG�^����[� ����ͯ߯���'� 9�K�]�o����������ɿۿ�O��$AR�G_� D ?	����0���  	$�O�	[D�]D���O�e�#�SBN_C�ONFIG 
�0˃���}�CI�I_SAVE  �O�����#�TC�ELLSETUP� 0�%  O�ME_IOO�O�%?MOV_H���ώ��REP��J��U�TOBACK�����FRA;:\o� Q�o����'`��o���{� �� f� o�����*�!�3�`�����f������ ����o�{��&�8�J� \�n������������ ������"4FXj |������\끁  ��_i��_\ATBCKC�TL.TMP 6�.VD GIF .TP D_q��NLQ���fЗINI�P�Օ�~c�MESSAG�����8��ODE_!D����z��O�0��c�PAUSM!!�~0� (73�U/g+(Od/�/x/ �/�/�/�/�/�/??�?P?>?t?1�0$: TSK  @-��Tߞf�UPDT��d��0
&XWZD_�ENB����6ST�A�0��5"�XIS~��UNT 20���� � 	 ���z���eng�-�뷛�S�Ho�U@��H����PzF�Oo�}Cw�g�%^����.�O�Op�O�O/_2FMET߀�2CMPTAA���@�$A-��@���@����@���]5���5�(d5���P5�r�5�F*5�338]S�CRDCFG 1��6�Ь�Ź�_�_oo(o:oLo��o�Q���_�o �o�o�o�o�o]o�o >Pbt���o9�i�GR<@M/�s�/NA�/�	�i��v_ED�1��Y� 
 �%=-5EDT-�'��GETDATAU�o�9��?�j�H�
o�f�\��A��/  ���2�&�!�E���:IB���@~�ŏ׏m����3�� &۔��D��ߟJ�����9�ǟ�4���ϯ �(����]�o�����5N������(�w�@�)�;�ѿ_��6� ��gϮ�(�CϮ������+��7��V�3�z� (��z�����i����!8��&���~�]���@F�ߟ�5����9~������]����Y�0k�����CR�!� ����W�q���#�5����Y��p$�NO_DE�L��rGE_UN�USE��tIGALLOW 1���(*SY�STEM*S	�$SERV_GRp�V� : REG��$�\� NUMx�
��PMUB >ULAYNP\�PMPAL|�CYC10#�6 $\ULS�U�8:!�L�r�BOXORI��CUR_���PMCNV�10L�T4DCLI�0��	���� BN/`/r/�/�/�/�/��/���pLAL_OUT �;���qWD_ABOR=�f�q;0ITR_R�TN�7�o	;0NO�NS�0�6 
HC�CFS_UTIL� #<�5CC_�@6A 2#; �h ?�?�?O#O6]CE_OPTIOc8�qF@RIA�_Ic f5Y@�2�0F�Q�=2q&}��A_LIM�2].� ��P�]SB��KX�P
�PY�2O�Q��B�r
�qF�PQ5T1)T�R�H�_:JF_P�ARAMGP 1�<g^&S�_�_��_�_�VC�  C�d�`�o!o`U�`�`�`�Cd��Tii:a:e>eBa��GgC�`� D�� D	�`�w?퀗2HE ONFqI� E?�aG_P�;1#; �� �o1CUgy��aKPAUS�19�yC ,��� ������	�C� -�g�Q�w���������hя���rO�A�O��H�LLECT_b�B�IPV6�EN. �QF�3�NDE>�� �G�712�34567890���sB�TR����%
 H�/%)���� ���W���0�B���f� x���㯮���ү+��� ��s�>�P�b����� �����ο��K��@(�:ϓ�^�|��B!F�� �I|�IO ##��<U%e6߰'�9�K���TR�P2$��(9X�t�Y޼`�%�̓ڥH��_M[OR�3&�=��@XB��a��A �$��H�6�l�~���D~S��'�=�r_A?�a�a`��@K��R�d�P��)F�ha�A-�_�'�9�%
� k��G� ��%Z�%���`�@c.�P�DB��+���c?pmidbg��	L�`:�����p��|N  ��@���.���]�­@s<�^�
�@sg�$���fl�q��u�d1:��:J��D�EF *ۈ��)��c�buf.�txt����_�L64FIX ,������l/[Y/�/ }/�/�/�/�/
?�/.? @??d?v?U?�?�?�?��?�?�?,/>#_E -���<2ODOVO�hOzO�O6&IM��.zo�YU>���d�l
�IMC��2/��b��dU�C��20�M�QT:Uw�Cz  �B�i�A���A����Au�gB�3�*CG�B�<�=w�i�B.���B���B���5B�$�D��%B���ezVC��q�C�v�D����D-lE\D�n�j��ؤB9"��22o�DT|����� ����C�C����2
�xObi�D4cdv`�D��`/�`v`s]E��D D�` E�4�F*� E�c��FC��u[F����E��fE���fFކ3FY�F�P3�Z���@�33 ;���>L���Aw�n�,a@��@e�5Y����a���`A��w�=�`<#�*
��?�o�zJRSMOFS�T (�,bIT�1��D @3��
д��'�a��;��b�w?���<�{M�NTEST�)1O�CR@�4��>VC5`A�w�Ia+a��aORI`CTPB�fU�C�`4���rN��:d�*�qI?��5��qT_�P�ROG ��
�%�$/ˏ�t��NUSER  �U�������KEY_TBL � ����#a��	
��� !"#�$%&'()*+�,-./��:;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������������������������������������������������������������������������L�CK�
����ST�AT/��s_AUT_O_DO �	��c�INDT_EN�BP���Rpqn�`�T92����STOr`��v�XC�� 26��) 8
SONY? XC-56�"b�����@��F( �А�HRC50w���>�P�7b�t�Aff����ֿ� Ŀ����C�U� 0�yϋ�fϯ��Ϝ���������-ߜ�TRLޡ�LETEͦ ���T_SCREE�N ��k�cs���U�MM�ENU 17�� <ܹ���w��� ������K�"�4� ��X�j�������� ����5���k�B�T� z������������� ��.g>P�t ������ Q(:�^p�� ��/��;//$/ J/�/Z/l/�/�/�/�/ �/�/�/7?? ?m?D? V?�?z?�?�?�?�?�? !O�?
OWO.O@OfO�O�vO�O�O(y��REG� 8�y����`��M�ߎ�_MANU�AL�k�DBCOΊ�RIGY�9�DB�G_ERRL��	9�ۉq��_�_�_� ^QNUMLIT�pϡ�pd
�
^Q�PXWORK 1:���_5oGoYoko|}oӍDBTB_Nѧ ;������ADB_AW�AYfS�qGCP� 
�=�p�f_AL�pR��bbRY�[�
��WX_�P 1<{y�n�,�%oc�P�6�h_M��ISO��k�@L��sONTIM6X��
���vy�
��2sMOTNE�ND�1tRECO�RD 1B�� y���sG�O�]� K��{�b��������V� Ǐ�]����6�H�Z� ��������#�؟� �����2���V�şz� �������ԯC���g� �.�@�R���v�寚� 	���п���c�χ� #ϫ�`�rτϖ�Ϻ� )ϳ�M���&�8ߧ� \�G�Uߒ�߶�����@I������4�� �p 7�n���ߤ����� �����"���F�1��� |��������[����� i���BTf����bTOLEREN�C�dB�'r�`L���^PCSS_CC?SCB 3C>y�`	IP�t}�~� <�_`r�K�@����/�{�� 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�OX_�~�LL� D���&qET�c�a 7C[C��PZP\^r_ A� p� ��sp��QGPt[	� A�p�Q�_�[?� �_�[oU�p1�P�pSB�V�c �(a�PWoio{h+�o��X�o�oY��[	r�hLW���N:p�����}6ګ��c��aD@�VB��|�G����+��K� �otGhXGr��So����eB   =��Ͷa�>�tYB�� �pC(�p�q�aA"�H�S�Q -��q���ud�v���|��AfP ` 0����D^P��p@�a
�QXTHQ�$���a aW>� �a9P��b�e:�L�^�h�Hc�́PQ�RFQ� PU�z�֟�o\^�� -�?��c�u����zKCz�ů�b2᤼Щ�RD�����l)*����S̡0��]��0�.��@���EQ� �p��F�X�ѿUҁп��VSȺNSTCOY 1E��]�ڿ��K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߒ���DEVICE 1F5� MZ�۶a ��	� ��?�6�c����	{䰟���_HN?DGD G5�VP����R�LS 2H �ݠ��/�A�S�e�w������ ZPARAMG I�FgHe��RBT 2K���8р<��WPpC�*C��,`¢P�Z�z���%{�C�� 2�jMTLU,`"nPB, s��M� `}�gT�g��
B��!�bcy�[2D chz����/���/gT#I%D��C�` b!�R���A��A,�ͿBd��A��P���_C4kP�!2�C���$Ɓ�]�ffA��À��B�� ��| ���/�/�T ( ��54a5�}%/7/ d?/M?_?q?�?�?�? �?�?O�?OO%O7O IO�OmOO�O�O�O�O �O�O�OJ_!_3_�_�_ 3�_�_�_�_�_o�_ (ooLo^oЁ=?k_Io S_�o�o�o�o�o�o �o#5G�k} �������H� �1�~�U�g�y�ƏAo �Տ���2�D�/�h� S���go����ԟ���� ϟ���R�)�;��� _�q����������ݯ �<��%�7�I�[�m� ��������}�&�� J�5�n�YϒϤϏ��� ��ѿ������F�� /�Aߎ�e�w��ߛ߭� ��������B��+�x� O�a��������� ��,���%�b�M���q� ������������� �L#5�Yk} ��� ��6 1CUg��� �����	//h/ ���/w/�/�/�/�/�/ 
?�/.?@?I/[/1/ _?q?�?�?�?�?�?�? �?OO%OrOIO[O�O O�O�O�O�O�O&_�O _\_3_E_W_�_?�_ �_�_�_�_"ooFo1o joE?s_�_�om_�o�o �o�o�o0f= Oa������ ����b�9�K��� o���Ώ��[o��(� �L�7�I���m�������$DCSS_S�LAVE L����ё���_4D  �љ��CFG MMѕ��������FRA:\�ĐL-�%04d.wCSV��  }��� ���A i�CH
q�z������|���.��  �����Ρ�ޯ̩ˡҐ-��*�����_CRC_O_UT N�������_FSI ?}њ �� ��k�}�������ſ׿  �����H�C�U�g� �ϋϝϯ���������  ��-�?�h�c�u߇� �߽߫��������� @�;�M�_����� ����������%�7� `�[�m���������� ������83EW �{������ /XSew �������/ 0/+/=/O/x/s/�/�/ �/�/�/�/???'? P?K?]?o?�?�?�?�? �?�?�?�?(O#O5OGO pOkO}O�O�O�O�O�O  _�O__H_C_U_g_ �_�_�_�_�_�_�_�_  oo-o?ohocouo�o �o�o�o�o�o�o @;M_���� ������%�7� `�[�m��������Ǐ ������8�3�E�W� ��{�����ȟß՟� ���/�X�S�e�w� ������������� 0�+�=�O�x�s����� ����Ϳ߿���'� P�K�]�oϘϓϥϷ� ��������(�#�5�G� p�k�}ߏ߸߳�����  �����H�C�U�g� �������������  ��-�?�h�c�u��� ������������ @;M_���� ����%7 `[m���� ���/8/3/E/W/ �/{/�/�/�/�/�/�/ ???/?X?S?e?w? �?�?�?�?�?�?�?O 0O+O=OOOxOsO�O�O��O�O�C�$DCS�_C_FSO ?�����A P �O �O_?_:_L_^_�_�_ �_�_�_�_�_�_oo $o6o_oZolo~o�o�o �o�o�o�o�o72 DVz���� ���
��.�W�R� d�v����������� ��/�*�<�N�w�r� ��������̟ޟ�� �&�O�J�\�n����� ����߯گ���'�"� 4�F�o�j�|������� Ŀֿ������G�B�|T��OC_RPI�N_jϳ����ς��O�����1�Z�U��NSL��@&�h߱������� ��"��/�A�j�e�w� ������������ �B�=�O�a������� ����������' 9b]o���� ����:5G Y�}����� �///1/Z/U/g/ y/�/�/�/�/�/�/�/ 	?2?-???Q?z?u?�� ߤ߆?�?�?�?OO @O;OMO_O�O�O�O�O �O�O�O�O__%_7_ `_[_m__�_�_�_�_ �_�_�_o8o3oEoWo �o{o�o�o�o�o�o�o /XSew �������� 0�+�=�O�x�s����� ����͏ߏ���'��P�K�]�o����� �P�RE_CHK �P۪�A ��,8�2���� 	 8�9�K���+�q���a������� ݯ�ͯ�%��I�[� 9����o���ǿ��׿ ���)�3�E��i�{� YϟϱϏ�������� ���-�S�1�c߉�g� y߿��߯����!�+� =���a�s�Q���� �����������K� ]�;�����q������� ������#5�Ak {����� �CU3y� i������/ -/G/c/u/S/�/�/ �/�/�/�/??�/;? M?+?q?�?a?�?�?�? �?�?�?�?%O?/Q/[O mOO�O�O�O�O�O�O �O_�O3_E_#_U_{_ Y_�_�_�_�_�_�_�_ o/ooSoeoGO�o�o =o�o�o�o�o�o =-s�c�� �����'��K� ]�woi���5���ɏ�� ������5�G�%�k� }�[�������ן�ǟ ����C�U�o�A��� ��{���ӯ����	�� -�?��c�u�S����� ��Ͽ῿�����'� M�+�=σϕ�w����� m������%�7��[� m�K�}ߣ߁߳��߷� ���!���E�W�5�{� ��ϱ���e������� 	�/��?�e�C�U��� ������������ =O-s���� ]����'9 ]oM����� ��/�5/G/%/k/ }/[/�/�/��/�/�/ �/?1??U?g?E?�? �?{?�?�?�?�?	O�? O?OOOOuOSOeO�O �O�/�O�O�O_)__ M___=_�_�_s_�_�_ �_�_o�_�_7oIo'o moo]o�o�o�O�o�o �o!�o1W5g �k}����� �/�A��e�w�U��� ����я��o���� 	�O�a�?�����u��� ͟�����'�9�� ]�o�M���������ۯ ��ǯ�#�ůG�Y�7� }���m���ſ����� ٿ�1��A�g�E�w� ��{ύ�������	�� ��?�Q�/�u߇�e߫� �ߛ��������)�� �_�q�O������ �������7�I��� Y��]����������� ����!3WiG ��}���� %�A�1w�g ������/+/ 	/O/a/?/�/�/u/�/ �/�/�/?�/9?K? �/o?�?_?�?�?�?�? �?�?O#OOGOYO7O iO�OmO�O�O�O�O�O _�O1_C_%?g_y__ �_�_�_�_�_�_�_o �_+oQo/oAo�o�owo �o�o�o�o�o); U__q���� ����%��I�[� 9����o���Ǐ��� ��ۏ!�3�M?�i�� Y�������՟�ş� ���A�S�1�w���g� ���������ӯ�+��=��$DCS_S_GN QK�c���7m� 1�4-FEB-19� 11:37  � O�l�JANt�0O8:38}����� N.DѤ�࠱������h�x,�rWf*σ�^�M��  O�VERSION [��V3.5.1�3�EFLOGI�C 1RK���  	����P�?�P�N�!�PR�OG_ENB  ���6Ù�o�UL�SE  TŇ��!�_ACCLIM^����Ö��WRSTJNT��vc��K�EMOx�𘱋� ���INIT� S.�G�Z���O�PT_SL ?	�,��
 	Rg575��Y�74^ٵ6_�7_�50��1���2_�@ȭ��<�TO  Hݷ���]V�DEX��dc�����PATH ;A[�A\�g��y��HCP_CL?NTID ?��6� @ȸ�����IAG_GRP �2XK� ,`���� ��9�$�]�H������12345678�90����S�� �|�������!�� ��H���;�dC�S���6��� ��.�Rv �f��H��/ /�</N/�"/p/�/ t/�/�/V/h/�/?&? ?J?\?�/l?B?�?�? �?�?�?v?O�?4OFO $OjO|OOE��Oy� �O�O_�O2_��_T_�y_d_�_,
�B^ 4�_�_~_`Oo�O&o Lo^oI��Tjo�o.o�o �o�o�o �O'�_K 6H�l���� ���#��G�2�k� V���B]���Ǐُ��������(��L�B\D�rx�@��PC�����4  79֐�$��>� ��:�����ߟʟܟ����CT_CONF_IG Y���>��egU����STBF_TTS��
��b����Û�u�O�MAU��|�MSW_CF6�Z���  �OCV7IEW��[ɭ������-�?�Q�c� u�G�	�����¿Կ� �����.�@�R�d�v� ϚϬϾ�������� ��*�<�N�`�r߄�� �ߺ���������&� 8�J�\�n���!�� �����������4�F�`X�j�|����RC£	\�e��!*�B^�������C2g{�S�BL_FAULT� ]��ި�GP�MSKk��*�TD?IAG ^:�ա�I��UD1�: 6789012345�G�BSP�-?Qcu� ������//p)/;/M/� �
�@q��/$�TRECP��

��/ ?"?4?F?X?j?|? �?�?�?�?�?�?�?O�O0OBOi/{/xO�/U�MP_OPTIO1Nk���ATR¢l�:�	�EPMEj��O�Y_TEMP  È�3B�J��P�AP�DUNI�m�Q��YN_B�RK _ɩ�E�MGDI_STA�"U�aQSUNC_S1`ɫ �FO�_�_
�^
�^dpOoo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{�E���� �y�Q��� �2�D� V�h�z�������ԏ ���
��.�@�R�d� �z�������˟�� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i������� ��ÿݟ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�{�iߗߩ߻�տ�� ����'�9�K�]�o� ������������� �#�5�G�Y�s߅ߏ� ����i������� 1CUgy��� ����	-? Qk�}������� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?u? �?�?�?��?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_m?w_�_�_�_�? �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9Ke_W ����_�_��� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�]oy������� �ӟ���	��-�?� Q�c�u���������ϯ ����)�;���g� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�_�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�W� E�s������ߧ����� ��'9K]o �������� #5O�a�k}� E������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-?G Yc?u?�?�?��?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_Q?[_m__ �_�?�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ I_Sew��_�� �����+�=�O� a�s���������͏ߏ ���'�A3�]�o� ������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 9�K�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� �����ߑ�C�M�_� q߃ߝ��߹������� ��%�7�I�[�m�� ������������� !�;�E�W�i�{��ߟ� ����������/ ASew���� ���3�!O as������� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?+=G?Y?k?!?� �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	_#?5??_ Q_c_u_�?�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o -_7I[m�_ �������� !�3�E�W�i�{����� ��ÏՏ����%/� A�S�e�q������� џ�����+�=�O� a�s���������ͯ߯ ����9�K�]�w� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������'� 1�C�U�g߁��ߝ߯� ��������	��-�?� Q�c�u������� ����m��)�;�M�_� y߃������������� %7I[m �������� !3EWq�{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/�/+?=?O? i_?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O?� �$ENETM�ODE 1aj5��  
0054_F[P�RROR_PRO/G %#Z%6�_��YdUTABLE  #[t?�_�_�_�gdRSEV_NU�M 2R  ��-Q)`dQ_AU�TO_ENB  qPU+SaT_NO>a� b#[EQ(b�  *��`��`��`��`4`+�`�o�o�oZdHIS%c1+P�Sk_ALM 1c.#[ �4�l0+�o;M_q���o_b``  �#[aFR�zPTC�P_VER !�#Z!�_�$EXTLOG_REQ�fs�Qi,�SIZ5��'�STKR�oe��)�TOL  �1Dz�b�A '�_BWD�p��Hfܻ�D�_DI�� dj5SdDT1KRņSTEPя�P>��OP_DOt�Q�FACTORY_�TUN�gd<�DR_GRP 1e#YNad 	���FP���x̹ ���� �$��f?�� ���ǖ��ٟ� ԟ���1��U�@�y� d�v�����ӯ����LW
 J�ݖ�,��tۯ�j�U���~y�B�  B୰}���$  A@��s�@UUUӾ����|���E�� E�`�F@ F�5U�/�,��L���M���Jk�L�zp�JP��F�g�f�?�  �s��9�Y9}��9��8j�
�6��6��;��A����O ��� �� I �������[FEATU�RE fj5���JQHand�lingTool� � "
P�English� Diction�ary�def.4D St��ard�  
!� hAnal�og I/OI� � !
IX�gle ShiftI��d�X�uto S�oftware �Update  �rt sѓ�mat�ic Backu�p�3\st���ground �Edit��fd�
Came�ra`�Fd�e��CnrRndIm����3�Commo�n calib �UI�� Ethe��n��"�Moni�tor�LOAD�8�tr�Reli�aby�O�ENS�D�ata Acqu�is>��m.fd~p�iagnos���]�i�Docume�nt Viewe�J��870p�u�al Check Safety*�� cy� �hanc�ed Us��Fr�����C �xt.� DIO :�fi�� m8���end.��ErrI�L��S�������s  t KPa�r[�� ����J944F�CTN Menur��ve�M� J9l��TP InT�fa}c{�  744���G��p Mask� Exc��g�� �R85�T��Pr�oxy Sv�� � 15 J�ig�h-Spe��Sk}i
� R738�����mmunic��ons�S R�7��urr�T�d�0�22��aю�con�nect 2� {J5��Incr���stru,Қ�2 �RKAREL Cmd. L��{ua��R860h�Run-Ti��E[nvL�oa��KU�el +��s��S�/Wѹ�7�Lic�ense���ro�du� ogBoo�k(System�)�AD pMACROs,��/Offs��2�N�Ds�MH�� ����MMRC�?���ORDE� ech/Stop��t? �7 84fMi$�|� 13dx��]еи׏���Modz�w/itchI�VP��t?��. sv��2Optm�8�2��fil��I ��2�g 4 !+ulti-T������;�PCM f3unY�Po|���x4$�b&Regi� �r �Pri��F�K+7���g Numo SelW  �F�#�� Adju���60.��%|�� fe���&tat�u�!$6���%�� � 9 J6R�DM Robot�)�scove2� w561��RemUz�n@� 8 (S�>F3Servo��ҩ�)SNP�X b�I�\dcys�0}�Libr1Ӟ�H� �5� �f�0��58��Soz� tr�ssag4%^G 91�p ��d&0���p/I���  (ig TMI�LIB(MӋ�Fi3rm����gd7���Ns�Acc����0��XATX�Heln���*LR"1��Swpac�ArquzПimulaH��� �Q���Tou�Pa���I��T��c��&���ev. f.s�vUSB pYo��"�iP�a���  r"1Unexcept��`0i$/�����H59� VC"&�r��[6���Px{��RcJPRIN�V��; d T@�TS?P CSUI�� �r�[XC��#We�b Pl6�%d -c�1R�@4d��8���I�R66?0FVx�L�!FVGridK1?play C�lh�@����5RiR�R.�@���R-35iA����Asciip���"��� 51f��cUpl� � (�T����S��@ri�tyAvoidM� �`��CE��rk��Col%�@�GEuF� 5P��j}P�����
 B�L�t� 1+20C C� o�І!�J��P��y��� o�=q�b @DCS b ./��c��O��q���`�; ���qc�kpaboE4�DH�@�OTШ�main� N��1.�H��a�n.��A> aB!F#RLM���!i ��пMI Dev�  9(�1� h8j��spiJP��� �@��A"e1/�r���!hP� M-2� i��߂�^0i�p6�PC���  iA/'�Passwo�qT��ROS 4����qe�da�SN��Cli ����G6x Ar��G 47�!���5s��DER��Tsup�>Rt�I�7 (M��a�T2DV�
�3?D Tri-���H&��_8;�
�A�@�Def?����B�a: deRe p 4t0��e�+�V��st64MB DwRAM�h86�΢FRO֫0�Arc� visI�ԙ�yn��7| ), �b�Heal�wJ�\=h��Cell`��p� �sh[��� tKqw�c� - ��v���p	VCv�ty�y�s�"Ѐ6�ut��v�m���xs ���TD_0��J�,m�` 2��a[�>R� tsi�MAILYk�/F2�h���>�� 90 H��F0�2]�q�P5'���Ta1C��5����FC���U�F9�GigE�H�S�t�0/A� i�f�!2��boF�d�ri=c �O�LF�S����" H=5k�OPT ���49f8���cr�o6��@��l�Ap�A�Syn.(RS�S) 1L�\1y�rH�L� (2x5�5�d��pCVx9����es�t�$SР��> \p�ϐSSF�e$�tex�D o���A�	�� BP���a�(R00�Qirt��:���2)�D��1�e�VK�b@l Bui, n��WAPLf��0b��Va�kT�XCGM�ċD��L����[CR1G&a�YBU��Y�KfL��pf��k�\sm�ZTAf�@��
��Bf2�и��V#��s���� r���CB����
f���WEB��!��
���T�p���DT�&4 Y�V�`��EH����
F�61Z��
�R=2L�
�E (Np��F�V@�PK�B���#��Gf$1`?G���H�р�?I�e ����LDh�L��N��7\s@����`���M��d�ela<,��2�M.�� "L[P��`�?��_�%�����S���-F�TSO�W�J57��VGF܋|�VP2֥ 5\b�`0&�cV:����T;T� �<�ce�,?VPD��$�
T;F��DI):�<I�a\so<��a-�6Jc6s6�4L��M�V9R�h���Tr@i�� ���5�` �f�@ �������P
� ���|�`��Img PH��[l��I/A � VP�S��U�O�w��!%S�Skastd�pn)ǲt�� SW_IMEST�BFe�300��-Q� �_�P8B�_�Rued�_�T��!�_�S ��_bH'573o2c2��-o�NbJ5N�Iojb)�Cdo�cxE��o�_�lp� �o�TdP�o�c�B�or �2.rٱ(Jsp�EfrSEo�f1�}�r�3 RGoeELS��sL����s������B	��S\ $�F�r�yz�ftl�o~�g �o���������?�����P  �n�&�"�l ��T�@<�^��Y���e�u8Z���alib��Γ��ɟ3����埿�\v ��e\c��6�Z�f�T�v�R� VW���8S��UJ�91����i�ů[c9�1+o�w8���847�:��A4�j���Q��t6�m���vrc�.����HR���oqt�0ݿ��  ��28ޯ�460�>e3S0L�97���U�ЄϦ�60.� g�Ѐ��+��'�ܠ�Ϻ�8Lco��DM߱U"������ߕpi�߲T! L��na;�� �� �u%��ⅰI���loR�d��1a590gϱŭ���95�ϔ�	R����1��?��o�@#��1A�/���vt{UWeǟ���ￇ7�3[���7�ρ�C �W��62K�=fR���8��������d����2�ڔ����@��@" "http�����t7 ��� v R7��78����4�� ��TTPT�#	��eGPCV4/v߀�j�&Q�Fa7��$N�0�/2�rIO�)/;/M/6'.sv3�64i�oS�>l? torah?*�8|`�?��AM/�?
?�?.?0�k/��1 J`O��� ,O�tro��`�[P��OB4c.K?��g'�)�24g?�� c(B�Od�\iO�A5sb�?U_�?vi �/i��/�/Wn��`�o%�Fo�4l�$of8��oXF I)xo�cgmp\7��mp���duC��lh����o�(A�_Bt� �o]6P���m�I?�w�@���nIaO��4*O0wip�%P�?"�bsg?� ]7�YEM���8woV�J�/ե11?o��D�Ms�BC��7�J�\���(�52�XFa# AP�ڟ<�v�`/�şaqs����/�Of��1�9�VRK���ph�ք3H5+�=�IN/¤�SkiW�/�IF`��_�%��fs�$I�O�l����"<�0�$�`����\jԿz5�bO�vrouς�3(�ΤH (DϮ��? sG��|��F�Ou����@���D)O��*�3P $�FӅ�k��ϻ���럊�� �PL��ʿ��pgbox�ߦebo�&��Sh �>�R.�0w1T{����fx6�� P��D��3��#_I�\m;YEe�OԆMp�hxW�=Ete,����dct\���O$k R������Xm*��փro3��D�l�j�9��V'�  �FC���|@�ք <f?6KARE0�_��~ (Kh��.c1f���WpoO�_K�up��a���H/�j#- Eqd/�84���$qu�o��/  o2o?Vo<�7C�)��s�NJԆ�|?�3l\sy�?�40�?Τ�wio�u]?�w58�?,F�$OJ�
?Ԇ�"io�!�V��u&A���PR�ߩ5, �s��v1\  ?H552B�Q�21p0R7�8P510.R0�  nel �J614Ҡ/W?ATUP��d�8P545*�H8R6���9VCAM:�q97PCRImP\1�tPUIF�C8Q28  ingsQy0��,4P P63P @P P�SCH��DO�CVڀD �PCSUȾ��08Q0=PqpVEIOCr��� P�54Pupd�PR�69aP���PSET�pt\hPQ`Qt�8P�7`Q�!MAS�K��(PPRX�Y���R7B#POCO  \pppb36���PR�Q��b1P�d60Q$cJ539�.eHsb��vL�CH-`(�OP[LGq\bPQ0]`:��P(`HCR���4`S�aund�PM�CSIP`e0aPle5r=Ps�p(`DSW�  �  qPb0`�aPa��(`PRQ`Tq�RE`(Poas601P<cPCM�P�HcR0@q\j23�b�V�`E`�S`UPvisP`E` c�`UP�cPRS	a�bJ699E`sFRDmPs�RMCN:eH93<1PHcSNBARa�r7HLB�USM�qc�Pg52�fHTC<IP0cTMIL�e"P4�`eJ �PA�PdSoTPTX6p967PTEL�p��P�`�`4
Q8P8$Q48>a"PPX�8P95�P`[�s95qqbUEC-`wF
PUFRmP�fahQCmP90ZQV�CO�`@PVIP�%�537sQSUI�zVSX�P�SWEB�IP�SHTTIPth�rQ62aP�!tPGL���cIG؁�`c�wPGS�eIRC%�N�cH76�P�e Q��Q|�Ror��R51`P s:P�P,t53=PR8u8=Py�C�Q6]``�b�PI��q52]`sJ56E`s���P�DsCL�qPt5�\�rd�q75UP cR�8���u5P sR55]`,s� P8s��P��`CP�PP�SJ77.P0\o�6��cXRPP�cR6�ap�`��QtaT�79P`�6�4�Pd87]`�d90P0c��=P,���5�Y9ta�T91P� ���1P(S���Qpaiv�P06=P- C�PF�T	���!aLP PsTS�pL�CAB%�)I БIQ` ;�H��UPPaintPMS��Pa��D�IP|�ST�Y%�t\patPT�O�b�P�PLSR7�6�`�5�Q��WaN�N�Paic�qNN�E`�ORS�`�cR�681Pint'�FCB�P(�6x�-W`iM�r��!(`OBQ`�plug�`L�ao;t �`OPI-���rPSPZ�PPG�Q�7�`73ΒPRQ�ad�RL��(+Sp�PS��n�@��E`�� �PTS�-�� W��P�`a�pw�`��P`cFV9R�PlcV3D%�l��PBVI�SAPL��Pcyc+PAPVv1�pa_�CCGIP� - U��L�Pr;og+PCCR�`�JԁB�P �PԁK=�C"L�P��p��(h��<�P��h�̱�@g�Bـ
TX�%���7CTC�ptp��2��P927"0ҝPs�2�Qb��TC-�rm�t;�	`#1ΒTC�9`HcCTE�Per�j�EIPp.p/�Ep�P�c��I�use��-Fـvrv�F%��ăTG�P� CP��%�d� -h�H-�Tra��PCTI�p��TL� TRS���p�@Pנ��IP�PTh�M%��lexsQTMQ`vGer, �p�SC:�8��F��Pv\e�PF�IPSV"+�H�$cj�vـtr�aCTW-����CPVGF-��SV{P2mPv\fx����pc�b��e��bVP4�fx_m��-��S�VPD-��SVPF.�P_mo�`V� c�V��t\��LmPo�ve4��-�sVP�R�\|�tPV�Qe5.W`V6�*u"��P�}�o`���`��CVKd��N�IIP��CV����IPN9�Gene���D��D�R�D������  ��f谔�p�os.��inal"��n��DeR���`2��d�P��omB���on,���R�D�R��\��TXf��D$b��womp�� "N��dP��m���! ���=C-f����=F�XU�����g Fx��(��Dt II��hr�D��u�� "�<���Cx_ui X������f2��h	�Crl2��D,r9u�i�Ԣ� it2�c�0co��e"�����ا(.)�� ���� ���� IQnQ� �I[ ��{_= wo��,�bD� ��|�GG� ��݅��4 �{e� vʷ� &� 2���Z uz����{�� ��TW&wq~q 5�׷&��o? ;0��  �2� �w�y� ���W&���� ?�3�� A��e��/> �\�3&T���� 77߸� ���� ����� ֵ��&���8 �l1���S�) ����d *J� F�'s ~���� 6:0� ��,���s�- Q�{v� ��� �,�T �ZB�Lx6���6 ���6���ParD ��s>�E��j�6wdsq��F  ��p�����ЁDhel������ti-S`�� �Ob��Dbcf��O�����t OFT��P<A�_�V�Z I��D��V\�qWS��= dtle�Ea�n�(bzd��tiStv�Z�z�Ez :XWO H6�6����5 H�6H69�1�E4܀Tofkst�F� Y682�4܌`�f804�E91�g�`30oBkmon�_�E��eݱ�� q�lm��0 J�fh���B�_  ZDTrfL0�f(P7�EcklKV� �6|��D�85��ّ�m\b�����xo�k�ktq��g2.g���yL�bkLVts��IF��bk������IdG I/f��GR� �han�L��V0y��%��%ere���v��io�� ac�- A�n�h����cuACl�_�^i!r��)�g��	.�@�&� G��R630 ���p v�p�&H�f�f�un��R57v�OJavG�`Y��wowc��-ASF���O��7���SM`�����
af���rafLa�v(l�\F c�w a����?VXpoV �30��NwT "L�FFM���=����yh	a�G-�w:�� �m2.�,�xt��̹�6ԯ6��sd_�MC'V��➟D���fslm��isc.  H5522���21&dc.p�R78����0��708J6�14Vip �ATUu�@�OL�5�45ҴINTL�6��t8 (VC�A���sse�CRI��ȑ��UI����rt\rL�28�g��NRE��.f�,�63!��,�SC�H�d Ek�DOCV���p��C,�<�L��0Q�isp��EI1O��xE,�54��z��9��2\sl,��SET���lр�l�t2�J7�Ռ�MASK��̀�PRXY҇��7����OCO��J6�l�3�l�� (SVl�A�H�L�@Օ��7539Rsv���;#1��LCH����OPLGf�out�l�0��D��HCR.
svg��S@�hƌ�CSa�!�{�50���D�l�5!�lQ��DSW��S����̀���OP����7��PR����L�ұ�(Sg9d���PCM���[R0 \s��5PՄ����0���n�q� EAJ�1��N�q�2��gPRSa���69��� (AuFR�D�Խ��RMCN̪��93A�ɐC_SNBA�F9� 'HLB��� M��h4���h�2A�95z��HTCaԈ�TMI�L6�j95,��8�57.,PA1�i{to��TPTXҴ; JK�TEL��pIiL�� XpL�80ՃI)��.�!��P;�J{95��s "N�ܱ�H�UEC��7\cs�FR��<Q���C��57\{VC�Oa�,���IP1j�H��SUI�	CS�X1�AWEB�a��HTTa�8�RK62��m`��GP%v�IG %tutK�IPGSj�| RC�1_me�H76t��7P�ws_+��?x�R51�\iaw�N���H�53!���wL�8!�h�R66��H���Ԡ����@;J56��1���(N0��9�j��L��ӣR5`%�A|�5q�r��`,�8 5��{165�!��@�"5��H84�!�29��0��PJ����n B[�J77!Ԩ�R6�5h3n�d��y36P��3R6��-`;о Ԩ@��e;xeKJ87��#wJ90!�stu+��~@!䬵�k90�kop�B����@"!�p�@|BA�g*�n@!��Q��06!�@[�F�FaP�6��́,лTS� NC[�CKAB$iͰl1I���R7��@q�y�C�MS1�rog+QM��� �� TY$x�C;TOa�nv\+���1�(�,�6�con��~0��15��JN�N�%e:��P��9O�RS%x���8A�8�15[�FCBaUn�ZQ�P!��p{��CM�OB��"G��OL܀�x�OPI�$\lEr[�SŠ�T	D7�U޹�CPRQR9RL���S�V�~`���K�ETS�$1��0����3�Ԩ�FVR:1�LZQV3D$ ���BVa�SAPLn1�CLN[�PV���	rCCGaԙ��C�L�3CCRA�n� "W!B�H�CSKQn\0�p��,)�0CTPn�ЌQpe��p!$bCt�aqT0U�pCTC�tyЋRC1�1 (�s���trl,�r��
�TX��TCaerr9m�r�MC"�s���#CTE��nrr�REa�XPj�^��Grmc�^�a"�PQF!$���$p e"�rG1�tTG$�c8��QH�$SCT�I�! s��CTLqdACK�Rp)���rLa�R82��M`��YPk�.���OF��.���e�{�CN���^�1�"M�^�a�С@�Q`US��!$��M�QuW�$m�VGF�$oR MH��P2�� H5� ΐq��ΐn�$(MH[�VP�uAoY����$)��D���hg��VPF��"�MHG̑`e!�+�V/vpcm�N��ՙ�8N��$�VPRqd)�&�CV�x�V� "�X�,�1�($TIa�t�\mh��K��et!pK�A%Y�VP%ɠ�!PN���Gen=eB�rip���x�8��extt���Y�m�"�(� �HB���)��x�������Ȣ�r�es.�yA�ɠn@����*���p�@xM�_�NĀ6L�p��Ș�yAvL�0Xr�Ȉ2��"R;�Ƚ�\ra��	P�� h86��Gu+ʸ�φ��SeLɨm�9�69�P�Ȩr�Ȩ2�ɹ1&��n2�h� �0L�,XR}�RI{�e� L�x���c�Ș���N��vx�L��"��2\r@�]�N�82�d����b�ɉa��y1��/�kp�@���A��ruk��� L�sop��H�}�Cts{�����s�ʼ9��j965��S�c��h��5 J9��{�
�PL�J	e;en��t I[
x��com��Fh�L�4c J��fo��DIF+�6�Q���ڏrati|��p��1L�0�
R8l߾�M�����P��8� �j�mK�X�HZ�����N�oڠ��3̹q��vi���80�~�l Sl�yQ�F�tpk�xb�j� .�@�R�d������,/n(�8�8�0���
�:�O8�<�Q}�COt���PT��O (��.�Xp|�~H���?�ov �wv���8�22�pm���722��j7�^�@�̙���cf�=Yvr���vcu���O��O�O�O_#_5_7�3�Y_��wv4{_�_yw�ʈ�ust_�_�cus�_�Z��o�o,o>oPo�io��n�ge��(pLy747��jWelʨHM47ZKEq {���[�m�MFH�?�(ws K�8J�n���oΝ�fhl;��wm�f���? :�}(4�	<g J{��II�)̏މw��X�7714kﭏ/7ntˏ݊�e+���se�/�a!w��8�ɐ��EX \��!+: �p��~�002��nh�,:Mo+�xO���1 "K�O��\a��#0��.8���{�h�L?�j+�mond�:��t�/�st�?-�w�:���)�;��p(=h�;
d Pۻ��{:  ���� �J0��re�����STD�!t�reLANG����81�\tqd��������rch�.������ht�wv�WWָ� wR79��"Lo�51 (�I�W�h�8Ո�4�aww�� �vy �623�c�h a?�cti �֘!�X�iؠ�	t ��n,�։�����j��"AJ1P@�3p�vr{�H��6��!��- Se�T� E3�) G�J9�34��LoW�4 (S������ <����91 ��8!4�j9 �所+���y�
��	�btN�ite{�R  ��I@Ո�����P� ������	 ����Z�vol��X ��9�<�I�p���ld*���F�864{��?��K�	�k扐�֘1�/wmsk��M�q�Xa�e����rp��0RBT�1�ks.OPT�N�qf�U$ RTCamT��y��U ��y��U��UlU6L�T�1Tx����"SFq�Ue�6T���USP W�b DT�qT2h�T�!�/&+��TX�U\j6&�U U�UsfdO&�&ȁT����662DPN�bi��%�Q�%62V��$���%�� ��#(�(6To6e #St�%��#5y�$\�)5(To�%tT0�%5�W6T���%�#�#orc��#I���#���%cct�6ؑ?��4\W6965"8p6}"�#\j536�p��4�"�?kruO O,Im?Np�C �?�t�0<O�;�e ��%���?
;gcJ7 �"AV�?�;avs�f�O__&_8Wtp�D_V_0GT�F|_:Uc�K6�_�_r�O�3e\�s�O2^y`O:�miugxGvgW! m�%��!�%T�$E A`{6�po6��#37N��)5R5_2E���$0\���$Ada�Vd�Ѐ�V�?;Tz7�_�e7DCDTF9���#8�`��%��4y�te�d Z@�A}�@�}�0�4N�}�}���}�d�c& }����u 6��v��v1�u1\b��u$2}���}� R8�3�u�"}��"}�vaClg���Nrh�&�8�J�Y�o�ue���� j70�v=1��M{IG�uerfa��{q���E�N�ء���EYE�ce A ���񁏯pV�e�A!�� �2Յ�Q�%��u1�e�i�@��H�e����J0�� '��b��T��E In�B�  W�|��537g�����(MI�t�Ԇr��ݟ�am���n�ҵv!g�U -�v J�߆8⹖F���P�y�a�c���2���Rɏ j�o��2�� djdx�8r}� og\k��0��g��wmf��Fro/� Eqx'�4"}�3 J8��oni[��ᅩ}Ĵ�� o� ��ʛ���m@�R�e��{n�Д�V�o�������  �������"POS\����ͯ menϖ�⑥OMo�43��� �w(Coc� An[�0t���"e�a\�vp�z��.��cflx$�le��8�hr�trᅻNT� CF+�x E/�t	qi�M�ӓcxc��p�f�lx��,��Z�cx��
0 h�6��h8��mo��=�c H���)� (�vSER,���g�0߆0\r�vX�= ���I � - �tiغ�H��VC�82�8�5��L"�RC���n G/���w�P��y�\v�vm " o�lϚ�x`��=e�ߠ-�R-3?�����x�vM [�AX/2�\)�S�rxl�v#�0氆h8߷=� RA�X�A�����9�H��E/Rצ����hN߶"RXk��F�v˦85��2L/�xNB885_�q�Ro��0iA��5\r�O�9�K��v����88���.�n "�v��88��8s�i ?�9  ��/�$�y O��MS"���&�9R� H74&�`�74�5�	p��p��yc�r0C�c�hP0� �j�-�a%?o��6D95�0R7trl��c;tlO�APC����j�ui"�L���  ]����^棆!�A���qH��&-^7�w��� ���616C�q�794h���� M�ƔI���99��(���$FEAT_A�DD ?	����Q%P  	�H._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����������& 8J\n���������TDE�MO fY   WM_ �������� //%/R/I/[/�// �/�/�/�/�/�/�/? !?N?E?W?�?{?�?�? �?�?�?�?�?OOJO AOSO�OwO�O�O�O�O �O�O�O__F_=_O_ |_s_�_�_�_�_�_�_ �_ooBo9oKoxooo �o�o�o�o�o�o�o >5Gtk}� �������:� 1�C�p�g�y������� ܏ӏ���	�6�-�?� l�c�u�������؟ϟ ����2�)�;�h�_� q�������ԯ˯ݯ�� �.�%�7�d�[�m��� ����пǿٿ���*� !�3�`�W�iϖύϟ� ����������&��/� \�S�eߒ߉ߛ��߿� ������"��+�X�O� a����������� ����'�T�K�]��� �������������� #PGY�}� ����� LCU�y��� ���/	//H/?/ Q/~/u/�/�/�/�/�/ �/???D?;?M?z? q?�?�?�?�?�?�?
O OO@O7OIOvOmOO �O�O�O�O�O_�O_ <_3_E_r_i_{_�_�_ �_�_�_o�_o8o/o Aonoeowo�o�o�o�o �o�o�o4+=j as������ ��0�'�9�f�]�o� ��������ɏ����� ,�#�5�b�Y�k����� ����ş����(�� 1�^�U�g��������� ������$��-�Z� Q�c������������ �� ��)�V�M�_� �σϕϯϹ������� ��%�R�I�[߈�� �߫ߵ��������� !�N�E�W��{��� �����������J� A�S���w��������� ����F=O |s������ B9Kxo ������/� />/5/G/t/k/}/�/ �/�/�/�/?�/?:? 1?C?p?g?y?�?�?�? �?�? O�?	O6O-O?O lOcOuO�O�O�O�O�O �O�O_2_)_;_h___ q_�_�_�_�_�_�_�_ o.o%o7odo[omo�o �o�o�o�o�o�o�o* !3`Wi��� �����&��/� \�S�e���������� ����"��+�X�O� a�{����������ߟ ���'�T�K�]�w� ���������ۯ�� �#�P�G�Y�s�}��� �����׿���� L�C�U�o�yϦϝϯ� �������	��H�?� Q�k�uߢߙ߫����� �����D�;�M�g� q����������
� ��@�7�I�c�m��� ������������ <3E_i��� ����8/ A[e����� ���/4/+/=/W/ a/�/�/�/�/�/�/�/ �/?0?'?9?S?]?�? �?�?�?�?�?�?�?�? ,O#O5OOOYO�O}O�O �O�O�O�O�O�O(__ 1_K_U_�_y_�_�_�_ �_�_�_�_$oo-oGo Qo~ouo�o�o�o�o�o �o�o )CMz q������� ��%�?�I�v�m�� �������ُ���>;�  2�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s��������'9  :>Ugy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������/=C6Yk }������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ������/�A��$FEA�T_DEMOIN�  E��q���>�Y�INDEX�f�u��Y�ILE�COMP gw�����t��T���SETUP2� h������  N ܑ��_�AP2BCK 1�i��  �)�B���%�C�>� ��1�n�E����)��� M�˯�������<�N� ݯr������7�̿[� �ϑ�&ϵ�J�ٿW� ��Ϥ�3�����i��� ��"�4���X���|ߎ� ߲�A���e����� 0��T�f��ߊ��� ��O���s�����>� ��b���o���'���K� ��������:L�� p����5�Y� }�$�H�l~ �1��g��  /2/�V/�z/	/�/ �/?/�/c/�/
?�/.? �/R?d?�/�??�?�? M?�?q?O�?O<O����P� 2��*.VRCO�O�0*�O�O�3�O�O�5w@�PC�O_�0FR6:�O=^�Oa_�KT���_�_&U�_�\h�xR_�_�6*.FzODo�1	(SoEl�_<io�[STM �b�oН^+P�o�m�0i�Pendant �Panel�o�[H �o �g�oYor�ZGIF|��e�O8a��ZJPG �*���e���z��JJS������0@���X�%�
JavaScrgiptُ�CSʏ�1��f�ۏ %C�ascading� Style S�heets]��0
�ARGNAME.SDT���<�`\���^���Д៍�АDISP*ן���`$��d��V�e��CLLB.ZI��=�/`K:\��\�����Collabo����	PANEL1[�C�%�`,�l��o�o�2a�ǿV���r����$�3�K�V�9���ϝ�$�4i���V���zό�!ߘ�TPEINS.XML(��@�:\<����Cu�stom Too�lbar}��PA?SSWORD���>?FRS:\���� %Passw�ord Config��?J���C�� "O��3�����i���� "�4���X���|��� ��A���e�����0 ��Tf����� O�s��>� b�[�'�K� ��/�:/L/�p/ ��/#/5/�/Y/�/}/ �/$?�/H?�/l?~?? �?1?�?�?g?�?�? O �?�?VO�?zO	OsO�O ?O�OcO�O
_�O._�O R_d_�O�__�_;_M_ �_q_o�_�_<o�_`o �_�o�o%o�oIo�o�o o�o8�o�on�o �!��W�{� "��F��j�|���� /�ďS�e�������� �T��x������=� ҟa������,���P� ߟ񟆯���9���� o����(�:�ɯ^�� ����#���G�ܿk�}� ϡ�6�ſ/�l����� ϴ���U���y�� � ��D���h���	ߞ�-߀��Q߻��߇��,���$FILE_DG�BCK 1i������� ( �)
S�UMMARY.DyG,���MD:`������Diag� Summary����
CONSLOG��y����$����Console� log%���	T�PACCN��%�g�����TP A�ccountin�F���FR6:I�PKDMP.ZI	P����
��)�����Exceptio�n-����MEMCHECK������8�Memory� Data��L�N�)�RIP�E���0�%�� Packe�t LE���$S<n�STAT*|#� %L?Status�i	FTP�/�/��:�mment� TBD=/� >�)ETHERNE�/o�/�/��EthernU~<�figuraL���'!DCSVRF�1//)/B?�0 �verify a�llE?�M(5DIFF:? ?2?x�?F\8diff�?�}7o0CHGD1p�?�?�?LO �?,sO~3&�
I2BO)O;O�O bO�O�O�GD3�O�O�OT_� �O{_
VUP?DATES.�P�_~��FRS:\�_��]��Updates List�_���PSRBWLD'.CMo���Ro��_9�PS_ROB�OWEL^/�/:G�IG��o>_�o��GigE ��no�sticW�N��>�)�aHAD�OW�o�o�ob��Shadow C�hange��� 8+"rNOTI�?=O��Notific�"���O�A�PMIO�o��h��f/��on�^U�*�UI3�0E�W��{�UI������B���f��_��� ����O��������� >�P�ߟt������9� ί]�򯁯�(���L� ۯp������5�ʿܿ k� Ϗ�$�6�ſZ�� ~��wϴ�C���g��� ߝ�2���V�h��ό� ߰���Q���u�
�� �@���d��߈��)� ��M���������<� N���r����%����� [����&��J�� n��3��i ��"�X�| ��A�e�/ �0/�T/f/��//�/=/�/�/�$�$FoILE_�PPR�P���� �����(MDO?NLY 1i5� ? 
 �z/Q? �/u?�/�?�?t/�?^? �?O�?)O�?MO_O�? �OO�O�OHO�OlO_ �O_7_�O[_�O_�_  _�_D_�_�_z_o�_ 3oEo�_io�_�oo�o �oRo�ovo�oA �oew�*�� `����&�O��*?VISBCK,81>;3*.VDV�����FR:\o�I�ON\DATA\�/��Vis�ion VD filȅ��&�<� J�4�n������3�ȟ W������"���F�՟ �|������m�֯e� �����0���T��x� �����=�ҿa�s�� ��,�>���b���� �ϼ�K���o��ߥπ:���^����ϔ��*M�R2_GRP 1�j;�C4 w B�}�	 71�������E�� E��  F@ F��5U������L����M��J�k�Lzp�JP��Fg�f�?�  S����9��Y9}�9���8j
�6��6�;���A�  ���BH���B���B���$�������������@UUU#����� Y�D�}�h����������������
C��_�CFG k;T M���]��NO :
�F0� � \�RM�_CHKTYP  0�}�000���OM_MI9N	x���50�X� SSBdl.5:0��b�x�Y���%TP_?DEF_OW0x��9�IRCOM���$GENO�VRD_DO*�62�THR* dz%d�_ENB�{ �RAVC��9mK�� ��՚�/3�/��/�/�� �M!OUW s��}��ؾ��8�g�;?�/7?�Y?[?  C��0�a���(7�?�<B�?B����2��*9�N SMTT#t[)��X��4�$HOSTC�d1ux��\�?�� MCx��;�zOx�  2�7.0�@1�O  e�O�O	__-_;Z �O^_p_�_�_�LN_HS�	anonymous�_�_�_oo1o yO��FhFk�O�_ �o�O�o�o�o�oJ_ '9K]�o�_� ����4o�Xojo G�~�o^�������ŏ �����1�T�� �y����������� ,�>�@�-�t�Q�c�u� ��������ϯ��� (�^��M�_�q����� ܟ� �ݿ��H�%� 7�I�[Ϣ�ϑϣϵ� ���l�2��!�3�E� Wߞ���¿Կ����
� ������/�v�S�e� w����������� ��+�r߄ߖ�s��� ���߻���������� '9K]����� ����4�F�X�j� l>��}���� ��//1/T� �y/�/�/�/�/.D\A�ENT 1v
;� P!J/?  ��/3?"?W??{? >?�?b?�?�?�?�?�? O�?AOOeO(O�OLO ^O�O�O�O�O_�O+_ �O _a_$_�_H_�_l_ �_�_�_o�_'o�_Ko ooo2o{oVo�o�o�o �o�o�o5�oY�.�R�v��z?QUICC0���3��t14��"�����t2��`�r�ӏ!?ROUTERԏ���#�!PCJO�G$���!19�2.168.0.�10��sCAMP�RTt�P�!d�1m�����RT폟������$NAME �!�*!ROBO����S_CFG �1u�) ��Auto-s�tartedFTP&��=?/ ֯s����0�B�� f�x���������S�� ����,�������� �ϼ�ޯ��������� ʿ'�9�K�]�oߒ�� �߷��������� (:~�k�Ϗ��� ���������1�C� f���y����������� �,�>�R�?��c u��`����� (�$M_q� ����� /H %/7/I/[/m/4�/�/ �/�/�/�~/?!?3? E?W?i?����?�/ �?/�?OO/O�/�? eOwO�O�O�?�ORO�O �O__+_r?�?�?�? �O|_�?�_�_�_�_o �O'o9oKo]ooo�_o �o�o�o�o�o�oF_X_ j_~ok�_��� ���o���1�T U��y���������U��)�_ERR w�3�я�PDUSI�Z  g�^�p����>�WRD �?r�Cq�  �guest b�Q�c�u�������"��SCDMNGRPw 2xr�����Cqg�\�b�K�� 	P01.�00 8(q  � �5p�5pz�}5pB  �{� ���H����L��L��L�����O8�����l������a4� x��jȤ�x��8���\�U��)�`�;��#�����d�.��@�R�ɛ_GROU�ېy�����	�ӑ���QUPD � ?u����İT�Yg����TT�P_AUTH 1�z�� <!i?Pendan��-��l���!KAREL:*-�6�H͇KC]�m��U��VISION SET���ϴ�g�G�U� �����R�0��H�B߀��f�x��ߜ߮���C?TRL {�����g�
S�FF�F9E3��AtF�RS:DEFAU�LT;�FAN�UC Web Server;�)�� ��9�K��ܭ����������߄WR_CONFIG |ߛ� ;��IDL_CPU_PCZ��g�B�Dpy� BH_�MINj�)�}�?GNR_IO���g���a�NPT_SOIM_D_������STAL_SCR�N�� ���TPM?ODNTOL������RTY��y����F �ENO���Ѳ]�OLNK 1}��M�������|�eMASTE���ɾeSLAVE �~��c�O_CcFGٱBUO�|O@CYCLEn�>T�_ASG 19ߗ+�
 �� ��//+/=/O/a/�s/�/�/�/�/��N�UM��
@I�PCH�^RTRY_CNZ���@P�������� @kI�+E�z?E��a�P_MEMBE�RS 2�ߙ� 5$���2���ݰ7��?�9a�SDT_I�SOLC  �����$J23_D�SM+�3JOB�PROCN��JOmG��1�+�d8�?��+D�O�/?
�LQ�O __/_�OS_e_w_�_`�O Hm@��E#?>&BPOSREQO��?KANJI_����a[�MON ����b�yN_goyo@�o�o�o�Y�`3�<�� ��e�_ִ��_L����"?`EYLO�GGINLE��������$LANGUAGE ��<T� {q�LeGa2�	�b���g��xP��  �J�g�'��b����>�MC:\RSCH\00\<��XpN_DISP �+G�J��O�O߃gLOCp�Dz����AsOGBOOK �������������X����� Ϗ����a�*��	p�����!�m���!���=p_BUFoF 1�p���2F幟���՟D�� Collaborativǖ��� F�=�O�a�s������� ֯ͯ߯���B�9��K���DCS �>z� =���'�f���?ɿۿ���H@{�I�O 1�� ~?9ü��9�I�[�m� �ϑϣϵ��������� �!�3�E�Y�i�{ߍ�@�߱��������E��TMNd�_B�T�f� x������������ ��,�>�P�b�t���p����L��SEVD0���TYPN�1�$6���QRS�"0&��<2FL 1�"�J0���������GTP�:pOF�NGN�AM1D�mr�tUP�S�GI"5�aO5��_LOADN@G� %�%TI~�pZUZAUN#��(MAXUALR�M�'���(��_P�R"4F0d��1�B�_PNP� V 2��C	MDR�0771ߕ�B�L"8063%�@ ��_#?�ߒ|/�C��z�6��/���/�Po@P 2��+� �ɖ	T 	t  ��/�% W?B?{?�k?�?g?�? �?�?O�?*OONO`O CO�OoO�O�O�O�O�O _�O&_8__\_G_�_ �_u_�_�_�_�_�_o �_4ooXojoMo�oyo �o�o�o�o�o�o0 B%fQ�u�� ������>�)� b�M�����{������� �Տ��:�%�^�p��S�������D_L?DXDISApB��MEMO_AP�jE ?C
 �,�(�:�L�^��p������� 1�C ����4��������4��X���C�_MSTR ����w�SCD 1���L�ƿH��տ� ��2��/�h�Sό�w� �ϛ��Ͽ���
���.� �R�=�v�aߚ߅ߗ� �߻�������<�'� L�r�]������� �������8�#�\�G� ��k������������� ��"F1jUg ������� B-fQ�u����h�MKCFG� ����/�#LT�ARM_��7"0�0N/V$� �METPUᐒ3�ퟎ�ND� ADC�OLp%� {.CMN�T�/ �%� ����.E#>!�/4�%_POSCF�'�.�PRPM�/9ST�� 1��� 4@��<#�
1�5 �?�7{?�?�?�?�?�? �?)OOO_OAOSO�O wO�O�O�O�O_�A�!�SING_CHK�  �/$MODAQ,#����.;U�DEV 	��	�MC:o\HSI�ZEᝢ��;UTA�SK %��%$�12345678�9 �_�U9WTRI�G 1���l3%% ��9o��"ocoFo5#�V�YP�QNe��:SE�M_INF 1��3' `�)AT&FV0�E0po�m)�aE�0V1&A3&B�1&D2&S0&�C1S0=�m)GATZ�o;"tH? g�a[o�xA�� z���� �o>� �o'��K��� ����я:�L�3� p�#�5���Y�k�}�� ����$�[�H���~� 9�����Ưد������ ��ӟ�V�	�z����� ��c�Կ����
��.� ��d��)�;��Ͼ� q�������˿<��� `�G߄ߖ�IϺ�m�� �ϣ����8�J��n� !ߒ�M�������h_�NITOR� G �?�[   	�EXEC1�/�2*5�35�45�55��P�7�75�85�9� 0�Қ�4��@��L� ��X��d��p��|�������2��2���2��2��2��2���2��2��22*3��3��3@�;Q�R_GRP_SVw 1��k (�A��z�4�~�Kａ������K:z�j]�Q_�D��^�PL_N�AME !3%�,�!Defa�ult Pers�onality �(from FD�) �RR2� �1�L6(L�?�,0	l d �������� //(/:/L/^/p/�/��/�/�/�/�/�/ZX2 u?0?B?T?f?x?�?�?�?�?\R<?�?�? O O2ODOVOhOzO�O��O�OZZ`\RD�?�N
�O_\TP�O :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo _)_~o�o�o�o�o�o �o�o 2DVh z�[omo���� 
��.�@�R�d�v����������Џ� �Ef  Fb� �F7���   ��!��d��@� R�6�t������l�๟ʝ�����  ݘ����"�@�F�d����� "𩯹�ݐAG�  ϩU[�$�n�B�E� �� � @oD�  �?��� �?�@��A@�;�f��FH� ;�	}l,�	 |���j�s�d�>�� ��� K(���Kd$2K ���J7w�KY/J˷�ϜJ�	�xܿ�� @I���_f�@�z���f�γ�N�������	Xl��������S��ĽÔ��I �����5���  �����A?oi#��;���� o���l� �π��-���ܛG�G�Ѳ���@n�@a �  �  ���ܟ*�͵	'�� � H�I� �  �Р�n�:�Èl�È�=��̈́�в@�ߚЕ����/������̷NP� � ',���-�@�
�@���?�=�@A���B� � Cj�a�Be�C<i��#�Bи��ee��^^ȹBР��P����0̠�����ADz՟� n�3��C�i�@�R�RиY����  �@�7 ���  ���?�ff������n� ɠ#ѱy9�G
(���I�(�@uP@~����t�t���>�����;�Cd;���.<߈<�g�<F+<L�������,�d�,�̠�?fff?��?&�&��@��@x���@�N�@�?��@T�H�� ��!-�ȹ�|�� 
`�������/ /</'/`/r/]/�/��eF���/�/�/�/@m?��/J?�(E���G�#�� F Y�T?�?P?�?�?�?�? �?O�?/OO?OeOk� �O�IQOG�?�O1?��OmO_0_B_T_������A_�_	_�_P�_�_ o��A��An0 bФ/o C�_Uo�_�Op��؃o�o�ol�o���W�����o;C�E� q�H�d��؜a@q��e��F�BµWB]��NB2�(A����@�u\?��D�������b�0��|�uR�����
x~�ؽ���Bu*C���$�)`�$ ����GC#����rAU�����1�eG��D�I�mH��� I:�I��6[F���C��I��J�:�\IT�H
~�QF�y��p���*J�/ I8�Y�I��KFjʻCe�o��s��� ��Џ���ߏ�*�� N�9�r�]��������� ���۟���8�#�\� G�����}�����گů ���"���X�C�|� g�����Ŀ������ �	�B�-�f�Qϊ�u� ���ϫ��������,� �P�b�M߆�qߪߕ� �߹�������(��L� 7�p�[����������s($���3:�����$���3���d�,�4��x@�R�wa����l�<~�wa���e����wa4 �{����@��(L:ueP�	P~�A�O�������	���� G2W}h� �����/�� �O�O7/m/[(d=�s/ U/�/�/�/�/�/?�/�1??U?C?y?�=  �2 Ef9gFb-��77�9fB)aa�)`C9A`�&`w`@ -o�?w`e�O)O�?MO�Ow`�?�?�O�O�OD�O9c?�0�A7ht4�w`w`!w`xn
 �O9_K_]_ o_�_�_�_�_�_�_�_��_o#ozzQ ���h��G���$M�R_CABLE �2�h t�a�T� @@�0`�Ae��a�a�a��`ɺ�0�`C�`�aO8��tB�n�d���`�aE�4�GE�#�o�f�#���0��0�DO���By`��Š���bED4E��c,��o�g8 [ ���C�07�d�4
vے�0 ��b��XE��Z&�l�`y`
qCܛp�bHE�
v#=g�5D�Ү�qz
�lҠ`��0�q�p�bw0�
v�%c����b=%	E;h��u/o�c-��4tH� \�?�9�K�]�o�ԏϏ ��
�ɏۏ@���?��e o �e\��8�������6�0���� ����*�,�** \cOM ��ii��3��P% �%%� 2345678'901i�{� f������������1����
��`�n�ot sent �5���;�T�ESTFECSA?LGR  e�qiG��1d.�š
:��� �DCbS�Q�c�u���� 9UD1:�\mainten�ances.xm�l��ֿqY�DEFAULT-��i4\bGRP 2�M�  =��a�7�E�  �%For�ce�sor c?heck  ���b��z��p����h5-���ϻ��������%�!1st cle�aning of� cont. v��ilation��}�Rߗ+��[��Дߦ߸���me;ch�cal`������0��h5k�@�R�d�v����>(�rolle_Ƶ����/���(��:�L��Basi�c quarte�rly�������,������������M��:C@"GpP�a�b`i4�������#C���M"��{Pbt����Suppq�grease���?/&/8/J/\/���C+ ge��. batn�y`/��/h5	/�/�/�/? ?X_�ѷen'�v��/�/��/��?�?�?�?�?�G=?O�qEp"CrB1O��0�/ `OrO�O�O�O�t$��Lf��C-m��A�O:�OO$_6_H_Z_l_z�t*cabl�Om���S<m��Q�_:�
_�_�_oo0o@o)(Ӂ/�_�_���_��o�o�o�o�o�O�@hau1�l��2r xm�<qC:���op������R/eplaW�fUȼ2�:�._4�F�X�j�|�m�$%���ߟ�� ��#���
��.�@��� d���ŏ׏����П� ���U�*�y�����r� ��������	�q��?� ߯c�8�J�\�n���ϯ �����ڿ)����"� 4�Fϕ�jϹ�˿��� ���������[�0�� ��fߵϊߜ߮����� !���E�W�,�{�P�b� t����߼����� A��(�:�L�^���� ����������  $s�H������q� ����9]o �Vhz���U �#�G/./@/R/ d/��/�/��//�/ �/??*?y/N?�/�/ �?�/�?�?�?�?�??? Oc?u?JO�?nO�O�Op�O�O+J�r	 H�O �O__6M2_@OBE:_ p_>_P_�_�_�_�_�_  o�_�_oHoo(oZo �o^opo�o�o�o�o�op �o :z �bA�?�  @�q _���Fw��� �H* �** @q>v�p2T�f��x�:�������ҏ��eO^C7�Տ#�5�G� 	�k�}���ُ���c� ����W��C�U�g� ��ß)�����ӯ��� 	��-�w�����9��� ����m�Ͽ��=�O��E	A�$MR_HIST 2�>u}N�� 
 \
B�$ 2345678901^�f�#��]�9O���φϸ� O�)�;����q߃� ��L�^߬����ߦ�� ��7�I� �m�$��� Z���~������!��� E�W��{�2�����h������:�SKCFM�AP  >u�Q��r5��������ONREL  .�3���EXCFENB8q
��QFNCX�JJOGOVLI�M8dNá ��KE�Y8��_P�AN7����RU�N����SF?SPDTYPxC���SIGN8JTO1MOT�G���_CE_GRP 1�>uV��@ �����/Ⱥ� �/�/U//y/0/ n/�/f/�/�/�/	?�/ ???�/c??\?�?P? �?�?�?�?�?O)OO�MO,���QZ_ED�IT5 )TCO�M_CFG 1����[�O�O�O 
>�ASI �y3�!
__+[_O_ċ�>O�_bHT_/ARC_U.Ń	�T_MN_MOD�E5�	UAP�_CPL�_gNO�CHECK ?^�� �� o .o@oRodovo�o�o�o �o�o�o�o*!�NO_WAIT_�L4~GiNT�A���EUwT_ERMRs2���3��Ʊ J�����>_)�V�|MO�s��}x:O�v���8�?������ l��rPA�RAM�r�����j���5�5�G� = ��d�v�~�X� �����������֟�0����b�t������SUM_RSPACE�����Aѯۤ��$ODRDSP��S7cOFFSET_CARt@�_��DIS��PEN_FILE:�7�A�F�PTION_�IO��q�M_P�RG %��%$�*����M�WORK� �yf C��춍����������	 �Ћ����gT��RG�_DSBL  Ľ�C�{u��RI_ENTTO7 ��C� A �UT_SIM_Dy����V�LCT ��}{B �٭��_PEX�P=�ԷRAT�W dc|��UP ���
`���e�w�]ߛ�֩��$�2r�L6(L?���	l d����� �&�8�J�\�n��� ������������"�4�F�X���2�߈��� ����������*�<w�Tfx�� �����J`�ˣG���Tz�Pg��� ���/"/4/F/X/ j/|/�/�/�/���/ �/??0?B?T?f?x? �?�?�?�?�?�?�?�/ �/,O>OPObOtO�O�O �O�O�O�O�O__(_0:_��O��y_�]2ӆ��_�^�_�_�W�^]^]��/ooSog �Hgrohozo�o�o�o��o�oF`�#|`��A�  9y����O�K�1�!k��!����<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	O |�Q�s�r^�q>��u �s�F`H<zH~��H3k7GL��zHpG㎁99l7�k_B�T�F`C�4��k�H���t���-�Ae���k������s���  ��ሏ����EeBV�T���dZ���π���ڏ  ���q-�Fk�y�{Fb�U���n@6��  ����z�Fo��Be	'� �� ��I� ?�  �:p܋�=���ڟ웆�@���B�,���"B���g�AgN�����  '|���g��BU��p�BӀC׏�����@  #�yBu�&�ee�/^^މB:p2����>�m�6p�Z���Dz?o}�܏������׿@������Ǒ��� f�?  � �M���=*�?�ff�_8�J�ܿ 3pϑ�ñ�8�Чϵʖq.·�(����P���'��s�t�L�>��/�;�Cd�;��.<߈�<�g�<F+�<L ��^oiΚrd�@��r6p?fff?��?&�п�@���@x��@�N��@���@T����Z���ћtމ�u �߈w	�x��ti�>�)� b�M��q������� ������:�%�^��������W���S�E� � G�aF�� Fk���������1 U@yd��� ���q��	��{� A��h�����"a��ird��A{/@w/J/5/n/vA��aA���":t�/ C^/��/Z/ ލ?��`�/�/1??���W�����g��pE� ~1�?04�0
1�1�@IӀ��Bµ�WB]�NB2��(A��@�u�\?����������b�0�|�u�R����
�>��ؽ��B�u*C��$�)�`�? ����GC#����rAU�����1�eG���I��mH�� I:��I�6[F�﫹C4OI���J�:\IT��H
~QF�y��Ol@�*J��/ I8Y�I��KFjʻC�� -?�O�O__>_)_b_ M_�_�_�_�_�_�_�_ o�_(oo%o^oIo�o mo�o�o�o�o�o �o $H3lW�{ �������2� �V�h�S���w����� ԏ�������.��R� =�v�a�������П�� ��ߟ��<�'�`�K� ]���������ޯɯ�@�&�8�#�\��3(J�ϳ�3:a������J�3��c4�������������1�ǲ��ڿ��1����e���14 �{2�2�r�`ϖτϺϔ���%PR�P���! �h�!�K�6�o�Z�����u�|ߵߠ� ���������3��W� B�{�f�4���������d�A����!��1� 3�E�{�i��������������  2 E�f�7Fb�7�b�6B�!�!� C9� 	�� �0@�/`r� �����#x�� +=�3?, V*�8v��0�0�u�0�.
 D �����//%/ 7/I/[/m//�/�:�� ��ֻ�G����$PARAM_MENU ?2���  �DEFPU�LSE�+	WAITTMOUT�+�RCV? �SHELL_WR�K.$CUR_S�TYL� 4<OsPTJJ?PTB_?�Y2C/?R_DECSN 0�Ű<�?�?�? �?�?OO?O:OLO^O��O�O�O�O�O�!SS�REL_ID  �.����EUSE�_PROG %��*%�O0_�CCCR�0�B��#CW_HO�ST !�*!HT�_=ZT��O_�Sh_�zQ�S�_<[_TI�ME
2�FXU� GDEBUG�@�+�C�GINP_FLM3SKo5iTRDo5gWPGAb` %l��tkCHCo4hTYPE�,� �O�O�o #0Bkfx� �������� C�>�P�b��������� ӏΏ�����(�:��c�^�p�����7eWO�RD ?	�+
 �	RSc`���PNS��C4�J9Ov1��TE�P�COL�է�2��g�LP 3������OjTRACECToL 1�2��!� �� ��Қ�q�DT �Q�2�Ǡ��D� � :�����Ԡ� Ԡ��}�ׯ���;�4��4�� 4���;�u:�q:����;�8�	8�
8��8�8�8�8��8��@:�8�8�@��� ���ٱ޴���ؿ�$�6� ��
�l�~�@�R�dϞ� ����������
��V� h�zߌߞ߰������� ��
�,�>�P�*�<�v�܈�*� +8� (��)��*������ ����)�;�M�_�q� �������������� %,�>�P�b�t��� ���������С� *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6@u bt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� ��V�߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�?��?�?�1�$PGT�RACELEN � �1  ����0��6_�UP ���e�A@�1@��1_CFG ��E�3�1
@�
<D�0<DZO<C�0�uO$BDEFSPD� �/L�1�0���0H_CONF�IG �E�3� �0�0d�D�&�2 �1�APpDsAl�A�0��0IN'@?TRL �/MOA�8pEQPE�E��G�A<D�AIWLID(C�/M	bT�GRP 1ýI� l�1B � �����1A��33FC� F8� E�� @eN	�A�AsA�Y�Y�A�@?� 	 vO�Fg�_ ´8cokB;`baBo,o>oxobo��o�1>о�?B�/�o�o~�o =%<��
 C@yd��"�������  Dz@�I�@A0�q� � ������ˏ���ڏ� ��7�"�4�m�X���|����Ú)ґ
V7�.10beta1�HF @�����Aq��Q�  �?� �B���P�p �C��~&�B�EQA���Q�P�Q�� ß[�m����<CA��0�b�@p���f������ҡr�R�ܣ�Rљ����1�i�������t<B!CeQKNO?W_M  lE7F�bTSV ĽJ�BoC_�b�t��������������1�]aSM��SŽK ���	�NB�0����ĿK���-�bb��A�RP���`�0�Ŗ��bQMR�S��T�iN���d����V]ST�Q1 1=�K
 4MU�iǨj� K�]�oߠ� �ߥ߷�������2�� #�h�G�Y��}������
������,�2r7�I��1�<t�H��P3^�p�����,�A4��������,�5(:,�6Wi{�,�7����,��8�!3,�MA�D�6 F,�OV_LD  KD��xO.�PARNUM�  �MC/%�S+CH� E
9'!8G)�3Y%UPD/���E�/P�_CMP_0��0@�0'7E�$�ER_CHK�%05H�&�/�+RS����bQ_MO�+?=5_�'?O�_RES_G6��:�I�o�?�?�? �?O�?O7O*O[ONO OrO�O�O�{4]��<�?�Oz5���O__ |3 #_B_G_|3V b_ �_�_|3� �_�_�_|3 � �_�_o|3Oo>o<Co|2V 1�:�k1�!�@c?�=2T?HR_INRc0i!�}�o5d�fMASS6�o Z�gMN�o�c�MON_QUEUE �:�"�j0��UO�N� U1Nv�+DpENDFqd?`y�EXEo`u� BE�npPAsOPTIO�Mwm;DpPROGR�AM %$z%�Cp}o(/BrTASK�_I��~OCFG� �$��K�D�ATA��T���j12/ď֏��� ���+�=�O�a�����������͟��INFO�͘��3t��!� 3�E�W�i�{������� ïկ�����/�A�@S�e�w�����Θ�a '��FJ�a K_N���T��˶ENB�g ڽw1��2��G�N�2�ڻ P(O�=���]�ϸ�@���v� ��u�uɡdƷ_E?DIT �T���|��G�WERFL�x��c)�RGADJ {Ҷ�A�  $Ձ?j00��a�Dqձ���5�?�$�ʨ�<u�)%e��0����FӨ�2�R��+	H;pl�G�b_�u>�pAod�t$��*�/� **:�j0�$�@�5AY�T���^��q�� �b~�L��\�n��� ������������� 4�F�t�j�|������� ������bLB T�x����: ��$,�Pb ���/���� /~/(/:/h/^/p/�/ �/�/�/�/�/V? ?? @?6?H?�?l?~?�?�? �?.O�?�?OO O�O DOVO�OzO�O_�O�O �O�O�Or__._\_R_ d_�_�_�_�_�_�_�f	g�io�pWo�o{d� �o�~o�ozoB�PREF �R��p�p
�IOR�ITY�w[���M�PDSP�q��pwU�T6����ODUC-T3�����;OG��_TG��8���ʯrTOENT �1׶� (!?AF_INE�p,�~7�!tcp7�>_�!udN���?!icmv���֯rXYK�ض���q)� ,�����p��&�	��R�9� v�]�o�����П����@��*��N�`�*�s�K��9}�ߢ���Ư ,�/6쒯������خ�At�,  �Hp��P�b�t�����u�w�HANCE �R��:�w!d��连�2s�9Ks���PORT_N�UM�s�p����_CARTRE�P{p�Ω�SKST�A�w d�LGS6)�ݶ��tӁp�Unothin�g�������{��T?EMP ޾y���'e��_a_seiban�o\��ol� ��}߶ߡ��������� "���X�C�|�g�� ������������	� B�-�f�Q���u����� ��������,< bM�q��������(L�VOERSIyp�w}� disab�ledWSAVE� ߾z	26�00H768S?�!ؿ����/C 	5(�r)og+^/y�e{/�/�/�/�/�*�,/? �p���]_�p 1�Ћ� �����W�h?z?�W*pURGE«�B�p}vgu,�WFF�0DO�vƲ�vW%���4(�C�WRUP_�DELAY ��\κ5R_HOT �%Nf�q׿GO�5R_NORMAL&H��r6O�OZGSEMI�jO�O�O(qQSKI%PF3��W3x=_ 98_J_\_]�_�_{_ �_�_�_�_�_�_	o/o AoSoowoeo�o�o�o �o�o�o�o+= aOq����� ���'��7�]�K��������)E�$RAF{���K/�zĀÁ�_PARAM�A3���K @.�@�`�61�2C<��y��C�6$�B�ÀBTIF�4`�R�CVTMOUu�vc��ÀDCRF3}��I �+Q�;/�CC�Se�D�#�1=h�߶-0�t]�/{��ޅ�����1�0��_��k_����Cd;��.<�߈<�g�<F+<L���Ѱ��d�u�L����� ��ϯ����)�;��M�_���RDIO_TYPE  M=�U�k�EFPOS1w 1�\�
 x4/�����+�$/<� �$υ�pϩ�D���h� �ό��'������o� 
ߓ�.ߤ�Rߌ����� ��5���Y���i�� *�<�v���r����� ����U�@�y����8� ��\�����������?���c����2 1�KԿX�T�<x��3 1�����nY�S4 1�'9K�/��'/�S5 1� ���/�/�/�/:/S6 1�Q/c/u/�/-??Q?�/S7 1��/�/
?D?�?�?|�?d?S8 1�{?��?�?�?WOBO{O�?SMASK 1pL��O�D�GXNO���F&�^��MOTE�Z�Ż��Q_ǁ��%]pA݂��PL_R�ANG!Q]�_QOW_ER �ŵ�P�1VSM_DRYP_RG %ź%"O��_�UTART ��^�ZUME_P�RO�_�_4o��_E�XEC_ENB � J�e�GSPD�`O`WhՅjbTDB�ro�jRM�o�hIN�GVERSION7 Ź#o�)�I_AIRPUR�hP �O(�MMT�_�@T�P#_ÀO�BOT_ISOLEC�NTV@A'qhu/NAME�l��o�J�OB_ORD_N_UM ?�X#q�H768 � j1Zc@�r�
�rV�s���r�?�r?��r�pÀPC_T�IMEu�a�xÀS�232>R1��� LTEAC�H PENDANw�:GX�!O �Mainten�ance Con%sj2����"��No UseB� ׏������1�C�y��V�NPO�P@�YQ��cS�CH_�L`�%^ �	�ő��!UD1:�럒�R�@VAIL��q@�Ӏ�J�QSPACE1 2�ż ��YRs�i�@C�t�YRԀ'{��8�?��˯��� �"���7�2�c�u��� ��G���߯ѿ򿵿� (��u�AC�c�u��� ��Ͻ�߿���ϵ�� (��=�_�qσϕ�C� �������߱��$�� 9�[�m�ߑߣ�Q��� ���߭��� ���	�W� i�{���M������� 5���.S�e�w� ����I������� *?as�� E�����/&/ /;/]o���� ��/2/�/?"?�/7? Y/k/}/�/�/O?�/�/��?�?�?O0OOKA���*SYPpM*��8.30261� yB5/21/2�018 A �lWPfG|�H�_TX`�� !$COM�ME�$U�SAp $E�NABLEDԀ�$INN`QpIOR��B�@RY�E_SI�GN_�`�AP�AI�T�C�BWRK�BD�<�_TYP�CRINDXS�@W�@%V�FRI{�_GRP�Ԁ$UFRAM��rSRTOOL\VM�YHOL�A$L�ENGTH_VT�EBTIRST�T  $SECLP��XUFINV_P�OS�@$MA�RGI�A$WA3IT�`�ZX2�\�V[G2�GG1�AI�@��S�Q	g�`_WR�BN�O_USE_DI��BuQ_REQ�BC��C]S$CUR_�TCQP�R"a^f ��GP_STATU}S�A @ �A�3`�BLk�H$zc1��h�P@���@_�F�X �@E_M�LT_CT�CH_l�J�`CO�@OL�E:�CGQQ$W�@w��b#tDEADL�OCKuDELAY_CNT�a3qGt��a$wf 2+ R1[1$X<�U2[2�{3[3$Z wy�q%Y�y�q%V�@�cL�@�b$V�`�RV�U�V3oh>b�@ �� �d�0arMSKJ�LgWaZ�C`NRK�PS_RATE�0�$���S
`�Q�TAC��PRD���e��S*��a4�A�0�DG��A 0�P�flp3 bquS2ppI��#`
`�P 
�S�\`  �A�Ro_ENBQ ��$RUNNER�_AXI�<`ALPLx�Q�RU�THICQ?$FLIP7��D?TFEREN��R��IF_CHSU�I0W��%V)�G1�����$PřA�Q�Pݖ_�JF�PR_P�	��RV_DATA~�A  $��ETIM���$V�ALU$�	�OP_   ��A  2 ��SC*�	� ?�$ITP_!�SQ�]PNPOU}�o�TO�TL�o�DSP��J�OGLIb��PE_IPKpc�Of�i��P�X]PTAS�$KEPT_MIR��d¤"`M�b�APq�aE�@�y�q�g@١�c�q�PG�BRK�6�x���L�I�� � ?�SJ�q�P�ADyEz�ܠBSOCz��MOTNv�DUM�MY16Ӂ$S}V�`DE_OP���SFSPD_OViR
���@LD�����OR��TP8�L�E��F������OV���SF��F����bF��d�ƣ&c)�fQc�L�CHDLY��REGCOV���`��W�P1M��gŢ�RO����r��_F�?� @v�=S �NVER�@�`�OFS�PC,�CSWDٱc�ձ���B�����TRG�š�`E_�FDO��MB_CiM}���B��BLQ��¢	�Q�̄Vza�BU�P�g��G
��A�M���@`KՊ�e�_M!�d�AMf�Q��OT$CA����DF���HBKd�v���+IOU��I'R��PA����������p���і�DVC_DB �S!�x�Q�!�s�d�9�1A��9�3A��ATIO�0��͠��aUS����WaAB�� R+c�`tá`DؾA���_AUXw�SUB'CPUP���S�`�����3Եжc���3�F�LA�B�HW_C wp"�Ns&�]sAa���$UNITS�|M�F�ATTRIz��Z�CYCL�CN�ECA���FLT�R_2_FI��TARTUPJp��ь�A��LP������_�SCT*cF_F�F1_P���b�FS��+�K�CHA/Q��*�d�RSD��Q��ص�Q���_TH�PRqOr���հEMPJ�䢠G�T� ��Q�DI�@y�R�AILAC/�bM�X�LOf�xS��ځ`���拁���PR#�S`app�C� �	��FUNC���RIN`QQP�� ԱRA)]R ���AƠ��AWAR֓��BLZaWraAkg�ngDAQ�0B�rkLD�र�&q�M�K���TaI���j��$�@�RIA_SW��AF��Pñ#��%%p�p9r1��MOIQ����DF_~P(�PD�"LM-�FA�PHwRDY�DORG��H; _QP�s%MU�LSE~Pz���*��� J��Jײ��F�AN_ALMLV�G��!WRN�%HA#RDP��UcO�� �K2$SHADO�W]�kp�a02��� S�TOf�+�_^�w�A�U{`R��eP_SBR�z5���:F��| �3MPINF?��\�4��3REGLV/1DG�+cVm L�C�CFL(��?��DAiP���Z`�� q�����Z�	 �Pv(Q$�A$Z�Q� V�@�[�
� ��EG��o���kA#AR���㌵2�axGܘ�AXE��RO]B��RED��W�Q2D�_�Mh�SYA��AtF��FS�GWRI�P~F&�STR����E��˰EH�)��D�a�\2kPB6P��=V��D.v�OTO�1)���ARYL�tR�v�3�淡FI&�ͣ$LGINKb!\��Q��_3S���E��QX�YZ2�Z5�VOFIF���R�R�XxP	B��ds�G�cFI�03g�������_J��'�ɲ �S&qR0LTV[6���a#TBja�"�bC����DU�F7�TU�R� X��e�Q�2XP�ЊgFL�E���x@�`�U9Z8���� W1	)�K��Mw���F9��劂����OCRQj��G;W3�� �#�Ґd ���uz�����1�tOVE�q_�M ��ё?C�uEC�uKB�v '0�x-�wH��t� ��& `��qڠ�B�ё �u�q�wh�ECh����SER��K	�EPH����AT�K�6e�9e�W���AX s�'��v�/�R �� ��!�� ��P��`���`�3p�Yp�1 �p�� �� �� (� � 8�� H�� X�� h��� x�� ������DEBU�$%3�I��·RAB���ٱr�sV��� 
d� J、��@񘧕���� ���Q���a���a��3q���Yq+$�`%"<�cL�AB0b�u�'�G�RO���b<��B_s��"Tҳ*`�0A��u��uq�p1}�AND Gp�������U��p1�� �ѷ0�Qθuݸ���PNT0���SE�RVE �Z@ $�`EAV�!�PO����nP!�P@��$!Y@  ]$>�TRQ�b
=�d�BG�K�%"2\���� _  l8��5�D6ERRVb(��I��V0`;���TO	Q:�7�L�@
�R��Je G�%�Q�� <�50F� ,�`�z��>�RA� 2' d!�����S�  M��pxU �����OCuG� � ��COUNT�6Q��FZN_CFGF� 4#��6��TG4�_�=�����ü��VC ���M  �"��$6��q ��CFA E� &��X�@@�������A���r�AP��P@HEL�0~�� 5b`�B_BAS��RS)R�6�CSH��R��1�Ǌ�2��3��U4��5��6��7��98��}�ROO���̚P�PNLEA�cAB�)ë ��ACKu�IeNO�T��(B$UR08� =�_PU��!0��OU+�Pd�8j���� V��TPFWD_KAR��� ��RE(ĉ P�P�>7QUE�:RO�p�`r0P1I� x�j�Pp�f��6�QSEM���0��� A��STYfL�SO j�DIX��&�����S!_TM>CMANRQ��P�ENDIt$KEYSWITCH��ذ�kHE�`BE�ATM83PE{@L�E��>]��U��F���SpDO_H�OM# O�@�EF�pPRaB�A#PY��C� O�!���OV�_M|b<0 IOCqM�dFQ��h�;HKYA D�Q�7��UF2��M���p޸cFORC�3WA�R�"�OM|@ G @S�#o0U)SUP�@1�2&3&�4E���T�O��L����8UNLO�v�D4K$EDU1 � �SY�HDD�NF� M�BL�OB  p�S�NPX_AS��� 0@�0��81$�SIZ�1$VA�{���MULTIP�-��# A� � $��� /$4`�BS��0�C���&OFRIFBO�S����3� NF�ODBUP߰�%@3;9(Ÿ)"��Z@ x��S�I��TEs�r�cSKGL�1T�Rp&���3B��@�0STMTdq�3Pg@VBW�p��4SHOW�5@��SV��_G�� 3p$PCJ�PИ���kFB�PHSP 1AW�EP@VD�0WC�� ���A00��PB XG XG �XG$ XG5VI6VI7�VI8VI9VIAVIB�VI�XG�YF�0XGFPVH��XbI1oI1|IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1Y1YU2UI2bI2oI2|I2�I2�I�`�X�I2pT�X�I2�I2�I2�I2�I2Y2Y�p�h�bI3oI3|I3�I3��I3�I3�I3�I3��I3�I3�I3�I3��I3Y3Y4�i4�bI4oI4|I4�I4��I4�I4�I4�I4��I4�I4�I4�I4��I4Y4Y5�i5�bI5oI5|I5�I5��I5�I5�I5�I5��I5�I5�I5�I5��I5Y5Y6�i6�bI6oI6|I6�I6��I6�I6�I6�I6��I6�I6�I6�I6��I6Y6Y7�i7�bI7oI7|I7�I7��I7�I7�I7�I7��I7�I7�I7�I7��I7Y7TɁV5P� UD�y"ՠ���
<A62��:t�R��CMD� ���M5�Rv�]��Q_h�R���e����<��YSL���  � �%\2��+4�'�W�BVALU���b��'���FH�IgD_L���HI��9I���LE_���f��$0C�SACѿ! h �V?E_BLCK���|�1%�D_CPU5� � 5ɛ �����C�� ���R " � �PWj��#0��LA�1SBћì���RUN_FLG�� �����ĳ ��������B��H���ХĻ��TBC2��# � @ B��e �S�p8=�FTDC�����V���3d�Q�T!HF�����R�L�?ESERVE9��F��3�2�E��Н��X -$��LE�N9��F��f�RA���W"G�W_5�b�14��д2�MO-�T%	S60U�Ik�0�ܱF����[�DEk�21LgACEi0�CCS#0�� _MA� j��z��TCV����z�T�������.Bi�'AH�z�'AJh�#EM5�"��J��@@i�V�z���2Q �0&@o�h�6��JK��VK9��0{���щ�J0�����JJ��JJ��AAAL���������4��5�ӕ N1����딨�.�LD�_�1�* �CF�"% `�GROU���1��AN4�C�#m RE�QUIR��EBqU�#��6�$Tk�2$���zя #��& \�APPR� C� 0�
$OP{EN�CLOS"�St��	i�
��&' �MfЩ����W"-_MG�7C�B@�A���BBR=K@NOLD@�0RTMO_5ӆp1J��P�������������60��1�@ )!�>#�(� ������'��+#PATH''@!6#@!�<#� r� '��1SCA�؆�6IN��UChJ�[1� C0@UM�(Y ��#�"�����*����*��� PAYLO�A~J2LؠR_AN^�3L��91��)1AR_F2L3SHg2B4LO4�!�F7�#T7�#ACRL�_�%�0�'�$��H���.�$HA�2FWLEX��J!�) P�2�D߽߫����0��* : ����z�FG]D����z���%�F1]A�E�G�4�F�X�j�|���BE ������������ (��X�T*�A���@�X I�[�m�\At�T$g�QX<�=��2TX���e mX��������������@����+	�J>+ �-�K]o|��٠AT�F�4�ELPFPѪs�J� *� ;JEmCTR�!�A�TN�vzHAN/D_VB.��1��n$, $8`F2Av���SWu	#-� $$M*0 .�]W�lg��PZ����A��� 1�����:AK��]AkA�z��LN�]DkD�zPZ G��C�ST�_K�lK�N}DY ��� A����0��<7 ]A<7W1�'��d�@g`�P��������"EX1B$. M�2D%"��H����OASYMj%0�� Bj&-��-W1�/_� {8� �$�����/�/�/�/ 3J<�:9��/�89�D_VI��v����V_UNI�ӛ��cD1J����� ��W<��n5Ŵ�w=4�@�9��?�?<�uc�4��3��%�H���a/�j��0�DIz�uO�ĭ�k�>S0 �`��I��A� �#���@ģ���@���IPl� 1 � -/�ME.Qp��49�ơT}�PT�;pG �+ Gt� ����'��T�0 $DUMMY1���$PS_�@RF��@  G b�'FLA@ YP(c|��$GLB_TP� ŗ���9 P�q���2 X� z!ST�9�� SBRM M�21_V�T$S/V_ER*0O�p�Ӧ��CL����AGPOl��f�GL~�EW>��3 4H �$Y
rZrW@�x�A1+��A���"j� �U&�4� 8`NZ�"�$�GI�p}$&� �-� �Y�>�5 L�H {��}$F�E^��NEAR(PN�CyF��%PTANC�B�	!JOG�@� �6.@$JOIN�Twa?pd�MSET.>�7  x�E��HQ�tpS{r��up>�8׼ �pU.Q?��� LOCK_FOxV06���BGLV�s�GLt�TEST_sXM� 3�EMP�����_�$U&@%�w`24� Y��5��2�d��3��C�E- ���� $KA�R�QM��TPDRqA)�����VECn@���IU��6��H=Ef�TOOL�C2�V�DRE IS3�ER6��@ACH� 7?Ox �Q��29Z�H I� � @$RAIL_�BOXEwa�R�OBO��?��HOWWAR�1�_�zROLMj��:q�w�jq� �@ O_=Fkp! d�l�>�9�� �R OB8B: �@�	"�"�OU�;�Һ�3�ơ�r�q_�$PIP��N&`H�l�@���#@CORDE�Dd�p >Cf�fpO��� < D ��OB⁴sd����Kӕ���qSYS��ADR�qf��T�CHt� = ,�8`ENo��1Ak�_�{�-$Cq_�f�VW�VA��> � � &��PREV�_RT�$ED�ITr&VSHWRBkq�֑ &R:�v��D��JA�$�a$HEAD�6�� ��z#KE:�E�CPwSPD�&JMP��L~��0R*P��?���1%&I��S�rC��pNE; �q�wTISCK�C��M�1<��3HN��@ @p� 1Gu�!_GPp6���0STY'"xL�O��:�2l2?�A �t 
m G3%%$�R!{�=��S�`!�$��w`���ճ���Pˠp6SQU��E�Ҟu�TERC�Q2�{TSUtB �����hw&`gw�Q)�pO����@IZ��{��^�PR�kюB1�XPU���E_DO���, XS�K~�A�XI�@���UR �pGS�r� ^0�&��pY_) �ET�BPm��o��0Fo��0A|���Rԍ��a�;�SR�Cl>@P��b_�yUr��Y ��yU��yS��yS���U Ї�U���U���U�]���Ul[��Y�bXk�]C�m�����YRSC��� D h�D1S~0��Q�SP���eATހ���A]0,2~N�ADDRES<=B} SHIF{s��_2CH�p�I\��=q�TVsrI��AE"���a�Ce�
���
;�VW�A��F 	\��q��0l|\A@�rC�_B"R{zp����q�TXSCRE�E�Gv��1TICNA���t{�c�8�A�b?�H T1�� �B�����I��A��BE�y RRO������� B���T�UE�4I �g�!p�S���RSM]0�GU�NEX(@~Ƴ�j�S_S�ӆ��Á։񇣣��ACY�0� 2-H�pUE;�J���\��@GMT��Lֱ��A��O	�BBL�_| W8���K �Լ0s�OM��LE�/r��� TO!�s�RwIGH��BRD
�%qCKGR8л�T�EX�@����WIDTH�� �B[�|�<� �UI_��H>i� L 8K���!_�!=r���R:�_� ��Y�1�O6q�%Mg0紐U��h�9Rm��LUMh��F�pERVw��P����`�N��&�G�EUR��FP)�)&� LP��(RE%@�a)ק�a�!��f �U5�6�7�8Ǣ�#B�É@���tP�f�W�S@M�US=R&�O <����qU�Qs�FOC).��PRI;Qm� :�޹�TRIP�m��UN����Pv� �0��f%��'���@�0� Q����AG ��0T� �a>q�O	S�%�RPo���8�R/�A�H�L4N���U¡�SU�g��8¢5��OFF����T�}�O�� �1R�����S�G�UN��6�B_�SUB?���,�SR	TN�`TUg2��mCsOR| D�RAUrP�E�TZ�#'�VCCܵ�	3V AC3�6MFB1�%d�P=G �W (#��ASTEM����䦒0PE��T3G�X� �\ ��MOVEz�A��AN�� ����M���LIM_X ��2��2��7�,���`��ı�
�BVF�` E���~��04Y���IB�7���5S��_�Rp� 2��� WİGp+@��}СP|��3�Zx ���3���A�ݠ9CZ�DRID��B��Vy08�90� De�?MY_UBYd�� �6��@��!��X���P_S��3��L��KBM,�$+0DEY(#EX`�����_UM_MU� X����ȀUS�� ���=G0`PACI���� �@��:��:,�:�����RE/�3qL�+���:[��TAREG��P�r��R<�\ d`��A��$�i	��AR��SW2 $��-��@Oz�%qQA7p�yREU�U�0�1�,�HK�2]g0�qP� N� �sEAM0GWOR����MRCV3�^� ���O�0M�C��s	���|�REF_���x(�+T�  ���������3_RCH4(a�P �І�hrj�NA����0�_ ��2����L@��n�@@OU~7w6d���Z��a2[��cRE�p�@;0\�ct�a'2K�@SUL��e]��C��0�^��� NT��L�3��(6 I�(6q�(3� L��Q5���Q5I�]7q�}�T�g`4D`�0.`0�A�P_HUC�5SA.��CMPz�F�6�5�5�0_�aR��a�1�I\!X�9��GFS���ad ��M8��0p�UF_x��B� �ʼ,RO��Q��'l����UR�3GR�`.�3IDp���)��D�;��A��~�IN"��H{D���V@AJ���S͓UWmi`=�����TYLO*��5����bt� +�cPA� �cCACH�vR�U@vQ��Y��p�#CF�-I0sFR�XT���VNn+$HO����P !A3�XBf�(1 ����$�`VPy� ^b_'SZ313he6K3he12J�eh chG�ch�WA�UMP�j��IkMG9uPAD�i�iIMRE�$�b_SIZ�$P����0 ���ASYNBUF��VRTD)u5tq~ΓOLE_2DJ�(Qu5R��C��U��vPyQuECCUl�VEMV �U�r�WV�IRC�aIuVTP G���rv1s��5qMP#LAqa��v�V0��c��� CKLA�S�	�Q�"��d ! �ѧ%ӑӠ@}¾�q$�Q���Ue |�0!�rSr�T�#0! ���r�iI��m�vK�BG��VE�Z�P�K= �v�Q�&�_H�O�0��f � �>֦3�@Sp�SLO�W>�RO��AC�CE���!� 9�VR`�#���p:���AD������PAV�j�� D:����M_B"���N^�JMPG ��g:�>#E$SSC��F��vPq��hݲvQS��`qVN��LEX�c�i T`�sӂ�ܗQ�FLD �DEsFI�3�02����:��VP2�Vj'� �A��V�4[`MV_PIs��t`���A�@��FI��|�Z��Ȥ�����A����A��~�GAߥ1 LsOO��1 JCB�इXc��^`�#PLA!NE��R��1F�c�����pr�M� [`������S����f����A@f��R�Aw�״tU�΁pRKE��d�VA�NC�A���� �k���ϲ�BR_AA� l��2� �p�p�#Hć�m h����O K�$������kLЍ0OU&A�"A�Y
p�pSK�TM@F�VIEM 2l p��P=���n <<�x�dK�UMMYK1�P��`D�M�ACU��#AU���o $��TIT>�$PR�����OP���VSH�IF�r�p`�J�Qsԙ�fOxE$� _R�`U�#���� s��q������G�"�G�޵'�T�$�SC9O{D7�CNTQ i� l�>a�-�a�;�a�H�@a�V���1�+�2u1���D����  ]� SMO�Uq�d�a�JQ�����aI_�R[�r�n�*@�LIQ�AA/`�XV%R��s�n�TL���oZABC�t��t�c�
|!ZIP���u���LVbcL�n"�� r�MPCF�x�v:�$�� �~��DMY_LN��p�����@y�w Ђ�(a�u� MCM�@C>bcCART_�D�PN� $J71D��=NGg08Sg0�BUXW� ��UXEUL|ByX���	��zAZ��x 	����m�YH�Db  �y 80���0EgIGH�3n�?(� �H����$z ����|�����$B� K�d'��_��L3�RV�S�F`���OVC �2'�$|�>P&���
q���5D�TR�@ �V�1�SPHX��!{ ,� *�<�$R�B2 2� ���C!��  ��| V+@b*c%g!�`+g"�`V*�,8�?�V+�/V.��/�/?�/�/V(7%3 @/R/d/v/�/6?�/�/ �?�?�?O4OOION;4]?o?�?�?�?SO�? �?�O_�O0_Q_8_f_N;5zO�O�O�O�Op_ �O_o8o�_MonoUo�oN;6�_�_�_�_�_ �oo%o4Uj�r�N;7�o�o�o�o �o� BQ�r�5���������N;8��� ��Ǐ=�_�n���R�टş��ڟN;G �� џ�
����?���W�i�{� ������ï�.��� ����A��dW�<� N�|�������Ŀֿ� ޯ���0�B�_�R� d�꿤϶��������� ����*�L�^��r� ��
�������������&�8�J�l�~� `ҟ @W��� ��ߩ��-���� &�,���9�{����� a��������������� A'Y��� �������a#1�
��N;_MODE  �^�S ��[�Y�B���
/\/*�	|/�/R4CWOR�K_AD�	�%�LT1R  ����� �/� _INT�VAL�+$��R_OPTION6� �q@V_D�ATA_GRP �27���D��P �/~?�/�?�9��?�? �?�?OO;O)OKOMO _O�O�O�O�O�O�O_ �O_7_%_[_I__m_ �_�_�_�_�_�_�_!o oEo3oioWoyo�o�o �o�o�o�o�o /eS�w��� ����+��O�=� s�a�������͏��� ߏ��9�'�I�o�]������$SAF_DO_PULS� ��~������CAN�_TIM�����ΑR !��!Ƙ�W�5�;#U!P"�1!��� �?E�W�i�{��� ��.�ïկ�����V'(~�T"2F�D��dR�I�Y��2�o+@a얿����)��u��� k0ϴ��w_ ��  T� �� �2�D�)�T D��Q�zόϞϰ� ��������
��.�@� R�d�v߈ߚ�/V凷�����߽�|�R�;�o ��W�p��
�t��Diz$� �0 � �T"1!� ���������� ������*�<�N�`� r��������������� &8J\n� ������� "4FX ��࿁ �������/ `4�=/O/a/s/�/�/��/�/�/�/�!!/ �0 ޲k�ݵu�0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ ok$o6o HoZolo~o�o�o�o�o 1/�o�o 2DV hz�/5?���� ����&�8�J�\� n���������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u��� ���`Ò�ϯ�� ��)�;�M�_�q����������˿ݿ� �p���3� ���&2�,��	123�45678v�h!B!���`Ch���0�ϵ� ���������!�3�9� ��\�n߀ߒߤ߶��� �������"�4�F�X� j�|�h�K߰������� ��
��.�@�R�d�v� ������������� *<N`r�� �����& ��J\n���� ����/"/4/F/ X/j/|/;�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�/�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_�?L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o=_�o�o�o �o�o�o 2DV hz�����h������u�o.�@��R���Cz  B}��   ���}2&� � _��
���  	�_�2�Տ����_�Kp������ď i�{�������ß՟� ����/�A�S�e�w� ��������N����� �+�=�O�a�s����� ����Ϳ߿���'ψ9�K�_������<�v�_��$SCR_�GRP 1
!�� !�� t� ��� ���	 ������������ ����_������)�a�����&�DE� DW8���l�&�G��CR-35i�A 901234�567890���M-20��8���CR35 ��:�
��������������:֦�Ӧ�G���"&������	��]��o����:��G�H���>���� �������&���ݯ�a�j����g������B�t��������r��A����  @�`���@� ( ?	�=��Ht�P
��F@ F�`z �y������  �$H��Gs0^p��B��7 ��/�0//-/f/ Q/�/u/�/�/�/8��� P�� 7%?����"?�W?-2?<���@]? H�1�?t�ȭ7�������?-4AA, �&E@�<�@G�B�a 3OZOlO�-:HA�H�O�O|O P�B(�B�O�O_���EL_DEFA�ULT  ��_��`S?HOTSTR#]A�7RMIPOWER�FL  i�/U�YTWFDO$V �/URRVENT �1����NU� L!DUM_�EIP_-8�j!AF_INE#P<�_-4!FT�_->��_;o!��`o ��*o�o!RPC�_MAIN�ojh�8vo�o�cVIS�oiiy��o!TPp�PU�Ydk!�
PMON_PR'OXYl�VeZ��2r��]f��!RDM_SRV�r�Yg�O�!R��dk��Xh>���!
�`�M��\i���!?RLSYNC�-9�8֏3�!RO�S�_-<�4"��!�
CE4pMTCO�M���Vkn�˟!	���CONS̟�Wl캟�!��WAS�RC��Vm�c�!���USBd��Xn R���Noӯ������� !��E��i�0���W�RVICE_KL� ?%�[ (%�SVCPRG1���-:Ƶ2ܿ�˰3��	�˰4,�1�˰5�T�Y�˰6|ρ�˰7@�ϩ�˰�����9����ȴf�!�˱οI� ˱��q�˱ϙ�˱F� ��˱n���˱���˱ ��9�˱��a�˱߉� �7߱��_����� ���)����Q�� ��y��'���O��� �w�������� ����˰��İd�c� �����= (as^���� ��/�/9/$/]/ H/�/l/�/�/�/�/�/ �/�/#??G?2?k?V? }?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O�O�O�O	_�O-_���_DEV ~�Y�MC:5X�d�GTGRP� 2SVJ ��bx� 	� 
 ,
�PJ 5_�_�T�_ �_�_o�_'o9o o]o Do�ohozo�o�o�o�o �o�o5{�_g �������� ��?�&�c�u�\��� ����Ϗ���J\)� ��M�4�q���j����� ˟ݟğ��%��� [�B��f������ٯ �������3��W�i� P���t���ÿ���ο ���A�(�e�L�ί ��RϿ��ϸ������  ��O�6�s�Zߗߩ� ���ߴ������'�~� ��]���h���� ���������5��Y� @�R���v��������� @�	��?&cu \������� �;M4qX� ������/�%/ /I/[/B//f/�/�/ �/�/�/�/�/�/3?? W?�L?�?D?�?�?�? �?�?O�?/OAO(OeO LO�O�O�O�O�O�O�O��O_iV �NLy�6 * 		S=>��+c"_�VU@Tn_Y_B����B�2�J�j�@�´~_g_�_@�%�JOGGING��_�^7T(?VjZ��Rf��Y��A�/e�_%o7e�Tt�] /o�o{m�_�o�m?Qi �o�o;)Kq%��o�}os�� ����9�{`�� )���%���ɏ���ۏ �S�8�w��k�Y��� }���ş���+��O� ٟC�1�g�U���y��� ����'����	�?� -�c�Q���ɯ����w� ��s����;�)�_� ����ſOϹϧ����� ����7�y�^ߝ�'� ��ߵߣ�������� Q�6�u���i�W��{� ������=��M��� A�/�e�S���w����� �������=+ aO������u� ��9']� ��M����� �/5/w\/�%/�/ }/�/�/�/�/�/=/"? 4?�/?�/U?�?y?�? �?�??�?9?�?-OO =O?OQO�OuO�O�?�O O�O_�O)__9_;_ M_�_�O�_�Os_�_�_ o�_%oo5o�_�_�o �_[o�o�o�o�o�o�o !coH�o{� �����; �_ �S�A�w�e������� я���7���+��O� =�s�a������П� ����'��K�9�o� ������_���[�ɯ�� �#��G���n���7� ��������ſ���� a�Fυ��y�gϝϋ� �ϯ�����9��]��� Q�?�u�cߙ߇ߩ��� %���5���)��M�;� q�_���߼��߅��� ����%��I�7�m��� ����]����������� !E��l��5� ������_ D�we��� ��%
//��� =/s/a/�/�/�/��/ !/�/??%?'?9?o? ]?�?�/�?�/�?�?�? O�?!O#O5OkO�?�O �?[O�O�O�O�O_�O _sO�Oj_�OC_�_�_ �_�_�_�_	oK_0oo_ �_co�_so�o�o�o�o �o#oGo�o;)_ Mo����o� ���7�%�[�I�k� ���������ُ� ��3�!�W���~���G� i�C����՟���/� q�V������w����� ���ѯ�I�.�m��� a�O���s�������߿ !��E�Ͽ9�'�]�K� ��oϑ�����Ϸ� ���5�#�Y�G�}߿� ����m���i������ 1��U��|��E�� ��������	���-�o� T������u������� ����G�,k���_ M�q���� ���%[I m���	��� //!/W/E/{/��/ �k/�/�/�/�/	?? ?S?�/z?�/C?�?�? �?�?�?�?O[?�?RO �?+O�OsO�O�O�O�O �O3O_WO�OK_�O[_ �_o_�_�_�__�_/_ �_#ooGo5oWo}oko �o�_�oo�o�o�o C1Sy�o��o i�����	�?� �f�x�/�Q�+���Ϗ �����Y�>�}�� q�_�������˟��� 1��U�ߟI�7�m�[� }����ǯ	��-��� !��E�3�i�W�y�ϯ ��ƿ�������� A�/�eϧ���˿UϿ� Q���������=�� dߣ�-ߗ߅߻ߩ��� �����W�<�{��o� ]���������/� �S���G�5�k�Y��� }��������������� C1gU���� ��{����	? -c���S�� ����/;/}b/ �+/�/�/�/�/�/�/ �/C/i/:?y/?m?[? �??�?�?�?? O?? �?3O�?COiOWO�O{O �O�?�OO�O_�O/_ _?_e_S_�_�O�_�O y_�_�_o�_+oo;o ao�_�o�_Qo�o�o�o �o�o'ioN` 9������ A&�e�Y�G�i�k� }�����׏���=�Ǐ 1��U�C�e�g�y��� �֟���	���-�� Q�?�a���ݟ��퟇� �ϯ��)��M��� t���=���9���ݿ˿ ��%�g�Lϋ��� mϣϑϳ�������?� $�c���W�E�{�iߟ� �߯������;���/� �S�A�w�e������ �������+��O� =�s������c����� ������'K��r ��;������ �#eJ�}k �����+Q"/ a�U/C/y/g/�/�/ �//�/'/�/?�/+? Q???u?c?�?�/�?�/ �?�?�?OO'OMO;O qO�?�O�?aO�O�O�O �O__#_I_�Op_�O 9_�_�_�_�_�_�_o Q_6oHo�_!o�_io�o �o�o�o�o)oMo�o A/QSe�����%{,p�$S�ERV_MAILW  +u!��*q~�OUTPUT��$�@�RV� 2�v  $�� (�q�}��SA�VE7�(�TOP1�0 2W� d? 6 *_�π(_������#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u����������Ͽݷ��Y�P��'�FZN_C�FG �u�$�~����GR�P 2�D� ?,B   A[�*q�D;� B\���  B4~�R�B21��HELL���u��j�k��2�����%RSR �������
�C�.�g� Rߋ�v߈��߬������	���-�?�Q��  �_�%Q���(_���,p��⦼�ޖ�g�2,pd�����HK 1�� ��E�@�R� d��������������� ��*<e`r����OMM ������FTOV_�ENB�_���HO�W_REG_UI��(�IMIOFW�DL� �^�)WAIT���$V�1�^�NTIMn���VA�|_)_UNIT����LCTRY�B�
�MB_H�DDN 2W� 2�:%0 �pQ/ �qL/^/�/�/�/�/�/��/�/�"!ON_ALIAS ?e�	f�he�A?S?e? w?�:/?�?�?�?�?�? OO&O8OJO�?nO�O �O�O�OaO�O�O�O_ "_�OF_X_j_|_'_�_ �_�_�_�_�_oo0o BoTo�_xo�o�o�o�o ko�o�o,�oP bt�1���� ���(�:�L�^�	� ��������ʏu�� � �$�Ϗ5�Z�l�~��� ;���Ɵ؟����� � 2�D�V�h�������� ¯ԯ���
��.�ٯ R�d�v�����E���п ���ϱ�*�<�N�`� r�ϖϨϺ���w��� ��&�8���\�n߀� �ߤ�O���������� ��4�F�X�j�|�'�� �����������0� B���f�x�������Y� ��������>P bt����� �(:L�p ����c�� / /$/�H/Z/l/~/)/ �/�/�/�/�/�/? ?�2?D?V?]3�$SM�ON_DEFPR�O ����1 �*SYSTEM*�0m6RECAL�L ?}9 (� �}tpdi�sc 0=>14�7.87.149�.40:1253�2 2 �>314�8 �1�95172�]?O+M}tpc?onn 0 �?�?��?�?�O�O4G
xy�zrate 11 JO\OnO�O_#_6E�E61�?�A�O�O _�_�_�NJ_\_n_�_ o#o6_H_�_�_�_�o �o�_F`�_[omoo�"5F?o�E2896 �o�o��8C�?Sx\n��#� 6O���������o �NW�i�{���1C U����������_S� e�w����-�?�џ� ���������O�a�s� ���(�;�ͯ߯�� ������K�]�o���� $�7�I�ۿ����Ϣ��5�8copy f�rs:order�fil.dat �virt:\tm?pback\I�[��y�
��/�/��mdb:*.*�����ϰߒߤ�7�3x��:\H���Z�[�s߅��(�;�4��a����V� ��������W�r� ���'�:���^���� ������K�]��߀� #6�����l����� ���aJ\n�#<6�H�844 �� ���J\n�0/#/6oHo02[�� �/�/�/9�9����@I/[!y/
??/�0?� �/R*�/?�?�?8H��V&t?�?O)O }5?�?�?�?O�O�O �/�/X?s?�O_(_;? �O_?�O_�_�_�?LO ^O�?�_o$o7O�_�_ mO�_�o�o�O�OP_�O }o 3_E_�oi_�o����y�$SNP�X_ASG 2�����q�� P 0 �'%R[1]�@1.1��y?��c%�!��E�(�:� {�^�������Տ��ʏ ���A�$�e�H�Z� ��~���џ����؟� +��5�a�D���h�z� ����ů�ԯ���
� K�.�U���d������� ۿ������5��*� k�N�uϡτ��ϨϺ� �����1��U�8�J� ��nߕ��ߤ������� ���%�Q�4�u�X�j� ������������� ;��E�q�T���x��� ��������% [>e�t��� ���!E(: {^������ /�/A/$/e/H/Z/ �/~/�/�/�/�/�/�/ +??5?a?D?�?h?z? �?�?�?�?�?O�?
O KO.OUO�OdO�O�O�O �O�O�O_�O5__*_ k_N_u_�_�_�_�_�_ �_�_o1ooUo8oJo��ono�o�o�d�tPA�RAM �u}�q �	��jUP�d9p�ht���pOFT_KB_CFG  s��u�sOPIN_S_IM  �{v�n��p�pRVQSTP_DSBW~�r"t�HtSR �Zy � &�!pINGS EL�_5SEM����vTOP_ON_?ERR  uCy~8�PTN Zu�k�A4�RN�_PR�D��`�VCNT_GP �2Zuq�!px 	r��ɍ���׏���wVD��RP 1	�i p�y��K� ]�o���������ɟ۟ ����#�5�G�Y��� }�������ůׯ��� ��F�C�U�g�y��� ������ӿ��	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�qߘߕߧ߹��� ������%�7�^�[� m����������� ��$�!�3�E�W�i�{� �������������� /ASew�� �����+ =Ovs���� ���//</9/K/ ]/o/�/�/�/�/�/�/ ?�/?#?5?G?Y?k? }?�?�?�?�?�?�?�?�OO)�PRG_CoOUNT8v�k��GuKBENB��FEM�pC:t}O_UPD �1�{T  
 4Or�O�O�O__!_ 3_\_W_i_{_�_�_�_ �_�_�_�_o4o/oAo So|owo�o�o�o�o�o �o+TOa s������� �,�'�9�K�t�o��� ������ɏۏ���� #�L�G�Y�k������� ��ܟן���$��1� C�l�g�y��������� ӯ����	��D�?�Q� c���������ԿϿ� ���)�;�d�_�q��=L_INFO 1��E�@ �2@����������� �ٽ`y*�d��h'��¿���=`y;MY?SDEBUGU@�@����d�If�SP_�PASSUEB?~x�LOG  �ƕ�C��*ؑ� � ��A��UD�1:\�ԘΥ�_M�PC�ݵE&�8�A���V� �A�SAV !�������X����SVZ�TE�M_TIME 1�"���@ 0 � ���X��X����$T1SV�GUNS�@VE'��E��ASK_OPTIONU@�E�A:�A+�_DI��qO�G�BC2_GRP� 2#�I�����@�  C���<Ko�?CFG %z���� �����` ��	�.>dO� s������� *N9r]�� �����/�8/ #/\/n/��Z+�/Z/�/ �/H/�/?�/'??K? ]�k?=�@0s?�?�?�? �?�?�?O�?OO)O _OMO�OqO�O�O�O�O �O_�O%__I_7_m_ [_}__�_�_�X� �_ �_oo/o�_SoAoco �owo�o�o�o�o�o�o =+MOa� �������� 9�'�]�K���o����� ����ɏ���#��_;� M�k�}��������ß �ן��1���U�C� y�g������������� ��	�?�-�c�Q�s� ���������Ͽ�� ��)�_�Mσ�9��� ��������m���#� I�7�m�ߑ�_ߵߣ� ����������!�W� E�{�i�������� ������A�/�e�S� u�w������������� +=O��sa� ������ 9']Kmo�� �����#//3/ Y/G/}/k/�/�/�/�/ �/�/�/??C?��[? m?�?�?�?-?�?�?�? 	O�?-O?OQOOuOcO �O�O�O�O�O�O�O_ _;_)___M_�_q_�_ �_�_�_�_o�_%oo 5o7oIoomo�oY?�o �o�o�o�o3!C iW����� ����-�/�A�w� e����������я� ��=�+�a�O���s� ������ߟ͟��o� -�K�]�o�ퟓ������ɯ���צ��$T�BCSG_GRP� 2&ץ��  �� 
? ?�  6�H� 2�l�V���z���ƿ��������(�d��E+�?�	� HC���>�㙚G����C� � A�.�e�q�C���>ǳ33��S�/�]϶�Y��=Ȑ� C�\  Bȹ��B=���>����PŖ��B�Y�z��L�H�0�$����J�\�n�����@�Ҿ���� �����=�Z�%�7��L���?3�����	V3.00.��	cr35��	*����
�������� 3��4� o  {�CT�Xv�}��J2�)�������CFG -+ץ'� *���+���I����.<
�< bM�q���� ���(L7p [������ /�6/!/Z/E/W/�/ {/�/�/�/�/.�H��/ ??�/L?7?\?�?m? �?�?�?�?�? OO$O �?HO3OlOWO|O�O� ���Oӯ�O�O�O!__ E_3_i_W_�_{_�_�_ �_�_�_o�_/oo?o AoSo�owo�o�o�o�o �o�o+O=s �E���Y��� ��9�'�]�K�m��� ����u�Ǐɏۏ��� 5�G�Y�k�%���}��� ��ßşן���1�� U�C�y�g�������ӯ ������	�+�-�?� u�c����������Ͽ ���/�A�S����� qϓϕϧ�������� %�7�I�[���mߣ� �߳������߷��3� !�W�E�{�i���� ����������A�/� e�S�u����������� ����+aO �s��e���� �'K9o] �������#/ /G/5/k/}/�/�/[/ �/�/�/�/�/??C? 1?g?U?�?y?�?�?�? �?�?	O�?-OOQO?O aO�OuO�O�O�O�O�O �O___M_�e_w_ �_3_�_�_�_�_�_o o7o%o[omoo�oOo �o�o�o�o�o!3 �o�oiW�{�� �����/��S� A�w�e�������я�� �����=�+�M�s� a���������ߟ�_ 	���_ן]�K���o� ������ۯɯ���#� ��Y�G�}�k����� ſ׿�������� U�C�y�gϝϋ��ϯ� �������	�?�-�c� Q�s�u߇߽߫����� ���)��9�_�M�� ��/����i������ %��I�7�m�[����� �������������� EWi{5��� �����A/ eS�w���� �/�+//O/=/_/ a/s/�/�/�/�/�/�/ ?'?��??Q?c??�? �?�?�?�?�?�?O�? 5OGOYOkO)O�O}O�O8�O�O�N  �@S� V_R�$�TBJOP_GR�P 2,�E��  ?��V	-R4S.;\��@|u0{SPU? >��UT� @�@LR	 ߐC� �Vf  C���ULQLQ�>�33�U�R�����U�Y?�@=�ZwC��P��ͥR}��P  B��W�$o/gC��@g��dDb�^��q�eeao�P&ff�e?=�7LC/ka#B o�o�P��P�efb-C�p��^!g`�d�o�PL�Pt�<�eVC\  ֥Q@�'p�`� G A�oL`�_w�C�BrD�S��^�]�_�S�`<PB��P�anaa`#C�;�`L�w�a�Qoxp�x�p:�O�XB$'tMP@�P�CHS��n���=��P����trd<M�gE�2pb����X� 	��1��)�W���c� ������������ ��7�Q�;�I�w���;d�Vɡ�U	V�3.00RScr35QT*�QT�A��� E�'�E�i�FV�#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F����F��3F����F�{G
�GdG߶G#
�D���E'
EM�KE���E��ɑE�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F���vF�u�<#��
<t���Dٵ=�_��V �R�p�V9� ]�ESTPARtp��HFP*SHR\�AB_LE 1/;[%�SG�� �W�GǅG�G� WQG�	�G�
G�GȖ�Q�G�G�G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{� �ߟ߱���w�S]�CS !ڄ�������� ����&�8�J�\�n� ������������ ]\� `��	��(�:��π��
��.�@�w�N�UM  �E*EQ�P	P ۰ܰ�w�_CFG 0���)r-PIMEBF_TTb��CSo��,VERڳ-B�,R 11;[ �8��R�@� �@&  ���� ���//)/;/M/ _/q/�/�/�/�/�/? �/?J?%?7?M?[?m? >�@�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_Rl_�Y@cY�MI_CHAN8� c cDBGL�V��:cX�	`E�THERAD ?Uf�\`��?�_uo�oQ�	`ROUmTV!	
!�d��o�lSNMASK�Qhcba255.�uߣ'9ߣY�O�OLOFS_DI�b��U;iORQC?TRL 2		�	Ϸ~T���� �#�5�G�Y�k�}��� ����ŏ׏������.��R�V�PE_D�ETAI/h|zPG�L_CONFIG� 8�	����/cell/$C�ID$/grp1�V�̟ޟ����Ӏ �o?�Q�c�u�����(� ��ϯ������;� M�_�q�����$�6�˿ ݿ���%ϴ�I�[� m�ϑϣ�2������� ���!߰���W�i�{��ߟ߱�%}F����� ��/�A�C�i�H��Eߞ���������� ?��.�@�R�d�v�� �������������� *<N`r�� �����&8 J\n��!�� ���/�4/F/X/ j/|/�//�/�/�/�/ �/??�/B?T?f?x? �?�?+?�?�?�?�?O O�?>OPObOtO�O�O��O���User View ���}}1234567890�O�O�O_�#_5_=T�P��]_���I2�I:O�_�_�_�_ �_�_X_j_�B3�_Go Yoko}o�o�o o�op^46o�o1CU�ovp^5�o���@��	�h*�p^6� c�u����������ޏp^7R��)�;�M�_�q�Џ��p^8�˟ݟ����%���F�L� �lCamera�J��������ӯ���E~��!� 3��OM�_�q��������y  e��Yz���	� �-�?�Q���uχϙ� 俽���������>��e�5i��c�u߇ߙ� �߽�d������P�)� ;�M�_�q��*�<��i ���������)��� M�_�q���������� ������<�û��=O as��>���� *'9K] f�Q������� /�%/7/I/�m// �/�/�/�/n<��^/ ?%?7?I?[?m?/�? �?�? ?�?�?�?O!O 3O�/<׹��?O�O�O �O�O�O�?�O_!_lO E_W_i_{_�_�_FOXG9+_�_�_oo(o:o �OKopo�o)_�o�o�o��o�o ��	g�0 �oM_q���No ����o�%�7�I� [�m�&l�n��Ə ؏���� ��D�V� h���������ԟ� ��g�ڻ}�2�D�V�h� z���3���¯ԯ��� 
��.�@�R���3uF� 鯞���¿Կ����� �.�@ϋ�d�vψϚ� �Ͼ�e�w���U�
�� .�@�R�d�ψߚ߬� ����������*��� w���v����� ��w�����c�<�N� `�r�����=�w��-� ����*<��` r��������<��  ��1 CUgy����x���    -/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_��  
��(  ��%( 	  y_�_�_�_�_�_�_o 	o+o-o?ouoco�o�ot�o�Z* �Q &�J\n� �����o���9 �(�:�L�^�p���� �����܏� ��$� 6�}�Z�l�~�ŏ���� Ɵ؟���C�U�2�D� V���z�������¯ԯ ���
��c�@�R�d� v�����᯾�п�)� ��*�<�N�`ϧ��� �ϨϺ�������� &�8��\�n߀��Ϥ� ����������E�"�4� F��j�|������ ������e�B�T� f�x������������� +�,>Pb�� �������� (o�^p�� ����� /G$/ 6/H/�l/~/�/�/�/ �//�/�/?U/2?D?�V?h?z?�?�/�`@ A�2�?�?�?�3�7��P��!frh:�\tpgl\ro�bots\m20�ia\cr35ia.xml�?;OMO _OqO�O�O�O�O�O�O�O ���O_(_:_ L_^_p_�_�_�_�_�_ �_�O�_o$o6oHoZo lo~o�o�o�o�o�o�_ �o 2DVhz ������o�
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟�ݟ��&�8�J� \�n���������ȯߟ ٯ���"�4�F�X�j��|�������Ŀ־�8�.1 �?@88�?�ֻ�ֿ �3�5�G�iϓ�}ϟ� �ϳ��������5���A�k�U�wߡ߿��$�TPGL_OUT?PUT ;�!�!_ ���� ����,�>�P�b�t� ������������ �(�:�L�^�p�������������2345?678901���� �����"��B Tfx��4�� ���
}$L ^p��,>�� � //$/�2/Z/l/ ~/�/�/:/�/�/�/�/ ? ?�/�/V?h?z?�? �?�?H?�?�?�?
OO .O�?<OdOvO�O�O�O DOVO�O�O__*_<_ �OJ_r_�_�_�_�_R_ �_�_oo&o8o�_�_ no�o�o�o�o�o`o�o �o"4F�oT|@����\��}������0�B�T�e�@�������� ( 	 ��Џ���� ��<�*�L�N�`��� ������ޟ̟��� 8�&�\�J���n����������ȯ���"���� ���*�X�j�F����� |�¿Կ��C���ϱ� 3�E�#�i�{�忇ϱ� S����������/ߙ� S�e�߉ߛ�y߿��� ;�������=�O�-� s���ߩ��]����� ���'����]�o�� ����������E��� ��5G%W}���� ��g���1 �Ug	w�{� �=O	//�?/Q/ //u/�/��/�/_/�/ �/�/�/)?;?�/_?q? ?�?�?�?�?�?G?�? O�?OIO[O9OO�O �?�O�OiO�O�O�O!_ 3_�O_i_{__�_�_��_�_�_�R�$TP�OFF_LIM �>�op:���mqbN_SV` � l�jP_M�ON <6��dopop2l�aS�TRTCHK �=6�f� bVT?COMPAT-h�a�fVWVAR �>Mm�h1d R�o �oop`ba�_DEFPROG� %|j%ZE�RO ZUZAU�N	�j_DISP�LAY`|n"rIN�ST_MSK  �t| ^zINU�SER�odtLCK��|}{QUICKM�EJp�"rSCRE��p6��btpscdt�q��b�*�_.�ST�jiR�ACE_CFG �?Mi�d`	��d
?�u�HNL 2@|i����k r͏ߏ���'��9�K�]�w�ITEM� 2A�� �%�$1234567�890����  =�<��П��  !���p��=��c ��^���������� .���R��v�"�H�ί ��Я������*�ֿ ���r�2ϖ�����4� ޿�ϰ���&���J�\� n���@ߤ�d�v��ς� �����4���X��*� ��@�����ߨ�� ������T���x��� ���l��������,� >�P�������FX�� d������:� p"��o�� ���F6HZt ~��N/t/�/��/ / /2/�/V/?(?:? �/F?�/�/�/j?�?? �?�?R?�?v?�?QO�? lO�?�O�OO�O*O|O _`O _�O0_V_h_�O t_�O__�_8_�_
o o�_@o�_�_�_Lodo �_�o�o4o�oXojo3 �oN�or��o�(�s�S�B���z��  h��zq ��C�:y
 P��v�]����UD1�:\�����qR_�GRP 1C��� 	 @Cp ���$��H�6�l�Z��|�����f���˟x���ڕ?�  
� ��<�*�`�N���r� ������ޯ̯��&�`�J�8�Z���	�u������sSCB 2D� ���� �(�:�L�^�pς��|�V_CONFIG E���@��������OUTPUT �F����� ��6�H�Z�l�~ߐߢ� �������������#� 6�H�Z�l�~���� ����������2�D� V�h�z����������� ����
�.@Rd v������� )<N`r� ������// %8/J/\/n/�/�/�/ �/�/�/�/�/?!/4? F?X?j?|?�?�?�?�? �?�?�?OO/?BOTO fOxO�O�O�O�O�O�O �O__+O>_P_b_t_ �_�_�_�_�_�_�_o o'_:oLo^opo�o�o �o�o�o�o�o $ ����!�bt��� ������(�:� -o^�p���������ʏ ܏� ��$�6�G�Z� l�~�������Ɵ؟� ��� �2�D�U�h�z� ������¯ԯ���
� �.�@�Q�d�v����� ����п�����*� <�M�`�rτϖϨϺ� ��������&�8�J� [�n߀ߒߤ߶����� �����"�4�F�W�j� |������������ ��0�B�S�f�x��� ������������ ,>Pa�t��� ����(:|L/x���k }gV�K��� //&/8/J/\/n/�/ �/�/W�/�/�/�/? "?4?F?X?j?|?�?�? �?�/�?�?�?OO0O BOTOfOxO�O�O�O�? �O�O�O__,_>_P_ b_t_�_�_�_�O�_�_ �_oo(o:oLo^opo �o�o�o�o�_�o�o  $6HZl~� ���o���� � 2�D�V�h�z������� �ԏ���
��.�@� R�d�v���������Ϗ �����*�<�N�`� r���������˟ޯ� ��&�8�J�\�n���𒿤���Ż�$TX�_SCREEN �1G�g�}ipnl�/��gen.htmſ�*�<�N�`Ͻ�Panel �setupd�}��dϥϷ��������� �ω�6�H�Z�l�~ߐ� ߴ�+�������� � 2�߻�h�z���� ��9�g�]�
��.�@� R�d����������� ����}���<N` r��;1�� &8�\��������QȾU�ALRM_MSG� ?���  �Ȫ-/?/p/c/�/�/ �/�/�/�/�/??6?�)?Z?%SEV  �-�6"EC�FG I���  ȥ@� � A�1   B�Ȥ
 [?ϣ��? OO%O7OIO[OmOO�O�O�G�1GRP �2J�; 0Ȧ	� �?�O I_B�BL_NOTE �K�:T�G�lϢ�ѡ�0~RDEFPRO =%+ (%N?u_ Ѡc_�_�_�_�_�_�_ o�_o>o)oboMo�o�\INUSER � R]�O�oI_M�ENHIST 1}L�9  (�0� ��)/SO�FTPART/G�ENLINK?c�urrent=m�enupage,?1133,1�oD8Vhz~�� }9361���� �r�$�6�H�Z�l�~� �����Ə؏�����  �2�D�V�h�z�	��� ��ԟ���
���.� @�R�d�v�������� Я�����9Rq�� B�T�f�x��������� ҿ����ϩ�>�P� b�tφϘ�'�9����� ����(߷�L�^�p� �ߔߦ�5������� � �$����Z�l�~�� ���C�������� � 2��/�h�z������� ��������
.@ ��dv����� _�*<N� r�����[� //&/8/J/\/��/ �/�/�/�/�/i/�/? "?4?F?X?C�U��?�? �?�?�?�?�/OO0O BOTOfO�?�O�O�O�O �O�O�O�O_,_>_P_ b_t__�_�_�_�_�_ �_�_o(o:oLo^opo �oo�o�o�o�o�o  �o$6HZl~i? {?������ 2�D�V�h�z����-� ԏ���
����@� R�d�v�����)���П ���������N�`� r�������7�̯ޯ� ��&���J�\�n�����������$UI�_PANEDAT�A 1N����ڱ  	�}�����!�3�E�W� )Y�}�7�� �Ϻ��������i�&� �J�\�C߀�gߤߋ� ����������"�4��\X�7�� �q}� �ϕ���������B� ���%�I�[�m���� ��
�����������! E,i{b�� ����l�ܳ 7�<N`r��� �-���//&/8/ �\/n/U/�/y/�/�/ �/�/�/?�/4?F?-? j?Q?�?�?%�?�? �?OO0O�?TO�xO �O�O�O�O�O�OKO_ �O,__P_b_I_�_m_ �_�_�_�_�_oo�_ :o�?�?po�o�o�o�o �oo�o sO$6H Zl~�o���� ��� �2��V�=� z���s�����ԏGoYo �.�@�R�d�v�ɏ ����П����� �<�N�5�r�Y����� ��̯���ׯ�&�� J�1�n�������ȿ ڿ����c�4ϧ�X� j�|ώϠϲ���+��� �����0�B�)�f�M� �ߜ߃��ߧ������� ��P�b�t��� ��������S���(� :�L�^����i����� ������ ��6 ZlS�w�'�9�}���"4FX)�}��l�� ���/j'//K/ 2/D/�/h/�/�/�/�/ �/�/�/#?5??Y?���C�=��$UI_P�OSTYPE  �C�� �	 e?�?�2QU�ICKMEN  ��;�?�?�0RE�STORE 1O�C�  '�L?��6OCC1O��maO�O�O�O�O �OuO�O__,_>_�O b_t_�_�_�_UO�_�_ �_M_o(o:oLo^oo �o�o�o�o�o�oo  $6H�_Ugy �o������ � 2�D�V�h�������� ԏ����w�)� R�d�v�����=���П ������*�<�N�`� r��������ޯ� ��&�ɯJ�\�n��� ����G�ȿڿ������7SCRE�0?��=u1sc�+@u2K�3K�4�K�5K�6K�7K�8<K��2USER-�2ϦD�ksMì�3��4���5��6��7��8����0NDO_CFG P�;� ��0PDATE ����None��2��_INFO �1QC�@��10% �[���Iߊ�m߮��� �����������>�P�3�t��i���<-�O�FFSET T�=�ﲳ$@����� �1�^�U�g������� ���������$-�ZQcu���?�
�����UFRAM/E  ����*��RTOL_ABRqT	(�!ENB*~GRP 1UI��1Cz  A� �~��~����B����0UJ��9MSK  hM@�;N%8��%��/�2VCCMf��V�ͣ#RG�#EY�9���/����-D�BH�p71�C���3711?�lC0�$MRf2_�*PS�Ҵ�	����~XC56 *ȋ?�6���1$�5ڴ��A@3C�N�. ��8�? ��OOKOx1FOsO�5�51��_O�O�� B����A 2�DWO�O7O_�O8_ #_\_G_�_k_}_�__ �_�_�_�_"o�OFoXo.�%TCC�#`mI1��i������ G�FS��2aZ; ��| 2345678901�o�b��� ��o��!5a�4�BwB�`56 311:�o=L�Br5v1 �1~1�2��}/��o�a ��#�GYk} �p�������ُ �1�C�U�6�H���5� ~���ߏ���	���4>�dSELEC)M!�v1b3�VIRToSYNC�� ����%�SIONTM�OU�������F��#bU��U��(u F�R:\H�\�A\��� �� M�C��LOG��  � UD1��EX�����' B@ ����̡m���̡  OBCL�1��H� �  �=	 1- n6  -�������[�,S�A�`=�S�͗��ˢ��TRAIN⯞b�a1l�
0d�$j�T2cZ; (aE2� ��i��;�)�_�M�g� qσϕϧ���������	��F�STAT dm~2@�zߌ��*j$i߾��_GE��#eZ;�`0��
� 02��HOM�IN� fU��U� ~�����Б�C�g�X���JMP�ERR 2gZ;
  ��*jl�V�7� �������������
���2�@�q�d�v�B�_�ߠRE� hWޠ$L�EX��iZ;�a1-�e��VMPHASOE  5��c&���!OFF/�F�PU2n�j�0��
��E1@��0ϒE1!1?s33�����ak/�kxk䜣!
W�m[�䦲�[�����o3;�  [i{�� ��/�O�?/ M/_/q/��/��// �/'/9/�/=?7?I?s? �/�?�/�/�?�??O m?O%O3OEO�?�?�O �?�O�O�?�O�O�O_ _gO\_�OE_�O�_�O �O/_�_�_�_oQ_Fo u_�_|o�o�_�oo�o �o�o�o;oMo?qof -�oI���� �7�[P��� ������ˏ��!�3� (�:�i�[�ŏg�}�������TD_FIL�TEW�n�� �ֲ:���@���+� =�O�a�s�������� �֯�����0�B��T�f�x���SHIF�TMENU 1o[�<��%��ֿ�� ��ڿ����I� �2� �V�hώ��Ϟϰ��������3�
�	LIVE/SNAP'�vsfliv���E����ION� * Ub�h�menu~߃�����ߣ�6��p���	����LE�.�50�s�P��@� ��AɠB8
z�z��}��x�9�~�P�� ����MEb���<�Z0���MO��q����z�WAITD_INEND�������OK1�OU�T���SD��TI]M����o�G� ��#���C���b�������RELEASE�������TM����=���_ACT[������_DATA r��%L�����xRDISb�E_�$XVR�s����$ZABC_G_RP 1t�Q��,#�0�2���ZIP�u'�&�����[MPCF_OG 1v�Q�0��/� w�ɤ�� 	�Z/  85�/�/H/�/l$?��+�/�/�/?�/��/???r?�?  �D0�?�?�?�?�?�;���x�]h_YLIND֑y�� ��� ,(  *VOgM.�SO�OwO�O�M i?�O�O ^PO1_�OU_<_N_�_ �O�_�_�__�_�_x_ -ooQo8o�_�o�oY�&#2z� � ��oC�e?a?>N|h�oq����qA�$D�SPHERE 2{6M��_�;o�� �!�io|W�i��_�� ,��Ï���Ώ@�� /�v���e�؏��p�����������ZZ�� �N