��   m�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING,��<$1_8k	  �FMS*�t *v M_LIF��u,(8*x��M(DSTB0+_0>*_���*#�z&+CL_TIM>�PCCOMi��FBk M� �MAL_�EC�S��P!Q%XO �$PS� �TI����%�"r $D�TY?R. l*1E�ND14�$1�ACST1#4V22\93\9�4\95\96\6_O3VR\6� GA[7�2 h7�2u7�2�7�2�7�2ޜ8FRMZ\6DE��DX\6CURL� HSZ27Fh1DG u1DG�1DG�1DG�1DC�NA!1?( �sPL� + ���STA23TRQ_�M��/@K"�FSUX�JY�JZ�II�JuI�JI�D �$U1�SS  ����6Q����+PV�ERSI� 4W  �5GQ?IRTUAL3_EQ�' 1 TX W ��(P���_�_�_�Vm���څ �!� ���~����������R?����?��J�B�y4���=�t��7�Q��]�����V���u������?�� ��_�P�eieoAQ�o�l	��\�鉵 ��� 
H 	?ȥ�ma͌o�o �_�l/VSetc�$�w�gAPB�w��un�Q� �Su���g`�� ��`���	 j�����& ~����_j��b%��d�op#�5�G���=L��k�t���?�z���@� ����я�����+��=�O�a�s���� �rU������ޟ:T  2��!�3�E�W�i� {���������<��ۯ ����#�5�G�Y�k��}��������$$ �1�\�aO��ԪJ=�;J$��oTP�P����N7��mD��J��:H�a�@�J`BB��@G(�moA���1����m�B�@kB�����`��C+����Pk��.dP �o�Ϙ�ϸ�+�=ϟ�<��M�x���2���V�A�z��� @P�� �֠՞ժ�� ���{Ђ��K�}gL��_3L�X�������L�c�M�ZQ�MZR<MZS�MZZ�U�3�8�H��L�VM]+N�2��q�td �x��t������6Q��Q� ������8NS$�T�i��i�����/U � ���� x
� �x������W��NQ��Q�sQ��WQ�BM�C�T��C���C���������E����������������Ə����%���^���p��C���C�F�C�4�C���C������� �6g��� �7 4�7� m�t �ZN� �X� �W� �Ts �1��5��&N�� �sW� �/4 �4�� �59�m9�z�����{��M���Q�� �_�r�Na�,a��$a� 2���ړ���� ����vc+�W{��M��M��M���M��M�I�������š���}�� t�� 0q�� 1� 1�L� 1ح�ρu���EA��@���s�����������������z��N�w���M�Ƞ7���9��O�K͋ w�3��n	 �1	 i	 � ������1g����F Av��qU�����#��+��&��8��'��>�H)dUc

eAIH�J��`K��k}+*����1sP���RxtesP�E�QV���`hsP�td���8f���ߔ���� 2 ' ��?S	-��TsewasP!?PO��sP�����9�������l>�����hi�AV�s�sP쩀>������ ����+�{� ⩀��H欥���ssP�b�sP�sP�sP���(�����������sPd��ͭ�M��AQ����4-8��P��Ǡ_� =��WS�sP��эiF.D�'ce�+�/`,�/ �$����??���*���I�ڭD�@�^�0g�0p��D��=�.��Ħ^�ħ���0��0�?������&J��L���.c��/mį@�z�0��06��0G�0P�0Y�?��s��0�?�t�_?�.k�����?-��?-���?-��?-��x?���@���?���?)���?�~�?����?�q`!@�?W�r")@�)@���z�w9@��z����鬾��b?��>����I.��\ž��v�u�l���ſ��]�2����!�{�.��zۮ�z+�;y@�y@�9@��@?���@��B�A�=��@K���@5�@D�@N�=%��>y�"�>�w�ޠ��@Gh�@�@?��E�@ߍ@ԍ@���@�5Bh�b�h�Ϊ�@��"�V���>����,����m��;B����f��/�?���?�׫��M?�:E��i�_�hճ��h�9�h�W��hѻ)Pm��B��B��9Q��ݫ�?�K���Jvh�Ju��MP}MP8?�����i��C͆�?+��uߪ9P!5P
5P5P �5P9P�� ,($�not a program|?���_��_�_�_�_PLAC�E�_%o�_Io0hZERXmoTofo�o�o�o�o�o�o4dFRAM��o,7oP7I�(�$A�q_POSP#IC���xA�� _q����#�`� G���k�}�����ޏ���PLCLų��� D�1�ѐ?�  �>���?C�� q�T�m�x�c������� ���������>�P�