��   /8�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CCHG_�LIM_T  � �
$COM�MENT �$CTRL_STATE  M�IO_TYPX
I�DXXUFRAM�E_NUMxTO�OL�INSID~WMARGINX �$UPP_XY�Z4   �$LOW� /C�FG8` Z�$KNOB_MO�UGZ �SE�L�EF�GRIP_wENBOPE� <K CLOSW K �LEVER�;U�gBTN_OUT�XeXuONE�_HANDXAV�G_F�� ROT�_]TRNS� T�R �b�uSFD�OD�  �$ORG_PTH�_RES�TOUCH�OC�*��$JNT4MR�G�2$+$�F+B"2a3�T"k(�SP�8t#�)�WPR�*�)RECa�$e�$�uTEACH_P�AT#MULTI��'�!�&CUST�O�GEN_TPO_PRO< K T�*��� �E=�� =1D�EV�m5���_�AR 2  
�$SB~2+$�0_�RIGH�.!HD_L_MAS��2�C61��1�2�V �1��5�7�5�<�:�<��7m1F_1 x7JFF�_VALID_M��MAX_RUNx� * � GAIN� |G� �2!� I(j!�F� SNGL��B:"H�qB� P��Xp2�D�!u0_R�3�!��T=1C�CUR_F5TSMG@(XqA?PUSH_FlC�@@GYDU=TSU�3;T�C�: �&�!�YJ1_нB�V�@�Z5�[SI�MPLE�AXOF��F�Q�ERSV Nt� �2bREA�0ܻcSTRa?>�0DEBUG� ��/DATA8� N�6�@ ^c@`ce$P� T�PO� -*�#Q2!�g�bk �b�z1�"S R$NE��REBO�2�I�T�OK�cON_�RSThFSA�RI9Tg�cORCW -"x!rJC-"MEAN z�HDGD_ACT�IVWSAFE_WDI1�]tOeu�Nru@�$`GX�P PSKTbNE�`�y3 0LSGS"xGS_WLP-"EX{�q�r+$��@ =`�V\�2!�Q �k  ,��T ��T ��T��rx��t�SMALGA��@OVR������FO=�r�@k ɉ14Ȋ֋5ȉBE|���fAF*��gESCwAPE��TOP<f_$CLAL_aAT�DDSB#QDCS_TCg �|e�% #Q�)#S�Wk��%��� �e�"�j���g�1��@�#Q�H-3�F�eEg�SUB30GtNOc_M�E�b�DB<!8`�I�b�WAI�dc��P�A�rb�'��NT��b��!pP�ڢCN�DOW�C�Nv�fבjד2��M|10�   pB�F�A��F�bDa2�G�RP8 � hA
2�46D�`IL5eIРR��m1DI��{3A�@W{3�5VEN ITYXUR 0MD�'�ΰ꽠128�f}� �$M��0? ���F����Y��Y;�=SIO�NC�  ��5W�IRTU�s`D�V��� d�Y����o���#���1�����ƭ�BȊ������������@���2�C3��B���C��CBWд_��~��1��V��s�� � �b��f��j�B_�  �d_�H��dNЕ�@�Ϩ�
2 N41_01������} K�
 P���������B��X E';� ����-� ������1�C�U�g� y������������ 	��|�?�Q�c�u��� ������������ );M_q���61�B�G�B�f��
?�33~���  �X/4�� ��A�?QcW����f�������V�ba� =�k��aBbC��2&p/� BN�� �������U�M� u?0  �?��!���d��>� @�?L��<#�
�Ҁ�ԭ��#�* "2 3�h/z/�/�/�/�/�/ �/�/
?H�V/3?E?W? i?{?�?�?�?�?�?G�O
 M��? �? OO>O9OKO]O�O�O �O�O�O�ѓ�KaQ`����$1��_ _:_���2��]_�_��8 �����|Q�B����X�@�$E����=����)��|Q>���> � >H�� ;���S����|Q�������B#6迶f�l?]p����H�.Vk_��	cm�<�B�@����A7�@�\��|Q�N  =3���m@����9�=5�B��|Q@2?�?�⾥��@ڱQ��>0?"ȉ@��Z�m�����-�@ɴ���o��o5l��� Cn}_<�o� M& sz������ �у�M�;o"?F�X�j� |�������ď֏�/� ��0�B�T�f�x���������L2�;���'�	!̕h� 2��2� l�O 	M���"�TP�@�� 0�?�KН����  UB؎��� �]�0�@��J�\�n�����3��@���ȯگ���4�@o�"�4�F�X���5q�@۸������Ŀ��6ݿ@G�����0���7I�@��f�xϊϜ���8��@����������9!�@��>�P�b�t�&�1  /��ت߼�������,� b��(�:�L��Ә��� ��������:���  ��$���p���Z�l� ~�����ܿ	������ ����H�~	2DVh �Ӵ��	������  �V
.@�ӌ�@�v���&�2�� .)��//*#d�) N/`/r/�/*#��9�/ �/�/�/*#<�r9&?8? J?\?*#���9�?�?�? �?*#JI�?O"O4O *#��IjO|O�O�O*# �"Y�O�O�O_*#X �YB_T_f_x_*#��Y �_�_�_�_&�30/fi o,o>oPobc�/�i�o �o�o�obc?>y�o (bct?�y^p� �bc�?���� � bcLO��6�H�Z�l�bc �O���Ə؏bc$_ Z�� �2�D�V��_ƙ z�������V��_2����
��V�4ho��R� d�v������o
���Я �����@v�*�<�N� `����⹖�����̿ ���N���&�8Ϛ� ����nπϒϤϚ��� &�������ߚ�\��� F�X�j�|ߚ�ȟ�ٲ� �����ߚ�4�j��0�B�T�V�5������ ��