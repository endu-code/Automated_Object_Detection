��  zE�A��*SYST�EM*��V8.3�0261 5/�21/2018 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� P �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f d PPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$VERSI3 ��!COUPLED�w $!PP_� OCES0s!_81F3�K2> �! � �$SOFT�T�_IDk2TOTAoL_EQs $�0�0NO�2U SPI�_INDE]�5X�k2SCREEN_�(4_2SIGE0�_?q;�0PK_F�I� 	$TH{KYGPANE�4� � DUMMYE1dDDd!OE4LA�!R�!R�	 � $TIT�!$I��N �Dd�DPd �Dc@�D5�F6�FU7�F8�F9�G0�G��GJA�E�GbA�E�G1B�G1�G �F�G2�B~!SBN_CF>"�
 8F CNV_�J� ; �"�!_CM�NT�$FLA�GS]�CHEC��8 � ELLSE�TUP � 7$HO30IO�0� �%�SMACRO��RREPR�X� D�+�0��R{�T UTOBACKU��0 �)DoEVIC�CTI*0��� �0�#�`B��S$INTERV�ALO#ISP_UsNI�O`_DO>f<7uiFR_F�0AIN�1���1c��C_WAkda�jO�FF_O0N�DEL�hL� ?aA�a1b�?9a�`C?���P�1E��#sAT9B�d��MO� �cOE D [M�c���^qREV�B3ILrw!XI� Qr�R  � O�D�P�q$NO^PM�Wp�t�r/"�w� �u�q�r��0D`S p =E RD_E�pCq�$FSSBn&$�CHKBD_SE�^eAG G�"$SLOT_��2=�� V�d�%��3 �a_EDIm  � � �"���PS�`(4%$EP<�1�1$OP�0�2��a�p_OK�UST1P_C� ��dx��U �PLACI4!��Q�4�( raCOsMM� ,0$D冀���0�`��EOWBn�I�GALLOW�� (K�"(2�0V�ARa��@�2ao�Lv�0OUy� ,K�vay��PS�`�0M_�O]����CC�FS_UT~p0 �"�1�3�#�ؗ`X�"�}R0  4F I'MCM�`O#S�`���upi �_�p�B�}�a���M/ �h�pIMPEE_F�N��N���@O���r�D_�~�n�Dry�F� dCC_��r0  T� '��'�DI�n0"��pu�P�$I�������F�t XF� GRP0��M=q�NFLI�7��0U�IRE��$g"� S�WITCH5�AX�_N�PSs"CF_�LIM� �; �0EED��!���qP�t�`PJ_dVЦMODEh�.Z`��PӺ�ELBOF � ������p� ���3���� FB/���0�>�G� �>� WARNM�`/���qP��n�NST�� COR-0bF�LTRh�TRAT�PT1�� $AC�C1a��N ��r$�ORI�o"V�RT��P_S� CHG*�0I��rT2��1
�I��T�I1��>� x i#�Q\��HDRBJ; TCQ�2L�3L�4L�5L�6L�7L� N��9s!V�'�CO`S <F +�=��O��#92��LLEC�y�"MULTI@�b�"N��1�!��O�0�T�� �STAY�"�R`�=l�)2�`����)�`T  |@� �&$��۱m��P��̱�UTO���E��EXT����ÁB���"2� (䈴![0������<�b+�� "D"���� �Q��<煰kcl�9�A#���1��ÂM���P��" '�3�$ L� E���P<�z�`A�$JOBn�xT���l�TRIG3�% dK�������<���\��+�Y�l�_yM��& t�p3FLܐBNG AgTBA� ���M��
 �!��p� �q��0�aP[`��O�'[����0tna*���"J���_R���CDJ���IdJk�D�%C��`�Z���0��P_��P��@ ( @F RaO.��&�t�IT�c�NOM�
���P�SY0�`T)w@����Z�P�d���RA��0��2b"����
$�T����MD3�TD��`U31���p(5!YHGb�T1�*E�7�c�KAb�WAb�cA�4#YNT���PD'BGD�� *(��PUt@X��W����AX��a��eTAI^cBUF��0!�+ � 7n�P�IW�*5 P�7M��8M�9
0�6F�7S�IMQS@>KEE�3PATn�^�a"� 2`#�"�L64F;IX!, ���!dĶ�D�2Bus=CCI��:FPCH�P:BAD�aHCEhAOGhA]H"W�_�0>�0_h@�f �Ak���F�q\'M`#��"�DE3�- l �p3G��@FSOES]FgHBSU�IBS9WC���. ` ��M�ARG쀳��FAyCLp�SLEWx�Qe�ӿ��MC�/�\pSM_JBM����QYC	g��e��0 �n��CHN-�MP�G$G� Jg�_� <#��1_FP$�!TCuf!õ#�����d�#a��V&��r�a;�fJR���rSEG�FR�PIO� S�TRT��N��cP!V5���!41�r�Ӏ
r>İ�b�B�O�2` +�[��� ,qE`�,q`y�Ԣ}t8��yaSIZ%����t�vT�s� �z�y,qRSINF}Oбc����k��`��`�`Lp�ĸ T`7�CRCf�ԣCC/�9��`a�ua8h�ub�MIN��uaPDs�#�G�D�YC��C�����e�q0��� ��EV�q�F�_
�eF��N3�s�ahƔ�Xa+p,5!�#=1�!VSCA?� �A��s1�"!3 ��`F/k��_�U��g���]��C�� a�s�.bR>�4� �����N����5a�R�HA;NC��$LG��P�6f1$+@NDP�t�AR5@N^��a�q���c��ME�18���}0f��RAө�AZ �𨵰�%O��FCT K��s`"�S�PFADIJ�OJ�ʠ� ʠ���<���Ր��qGI�p�BMP�dp�p�Dba��AES�@�	�K�W_��BAS��� �G�5  zM�I�T�CSX[@�@�!62�	$X����T9�{sC��N��`�~P_HEIG9Hs1;�WID�0�VT ACϰ�1�A�Pl�<���EXP�g���|��CU�0M�MENU��7�T[IT,AE�%)��a2��a��8 P�� a�ED�E  ��PDT��REM�.��AUTH_K�EY  ������ ��b�O	����}1E�RRLH� �9 \�� �q-�OR�DB�_�ID�@l �PUN_�O��Y�$SYSP0��4g�-�I�E��EV�#q'�PXW�O�� �: $S�K7!f2%�Td�TR�L��; �'AC��`��ĠIND9DIJ.D��_��f1�Ԭf���PL�A�RWAj���SD�A��!�+r|��UMMY9d�F�10d�&����J�<��}1PR�; 
3�POS��J�g= �$VS$�q�PL~�>��H�SܠK�?����CJ��@����ENE�@TƷ�A���S_�RE�COR��BH �5 O�@=$LA�>$~�r2�R��`��qU�`�_Du��0R	O�@V�T[�Q�U��������! }У�PA�US���dETURYN��MRU� v CRp�EWM�b��AGNAL:s2$�LA�!?$=PX�@$P�y #A �Ax�C0 #ܠDO�`X�k�W�v��q�GO_AWAYF��MO�ae���]��CSS_CCSCB C �'N��CERI��гJ`u�QA0�}��@�GAG� R�0�`�`�{`��{`OF�q`�5��#MA���X��>�LL~�D� �$�� �sU�D)E%!`���OVR10W�,�O�R|�'�$ESC�_$`�eDSBIO�Q��l ��B�VIB&� �c,����8�f�=pSSW���6f!VL��PL����ARMLO
��`0����d7%SC �bcALspH�MPC�h �Ch �#h �#h 5�UU���C�'�C�' �#�$'�d�#C\4�$�pH��Ou��!Y��!�SB���`k$4��C�P3Wұ46$oVOLT37$$`�*�^1��$`O1f*�$o��0RQY���2b4�0DH_THE����0SЯ4�7ALPH�4�`���7��@ �0�qb7�rR�5�88� ×���P"��Fn�M�B�VHBPFUAFLQ"�D�s�`�THR���i2dB�����G(��PVP�����������1�J2�B�E�C�E�CPSu�Y@��Fb3� ��H�(V�H:U�G�
X 0��FkQw�[�Na�'Bx���C INHBcFILT���$�� W�2�T1�[ ���$���H YАAF�sDO��Y�Rp� f g�Q�+�c5h�Q�iSh�QPL���Wqi�QTMOU�#c�i �Q\��X�gmb��vi�hҍbAi�fI�aHIG��ca	xO��ܰ��W�"vAN-u!��V	#AV�H!Pa8C$P�ד#p�R_:�QA�a��B�N0�X�MCN���f1[1�qVE�p��Z2;&f�I�QO�u�rx�w-GldDN{G|d�B�aF>!�9��aM:�NU�FWA�:�Ml� ��X�Lu��$!����!l�ZO����0%O�l1F�s�13�DI�W�@��Q���_��>!CURVA԰0rCR41ͰZ�C<�r� H�v���<�`U�<�(�f�CH�QR3�S��`�t���Xp�VS_�`H�ד�F��ژ���2�NST�CY_ E L����1�t�1��U��U24�2B�NI O7�x�����DEVI|� F��$5�R�BTxSPIB�P����BYX����T���HNDG��G H tn���L��Q�C���5��Lo0 H���f��FBP�{tFE{�5�t��T��I�DyO���uPMCS�v�>�f>�t�"HOT�SW�`s�&шE;LE��J T���e �2��25�� O� ���HA7�E��344�0�鵘�A�K �� M{DL� 2J~PE��	A��s��tː���s�JÆG!��rD"`�ó�����\�TO���W�	��/��SLA�V�L  \0I�NPڐ���`%ن_�CFd�M� �$��ENU��OG���b�ϑ]զP�0x`ҕ�]�IDMA�Sa��\�WR�#��"�]�VE�$a�SKIB�STs��sk$��2u���J�������	��Q܇��_SVh�EX�CLUMqJ2M!ON�L��D�Y��|�PE� ղI_V�AP�PLYZP��HIDX-@Y�r�_M�2��VRFY�0��r�1�cIOC_f�� �1������O��u�L�S���R$DUM�MY3�!���S� L_TP/Bv�"����AӞ�ّ N 9���RT_u��/ �G&r[��O D��P_BA��`�3x�!$F ��_5���H��]����� �� P $<�KwARGI��� �q�2O[�_SGNZ�Q �~P/�/P�IGNs�l�$��^ sQANNUN�@�T<�U/�ߴ�LAzp]	Z�dZ~�EFwPI�@_ R @�F?�IT�	$TOT�A%��d���!ڙM�NIY�S�+���E�A[�
D7AYS\�ADx�@���	� �EFF/_AXI?�TI��0�zCOJA �ADJ_RTRQ��Up��<P�1D D�r5̀Ll�T�p�? ]P�"p��P�A8tpd��V 0w��G��������SK��SU� ��CTR�L_CA�� W>�TRANS�6PIDLE_PW����!��A�V��V_��l�V �DI�AGS���X� �/$2�_SE�#TAC���t!�!0z*L@��RR��vPA��4�p ; SW�!�! �  ��ol�U��o3OH��PP� ��sIR�r��BRK'#��"A_Ak���x 2 x�9ϐZs2��%l��W�pt*�x%RQD�W�%MSx�t5AX��'�"��LIFEC�AL���10��N �1{"�5Z�3{"dp5�xZU`}�MOTN°9Y$@FLA�cZgOVC@p�5HE	>��SUPPOQ�ݑ�Aq� Lj (C�1_�X6�IEYRJZRJW�RJ�0TH�!UC��6�X�Z_AR�p��Y2��HCOQ��Sf6AqN��w$�ICTE��Y `��CACHE�C9�M�P�LAN��UFFIQ@�Ф0<�1	���6
�LN�MS�W�EZ 8�KEgYIM�p��TM~�SwQq�wQ#���Ґ����VIE� �[; A�BGL��/�}�?� 	�?��D�\p�ذST��!�R� �T� �T� �T<	��PEMAIf�ҁ���_FAUL��]�Rц�1�U|�КR�DTRE�^< $Rc��uS�% IT��BCUFW}�W��N_�N� SUB~d��C|�p�Sb�q�bSAV�e �bu �B��� �gX�^AP�d�u+p�$�_~`8�e�p%yOTT���
�sP��M��OtT�Lw#AX � ��X~`9#��c_G�3
�YN)_1�_�D��1� �2M���T��F��H@ g�`� 0p��Gbn-sC_R�AIK���r�t�RoQ�u7hN�qDSPq��rP��A�IM�c6�\����sB2�U�@�A�sM*`#IP���s�!DҐ6�CTH�@n�)�OT�!�6�HSDI3�AB#SC���@ Vy���� �_D�CONVI�G���@3�~`F�!�pd��psq�SCZ"���sMERk��qFB��k��p�ET���aeRFU&:@DUr`����x�CD,���@p;cHR�A!��bp�Ք�Ք+PSԕC��2�C��p�ғ|Sp�cH *�LX�:cd�Rqa�| �� ��W��U��U��U�P	�U�OQU�7R�8R��9R��0T�^�1k�1�x�1��1��1��1���1��1ƪ2Ԫ2T^�k�2x�2��2��U2��2��2��2ƪ�3Ԫ3^�3k�x�3P���o���3��3���3ƪ4Ԣ%�XTk!0�d <� 7h�p��6�pO��p����NaF{DRZ$eT^`�V�Gr����䂴2R�EM� Fj��BOV�M��A�TRO�V�DT�`-�MX�<�IN��0,�W!INDKЗ
w�׀�p$DG~q36��P�5�!D�6�RIVx���2�BGEAR�KIO�%K�¾DN�p���J�82�PB@�CZ_MCM�@�1��@9U��1�f ,②aO? ���PI�.�!?I�E��Q�!���`m���g� _05Pfqg RI9ej��k!UP2_ h � �cTD�p����! a����A�bBAC�ri T�P�b�`Z�) OG��%�8��p��IFI�!�p�m�>��	�PT�"���MR2��j ��Ɛ+"����\� �������$�B`x%��%_ԡ�ޭ_���� M������DGC{LF�%DGDY%LDa��5�6�ߺ4SCHB��UkM`��? T�FS#p�Tl P���e�qP�p$EX_����1M2��2� 3�5���G ���m ���Ѝ�SW�eOe6D�EBUG���%G�R���pU�#BKUv_�O1'� �@PO�I5�5�MS��OOfswSM��E�b�@�0�0_E n �p| P�TERM��o�! �OR�I+�p�2O ��SM_���b�q���A�r�U�IF�UP�Rs� -�1�2n$|�' o$SEG,*�> ELTO��$wUSE�pNFIA�U"4�e1���#$p$UFR���0ؐO!��0����OT�'�TqAƀU�#NST��PAT��P�"PTHJ����E�P rF�V"ART�``%B`�a�bU!REL:�aS�HFT��V!�!�(_�SH+@M$���� ���@N8r����OV9Rq��rSHI%0���UN� �aAYLO����qIl����!�@��@ERV]��1� ?:�¦'�2��%��5��%�RCq��EAScYM�q�EV!WJi'��}�E���!I�2��U@D��q�%Ba��
5aPo��0�p6OR��MY� `GR��t 2b5n� � ���aN�Uu Ԭ")���TOCO!S�1POP ��`�pC�����e��Oѥ`REP�R3��aO�P�b�"ePR�%WU.X1���e$PWR��IM�IU�2R_	S�$VI1S��#(AUD��O`�av" v��$�H���P_ADDR
��H�G�"�Q�Q�Q�БR~pDp1�w H� SZ�a��e�ex�e��SE��r���HS��MNvx ���%Ŕ��OL���p<P��-��ACROlP_!QND_C��ג�1�T� �ROUPT��B_$�VpQ�A1Q�v� �c_��i���i��hx�`�i���i��v�ACk�IOU��D�gfsu<^d�y $|�P�_D��VB`bPR�M_�b�QTT�P_אHaz (��OBJEr��P��[$��LE�#�s>`{ � ��u��AB_x�T~�S|�@�DBGLV���KRL�YHITC�OU�BGY LO: a�TEM��e�0>�+P'�,PSS|�P��JQUERY_F;LA�b�HW��\!�a|`u@�PU�b�PIO��"�]�ӂ�/dԁ=dԁ�� �IWOLN��}����CXa$SLZ�$INPUT_g�$IP#�P��'���SLvpa~��!�\�`W�C-�B�IO�p�F_ASv���$L ��w �F1G�U�B0m!���0�HY��ڑ���᎐U;OPs� `�������[�ʔ[�і"�[PP �SIP�<�іI�2�?�IP_MEMB��ni`� X��IP�P�b{�_N�`�����R�����bSP���p$FOCUS�BG�a~�UJ�Ƃ� �  � o7JO�G�'�DIS[�JY7�cx�J8�7� �Im!�)�7_LA�B�!�@�A��AP�HIb�Q�]�D�� J7J\���� _�KEYt� ��KՀLMONa���$XR��ɀ��?WATCH_��3L���EL��}Sy~�L��s� f �!V�g� �CTR3򲓥v��LG�D� �R����I�
LG_SIZ���J�q IƖ�I�FDT�IH�_�jV� GȴI�F�%SO���q  �Ɩ���v��ƴ��K�AS����w�k�N�
���E��\����'�*�U�s5��@L�>�4�DAUZ�EA`�pՀ�Dp�f�GH�B}�OGBOO�⟇� C���PI�T���� ��REC���SCRN����Dx_p�aMARGf� �`��:���T�L���	S�s��W�Ԣ�Iԭ��JGMO�MNCHL�c��FN��R�Kx�7PRGv�UF��p0n��FWD��HL��STP��V��+���,�Є�RS��H�@����Cr4��?B��� +�O�U�q��*�a28��d��Gh�0PO���������M8�Ģ��E]X��TUIv�I��(�4�@�t� x�J0J�~�P��J0��9N�a�#ANA��O"Ά0VAIA��dCL�EAR�6DCS_CHI"�/c�O�MO�SI��S��IGN_�vpq�u�r��T�d� DEV-�cLLA �°BUW�`��x0T<$U�EM��Ł���*��A�R��x0��σ�a�@OS1�2��3�a�`� �ࠜh�AN%-���.-�IDX�DP�2MRaO��Գ!�ST���Rq�Y{b! �$E&C+��p�.&A&����a� L ��ȟ%Pݘ��T\Q�U�E�`�Ua��_ � �@(��`������# �MB_PN�@ R`r��R�w�TR�IN��P��BAS�S�a	6IRQ6��ϠMC(�� ���CLDP�� ETRQLI��!D�O9=4FLʡh2�Aq3z1D�q7��LDq5[4q5ORG�)�2� 8P�R��4/c�4=b-4�t� �rp[4*�L4
q5S�@TO0Qt�0*D}2FRCLMC@D �?�?RIAt,1ID`�Dg� d1��RQQp=rpDSTB
`�c �F�HAXD2����G�LEXCESH?R�ёBMhPa�Ё�BD4`�B�q`�`�F_A�J�C[��O�H� K��� \ȶ��bTf$� ��LI��q�SREQUIR�E�#MO�\�a�XD�EBU��,1L� M䵔 �p���P�c�AA,1N��
Q�qa�/�&���-cDC���B�IN�a?�RSM�Gh� N#B��N�i�PST9� � �4��LOC�RI쀀�EX�fANGx��A,1ODAQ䵍��@$��9�ZMF�����f��"��%�u#ЖVSUP�' w�FX�@IGGo�� �rq�"��1� �#B��$���p%#by���rx���vbPDATAK�pE;����Rr��M��*� t�`+MD�qI��)�v� ��t�A�wH�`��tD�IAE��sANSW���th���uD��)p�bԣ(@$`� P�CU_�V6�ʠ�A� ��PLOr�$`�HR���B���B�p������$RRR2�E��ɀ ��V�A/A ?d$CALI�@��	G~�2��!V��w<$R�SW0^D�"��ABC�hD_�J2SE�Q�@�q_�J3M�
G�1SPH�,��@PG�n�3m�(u�3p�@��JkC��4�2'AO)IMk@{BCSKP^:ܔ9�wܔJy�{BQܜ��8���`_AZ.B���?�EL��YAOC�MP�c|A)��RT�j���1�ﰈ��@�1�������Z��S�MG��pԕ� ER�!���INҠACk�p����b�
n _�������D4�/R��DIU��C�DH�@
�#a�qc$V�Fc�$x�$���`@���b���̂�E�H ��$BELP����!A/CCEL���kA>°IRC_R�pG0��T!�$P)S�@B2LDp����W3�ط9� ٶPACTH��.�γ.�3���p�A_��_�e�-Br�`C���_MG�$DD��ٰ��$FW�@�p����γ칲��DE��PPA�BN�ROTSPEEu��O0���DEF>Q��Dp$OUSE_��JPQP�C��JY����-A 6qYN�@A�L�̐��L�MOU�NG̭�|�OL�y�INCU��a�¢ĻB��ӑ�AENCS���q�B������D�IN�I`�����pzC�VE��<���23_U ��b^�LOWL���:�O0��0�Di�B�P�Ҡ� ��PRC����M3OS� gTMOpp�@�-GPERCH  M�OVӤ ����� !3�yD!e�]�6�<�$� ʓA����LIʓ�dWɗ��:p3�.�I�T3RKӥ�AY���� ?Q^���m�b��`p�CQ�� MOM�B?R �0u��D���y�0�̂��DUҐZ�S_�BCKLSH_C ����o�n��TӀ����
c��CLAL�J��A��/PKCH�KO0�Su�RTY�� �q��M�1�q_�
#c�_UMCP�	C����SCL���LMTj�_L�0X����E�� �� � ��m�h���6��PC����H� �P��2�CN@�"XT����CN_��N^C�kCSF����V6�����ϡj���nCAT�SHs�����ָ1����֙���������P�A���_P���_ P0� e���O1u�$x�JG� P{#�OG|���TORQU(� p�a�~����Ry������"_W��^�����4Pt�
5z�
5I;I ;Iz�F�`�!��_8�1��VC��0�D�B�2�1�>	P�?�B�5JR�K�<�2�6i�DBL�_SM�Q&BMD`_sDLt�&BGRV4`
Dt�
Dz��1H_��8�31�8JCOSEKr�EHLN�0hK�5oDt� jI��jI<1�J�LZ1�51Zc@y��1MYqA�H�QBTHWMYTHE{T09�NK23z��/Rn�r@CB4VCBn�CqPASfaYR<40gQt�gQ4VSBt��RN?UGTS���Cq���a��P#���Z�C$DUu ��R䂥э2��Vӑ��Q�r�f$N	E�+pIs@�|� �	$R�#QA'UPeYg7EBHBALPHEE.b�.bS�E�c�E�c�E.b��F�c�j�FR�VrhV�ghd��lV�jV�kV��kV�kV�kV�kV�iHrh�f�r�m!�x��kH�kH�kH�kH��kH�iOclOrhOT��nO�jO�kO�kUO�kO�kO�kO�F�F.bTQ���E��egS�PBALANCEl��RLE�PH_'USP衅F��F��FPFULC�3���3��E��1�l�UT�O_p �%T1T2t���2NW������ǡ��5�`�擳�T��OU���� INSsEG��R�REV���R���DIFH��1ٟ��F�1���OB��;C��2� �b~�4LCHWAR���;�ABW!��$MECH]Q�@k�q��AXk�P��IgU�i�� 
���!����7ROB��CR��ͥ�:� �C��_�s"T � x $WEIGHh�F9�$cc�� Ih��.�IF ќ�LAG�K�8SK��K�BI�L?�OD��U��S	TŰ�P�; ���(�������
�Ы�<L��  2�`�"�/DEBU.�L&�n�=�PMMY9��qNA#δ9�$D&�ƪ�$��� Q   �DO_�A��� <	���~�H�L�BX�P�N�Ӣ+�_7�L�t�OH  ��� %��T����ѼT�����TgICK/�C�T1��%������N��c����R L�S���S��ž��PROMPh�E~� $IR� �X�~ ���!�MAI��0��j���_9�����t�l�R�0CO�D��FU`�+�ID�_" =�����G_�SUFF<0 h3�O����DO�� ِ��R��Ǔن�S���P�!{������	�H)��_FI��9��O�RDX� ����3�6��X�����GqR9�S��ZDTD����v�ŧ4 =*�L_NA4���|K��DEF_I[� K���g��_���i���0��š���IS`i  �萚����e��"��4�0i�Dg����D� O��LOCKEA!uӛϭ�0����{�u�UMz�K� {ԓ�{ԡ�{����}� ��v�Ա��g����� ��^���K�Փ����!w�N�P'���^����,`�W\�[R��7�TEFĨ ��OULOMB�_u�0�VIS�PITY�A�!O>Y�A_FRId��F(�SI���R��H����3���W�!W��0��0_,�EAS%��!�& �"���4p�G;穯 h ��7ƵC?OEFF_Om��H�m�/�G!%�S.��߲CA5����u�G�R` � � �$R� �X]�TME�$R�s�Z�/,)ËER�T;�:䗰��  ]�LL��S��_SV�($�~���0���� �"SETU��MEA��Z�x0�u���>��� � � �� ȰID�"���!�*��&P���*�F�'����)3��#�A��"�5;`*�ЧREC���!7�S�K_��� P~	�1_USER���,��4���D�0��VE�L,2�0���2�5S�I���0�MTN�CF}G}1�  ��z�Oy�NORE���3��2�0SI���� ��\�UX-�ܑ�PDE�A $�KEY_�����$JOG<EנSV�IA�WC�� 1DSW�y���
��CMULT��GI�@@C��2� 4 �#t�+�z�XYZ��쑡���zz� �@_ERR��C� ��S L�-����@��s0BB$BU�F-@X17ࡐMO�R�� H	�CU �A3�z�1Q�
��3���$��FV���2SbG�� � $SI�@� G�0VO B`נO�BJE&�!FADJyU�#EELAY' 4���SD�WOU�мE�1PY���=0QT� i�0�W�DIR�$ba�pےʠDY�NբHeT�@��R�^�X����OPWwORK}1�,��SYSBU@p 1SCOP�aR�!�jU�kb�PR��2�ePA�0��!�cu� 1OP��U�J��a'�D�QIMAG�A	��`i�3IMACrIN,�b~sRGOVRD=a�b�0�aP�`sʠ�P �^uz�LP�B�@|��!PMC_E,�Q��N@�M�rǱ��11Ų7�=qSL&�~0����$OVSL \G*E��*E2y�Ȑ�_=p�w��>p�s�� �s	����y��t�#�}1� @�@;���O&E�RI#A��
N��@X�s�f�7���PL}1�,RTv�m�ATU}SRBTRC_T(qR��B �����$ �pƱ��,�~0� D��`-CSALl`�SA���]1gqXE���%����C��J�
���U1P(4����PX��؆��q��3�w� �P�G�5� $SUB������t�JMPWAITO�,�s��LOyCFt�!D=�CVF	ь�y����R`�0��CC_C�TR�Q�	�IGN�R_PLt�DBTeBm�P��z�BW)�d���0U@���IG�az��Iy�TNLN��"Z�R]aK� N��B�0�PE�s���r��f�wSPD}1� L	��A�`gఠ�S��UN��{���]�R!�BDcLY�2���7�_PH_PK�E��2?RETRIEt��2f�b���FI�BǼ ����8� �2��0DBGLV~�LOGSIZ$C��KTؑUy#u�D�7�_�_T1@�EMB�@C\1A����R��|D�FCHECKK��R�P�0����@�&�(bLEc�" PA�9�T���P�C߰P4N�����ARh�0Ґ��Ӯ�PO�BORMATTnaF�f1�h���2�S��UX�y`	�tQPLB��4��  rEITC�H3�8PL)�AL?_ � $��XPRB�q� C,2D�!���+2�J3D���{ T�pPDCKyp���oC� _ALPH���BEWQo����� ��I�wp �� �b@PAYLOYA��m�_1t�2t���J3AR��؀�x�֏�laTIA4��u5��6,2MOMCP@�����������0Bϐ�AD��������PUBk`R��;���;����z��z4�` I$PI\Ds�oӓ1�yՕ�w�2�w�Z��I
��I��I���p����n���y�e`�9S|)bT�SPEED� G��(�Е��/���Е �`/�e�>��M��ЕSAMP�6V��/���ЕMO�@ 2@�A��QP���C��n� ����������LRf`kb`�ІE9h�EIN0 9��7S.В9
yxPy�GAMM%�S���D$GETH)bP�cD]��2
��IB�q�I�G$H�I(0;A��LRE�XPA8)LW VM8z)��tg���C5�CHKKp4]�0�I_��h` eT��n�q��eT�,���� �$^�� 1�iPI� RCH_D�313\��30LE�1�1\�o(�Y�7 �t�MSWFuL �M��SCRc��7�@�&��%n�f�SV���PB``�'��!�B�sS_SAV�&0ct5B3NO]�C \�C2^�0�mߗ�u� �a��u���u:e;��1���8��D�P����� ����)��b9�� e�GE�3��V�7���}Ml�� � ��YL��QNQS RlbfqXG�P�RR#@dCQp� �S:AW70��B�B[�CgR:AMxP�KCL�H���W�r��(1n�g�M�!o��� �F�P@}t$W P�u�P r��P5�R <�RC�R��%�6�`���� ��qsr X��O�D�qZ�Ug�ڐ>D�[ ��OM#w� J?\?n?�?�?��9�b"���e�]�_��� |��X0��bf��qf@��q`�ڏgzf��EڐN� Ag�"�ܰ���FdPB��PM��QU�� � =8L�QCOU!h 7QTHI�HOQBp7HYSY�ES��q�UE�`�"�O��ˋ  �P�@\�U)N���Cf�O�� P��Vu��!�����OGRAƁcB22�O�tVuITe �q^:pINFO����h�{�qcB�e�OI�r�� (�@SLEQ@S��q��p�vgqS�ލ�� 4L�EN�ABDRZ�PTIO�Nt�����Q���)�G�CF��G�$JX�q^r�� R����U�g�+&�_E9D����� �F��P�K��E'N9U߇وAUT$1܅COPY�����n��00MN���PWRUT8R �Nx�;OU��$G[rf�}e�RGADJ����*�X_:@բ$P�����P��W��P��`} ��)�}�EX�kYCDR|�NS.�9�F@r�LGO�#��NYQ_FREQ�R�W� �#�h�TsL�Ae#����ӄ �CcRE� s�IF�ᶕsNA��%a�_}Ge#STATUI`<e#MAIL������q t�������EwLEM�� �/0><�FEASI?�B ��n�ڢ�vA�]� � I�p��Y!q]�Lt#A�ABM���E�pr<�VΡY�BASR҈Z��S�UZ��0�$q���RMS_TR;�qb ���SY��	�ǡ��$���>C��Q`	� 2� _�TM������̲��@ �A��)ǅ�i$D�OU�s]$Nj���P�R+@3���rGRIyD�qM�BARS �sTY@��OTO�Rp��� Hp_}�!����d�O�P/�� �s �p�`POR�s���}���SRV��),����DI&0T��Ѡ�� #�	�#�4!�5*!�6!�7!�8�e��F�2��Ep$VALUt��%��ֱ��>/��� ;�1ėq�����(_�AN��#�ғ�Rɀ(���T�OTAL��S��P�W�Il��REG#EN�1�cX��ks0(��a���`TR��R��_S� ��1ଃV �����⹂Z�E��p��q��Vr���V_Hƍ�DA�S����S_�Y,1�R4�S� AR��P2� ^�IG�_SE	s����å_�Zp��C_�Ƃ�EN�HANC�a� T ;�������GINT�.��@FPs^İ_OVRsP�`@p�`��Lv��o��7�p}��Z�@�SLG�
AA�~�25�	��Dd��S�BĤDE�1U�����TE�P���� !Y��
��J��$2�IL_M`C�x r#_��`TQ�`���q���'�BV�CF�P_� 0�M�	[V1�
V1�2�U2�3�3�4�4�
�!���� � m�A�2IN~VIB�P���1�2�2��3�3�4�4��A@-�C2���=p� MC_Fp+0�0L	11d����M50Id�%"E� �S`�R/�@KEEP_HNADD!�!`$^�j)C�Q�� �$��"	��#O�a_$�A�!K��#i��#REM�"�$��½%�!��(U}�e�$HPW�D  `#SBWMSK|)G�qU�2:�P	�COLLAB� �!K5�B�� 4��g��pITI1{�9p#>D� ,�@F�LAP��$SYNT �<M�`C6���UP_DLYAA�ErDELA�0ᐢmY�`AD�Q���QSKIP=E� i���XpOfPNTv�A�0P_Xp�rG�p �RU@,G��:I+�:IB1 :IG�9JT�9Ja�9Jn��9J{�9J9<��RA=s� X���4��%1�QB� NFLIC�s�@J�U�H�LwNO_H�0�"?��R�ITg��@_PAz�pG�Q� �K�
^�U��W��LV�d�NGRLT�0_q���O�  " ��OS��T_�JvA V	�APPR�_WEIGH�sJg4CH?pvTOR��vT��LOO��]�+�"tVJ�е�ғA�Q�UL�S�XOB'�'���SJ2P���7�X�T�<a43DP=`Ԡ\"p<a�q\!��RDC�ѮL� �рR��R�`� �RV��jr�b�RGE��*��cNFLG�a�Z���SsPC�s�UM_<`>^2TH2NH��P~.a 1� m`�EF11��� �lQ �!#� <�p3AT� g�S�&�Vr�p�t�Mq�Lr���HO�MEwr�t2'r�-?Qcu��w3'r������
�w4'r�'�9�K�]�(o����w5'r뤏���ȏڏ����w6'r�!�3�E�W�i�{��w7'r힟��ԟ���
�w8'r��-�?�Q�Hc�u��uS$0�q�p!�� sF��`la�!,`P�����`/�L��-�IO[M�I֠z��*�POWE��� ��0Za�*��� �5��$�DSB GNAL����0Cpm�S23�23�� �~`���� / ICEQP��P1Ep��5PIT�����OPBx0��FLOW�@TRvP��!U�֤�CU�M��UX�T�A��w�ERFAiC�� U��)a�RSCH��� t�Q  _��>�Q$L����OM��A�`�T�P#UPD7 Ad�ct�T��UEX@8�ȟ�U EFA: X"΁1RSPT����)�T ��PPA�0o�l���`EXP�IOS���)ԭ�_���%Ќ�C�WR�A��ѩD�ag֕`ԦFRIE3NDsaC2UF7P��ޤ�TOOL��MY�H C2LENGT_H_VTE��I�<�Ӆ$SE����?UFINV_����RGI�{QITI5B��Xv��-�G2-�G17�w�S�G�X��_��UQQD�=#���AS��d~C��`��q�� �$$�C/�S�`������S0Ȱ����VERsSI� ��Ȱ�5��I��������AAVM_Y�2� � �0  �5���C�O�@�r� r�	 ����S0�!����������������
?QY�B�S���1��� <-�� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O�OiCC�@XLM�T��C�  ��DIN�O�A�Dq�EXE�HPV_���ATQz
��L�ARMRECOV� �RgLM_DG *�5���OLM_IF 	*��`d�O�_�_�_ �_j�_'o9oKo]onm, 
��odb���o�o�o�o^��$� yz, A   2�D{�PPINFO7 u[ �Vw��������`� ������*��&��`�J���n�����DQ� ���
��.�@�R��d�v���������a
P�PLICAT��?��P��`�Handlin�gTool 
� �
V8.30P�/40Cpɔ_LI
883��ɕ$ME
F0G��4�-

39�8�ɘ�%�z�
?7DC3�ɜ^
�NoneɘVr����ɞ@6�d� Vq_ACT#IVU��C죴�MODP���C�I��?HGAPON����OUP�1*�� i�m�����Қ_����1*� 	 �@����f���� ��Q���Կ�@�
������ ���5�Hʵl�K�HTTHKY_� �/�M�SϹ������� ��%�7ߑ�[�m�� �ߣߵ���������� !�3��W�i�{��� ������������/� ��S�e�w��������� ������+�O as������ �'�K]o �������� /#/}/G/Y/k/�/�/ �/�/�/�/�/�/?? y?C?U?g?�?�?�?�? �?�?�?�?	OOuO?O QOcO�O�O�O�O�O�O �O�O__q_;_M___ }_�_�_�_�_�_�_k�ƭ�TOp��
�DO?_CLEAN9�ꤾpcNM  !{ 衮o�o�o�o�o��DSPDRYRwo&��HI��m@�or ����������&�8�J���MAX@ݐWdak�H�h�XWd��d���PLUG�GW�Xgd��PRC*)pB�`�kaS��Oǂ2DtSEGF0�K� �+��o�o�r����������%�LAPOb�x�� �2� D�V�h�z�������¯�ԯ�+�TOTAL�����+�USENU
O�\� e�A�k­��RGDISPMM�C.���C6�z�@I@Dr\�OMpo�:��X�_STRING� 1	(�
�kM!�S�
���_ITEM1Ƕ  n������+� =�O�a�sυϗϩϻπ��������'�9��I/O SIG�NAL��Tr�yout Mod�eȵInpy�S�imulated�̱Out���OVERRLp =� 100˲In� cycl�̱�Prog Abo�r��̱u�Sta�tusʳ	Hea�rtbeatƷMH Faul	��Aler�L�:� L�^�p��������� ScûSaտ ��-�?�Q�c�u����� ����������)�;M_q��WOR .�û������ +=Oas� ������//'.PO����M � 6/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l?�~?�?�?�?�?H"DEVP.�0d/�?O*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_>n_PALT	��Q �o_�_�_�_�_oo )o;oMo_oqo�o�o�o��o�o�o�o�_GRIm�û9q�_as �������� �'�9�K�]�o�������'�R	�݁Q�� ��)�;�M�_�q��� ������˟ݟ����%�7�I�ˏPREG �^����[�����ͯ߯ ���'�9�K�]�o� ��������ɿۿ�Oݿ�$ARG_� D ?	���0���  �	$O�	[�D�]D��O�e�#�S�BN_CONFIOG 
0˃����}�CII_SA_VE  O������#�TCELLSETUP 0��%  OME_I�OO�O�%MOV�_H������REP���J��UTOBA�CK�����FRA:\o�c Q�o���'`�йo���� �� f�o�����*�p!�3�`�Ԉ��f� ����������o�{� �&�8�J�\�n���� ��������������" 4FXj|�������끁 � ��_i�_\AT�BCKCTL.T�MP 6.VD _GIF PHDp_q��N�t#\��f�INI�P�����c�MESSA�G�����8��OD�E_D����z��Ox�0�c�PAUSM!�!�0� (q73�U/g+(Od/ �/x/�/�/�/�/�/�/ ???P?>?t?1�0$~: TSK  @-x��T�f�UPDT��d�0
&XWZD_ENB����6�STA�0��5"�X�IS��UNT 2�0Ž� � 	� ��z���eng��-뷛�#S�o�U@��H��A��zF�Oo�}Cw쀕g�^����.��O�O�O�O/_2FME�T߀2CMPTAA���@�$A�-�@���@���@���]�5��5�(d�5��P5�r��5F*5�33�8]SCRDCFG� 1�6�Ь�Ź�_�_o@o(o:oLo��o�Q�� �_�o�o�o�o�o�o]o �o>Pbt��0�o9�i�GR<@MX/�s/NA�/�s	i��v_ED��1�Y� 
 ��%-5EDT-��'�GETDA3TAU�o�9��?�(j�H�o�f�\�ּA��  ���2`�&�!�E���:IB ���~�ŏ׏m����3��&۔��D��ߟ@J�����9�ǟ�4�� �ϯ�(����]�o�����5N������ (�w��)�;�ѿ_��6ϊ�gϮ�(�CϮ� ��ϝ�+��7��V� 3�z�(��z�����i߄���8��&���~� ]���F�ߟ�5����!9~������]�����Y�k�����CR �!ߖ���W�q���#��5���Y��p$�NO_�DEL��rGE_�UNUSE��tI�GALLOW 1���(*SYSTEM*S�	$SERV_�GR�V� : RE�G�$�\� N�UM�
��PM�UB ULAY�NP\PMP�AL�CYC1�0#6 $\ULSU�8:!��Lr�BOXO{RI�CUR_�~�PMCNV��10L�T4DLI�0��	����BN/`/r/�/�/�/�/�/���pLAL_OUT �;����qWD_ABO�R=f�q;0ITR/_RTN�7�o	;0�NONS�0�6 �
HCCFS_UT�IL #<�5CsC_@6A 2#; h ?�?�?O#O�6]CE_OPTI�Oc8qF@ROIA_Ic f5Y@j�2�0F�Q�=�2q&}�A_LIMv�2.� ��PM�]B��KX�Pe
�P�2O�Q��B)�r�qF�PQ5T�1)TR�H�_:JF�_PARAMGP7 1�<g^&S�_�_�_�_�VC� W C�d�`�oT!o`�`�`�`�Cd��Tii:a:e4>eBa�GgC�`� �D� D	�`��w?��2HE O�NFI� E?�aG_�P�1#;  ���o1CU�gy�aKPAUS�1�yC , ��������� 	�C�-�g�Q�w����������я���rO�A��O�H�LLEC�T_�B�IPV6�E�N. QF�3�NDE�>� �G�7�1234567890��sB�TR����N%
 H�/%)� ������W���0�B� ��f�x���㯮���ү +�����s�>�P�b� ���������ο�� K��(�:ϓ�^�|��B�!F� �I|�I�O #��<U%�e6�'�9�K���TR�P2$��(9X�t�Y޼`%�̓ڥH��o_MOR�3&�=}��@XB��a ��A�$��H�6�l�~���~S��'�=�r_AA?�a�a`��@K��R�dP��)F�ha�-�_�'�9�%�
�k��G� ��%�Z�%��`�@c..�PDB��+����cpmidbg���	�`:��@ �����p��N W ��@-+
��,�]ܭ@js<��^��@[sgX�$� ysf�l�q��ud1�:��:J��DEFg *ۈ��)��c�buf.tx�t����_L64FIX ,�� ����l/[Y/�/}/�/ �/�/�/
?�/.?@?? d?v?U?�?�?�?�?�?��?,/>#_E -���<2ODOVOhOzO��O6&IM��.o�YU>���d�
�I�MC��2/����dXU�C��20�M�QT|:Uw�Cz  B��i�A���A����Au�gB3��*CG�B<��=w�i�B.��B����B��5B��$�D�%B���ezVC�q��C�v�D����D-lE\D�n�j��B9"6��22o�D|���U'���C�C-����
�xObi�D4cdv`D��`/��`v`s]E�D D��` E4�F�*� Ec��F�C��u[F���E���fE��fF�ކ3FY�F��P3�Z��@�3�3 ;��>L̩��Aw�n,a@��@e�5Y���a���`�A��w�=�`<#����
��?�ozJRS�MOFST (X�,bIT1��D @3��
д����a���;��bw?����<�M�NT�EST�1O�CR�@�4��>VC5`A�w�Ia+a�aORI`mCTPB�U�C�`�4���r��:d�T���qI?�5��q�T_�PROG 	��
�%$/ˏ�t��NUSER  �U�������KEY_?TBL  �����#a��	
��� !"#$%&'�()*+,-./���:;<=>?@�ABC�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~��������������������������������������������������������������������������������͓���������������������������������耇���������������������9�����LCK�
�<���STAT/��s�_AUTO_DO� �	�c�IND�T_ENBP���R�pqn�`�T2����ScTOr`���XC��� 26���8
�SONY XC-�56�"b����@���F( А=�HR50w����>�P�7b�t�Af!f����ֿ� Ŀ� ���C�U�0�yϋ�f� ���Ϝ��������-���TRL��LET�Eͦ ��T_S�CREEN >��kcs����U�MMENU {17�� <� ����w�������� �K�"�4��X�j�� �����������5�� �k�B�T�z������� ��������.g >P�t���� ��Q(:� ^p����/� �;//$/J/�/Z/l/ �/�/�/�/�/�/�/7? ? ?m?D?V?�?z?�? �?�?�?�?!O�?
OWO .O@OfO�OvO�O�O(y~��REG 8�y�����`�M�ߎ�_?MANUAL�k��DBCO��RIG�Y�9�DBG_ER�RL��9�ۉq���_�_�_ ^QNOUMLI�pϡ�p�d
�
^QPXWO_RK 1:���_�5oGoYoko}oӍDBwTB_N� ;������AD�B_AWAYfS^�qGCP 
�=�p�f_AL�pR��bbR�Y�[�
�WX_�P +1<{y�n�,�%o`c�P��h_M���ISO��k@L��sOoNTIMX��
����vy
��2sM?OTNEND�1t�RECORD 1�B�� ���sG�O�]�K��{�b�� ������V�Ǐ�]�� ��6�H�Z������� ��#�؟������2� ��V�şz�������� ԯC���g��.�@�R� ��v�寚�	���п� ��c�χ�#ϫ�`�r� �ϖ�Ϻ�)ϳ�M�� �&�8ߧ�\�G�Uߒ� ߶�����I������4�� �p7�n���� ����������"� ��F�1���|������ ��[�����i���B�Tf���bTOL�ERENC�dB��'r�`L��^PCS�S_CCSCB �3C>y�`IP�t }�~�<�_` r�K�����/�{��5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O��O�O�O�O_�~�L5L� D��&qET|�c�a C[�C��PZP^r_ A�� p� �sp�x�QGPt[	 A�p�Q�_�[? �_�[oU�p�P�pSB�V�c�(a�PWoPio{h+�o�X�o�oY��[	r�h�LW��N:p����}�6ګ�c��aD@VB���|�G���+��K� �otGhXGr�So�����eB   =���Ͷa>�tYB��� �pC�p�q�aA"�H�S�Q-��q����ud�v�����AfP w` 0���D^P���p@�a
�QAXTHQ�z�a a"W>� �a9P��b�e :�L�^�h�Hc�́PQ�RFQ�PU�z�֟ �o\^��-�?��c��u����zCz��ů�b2�Щ�RD�;����l)*��� �S̡0��]�0�.��@���EQ�p��F�X� ѿUҁп�VSȺ�NSTCY 1E��]�ڿ��K� ]�oρϓϥϷ����� �����#�5�G�Y�k��}ߏߒ��DEVI�CE 1F5� MZ�۶a��	� ��?�6�c���	{䰟�����_HNDGD �G5�VP���R�LS 2H�ݠ��/��A�S�e�w����� ZPARAM I��FgHe�RBT [2K��8р<�߬WPpC�C��,`¢�P�Z�����%
{�C��2�jMTLU0,`"nPB, s ���M� }�gT�g��F
B��!�bc y�[2Dchz� ���/��/gT�#I%D��C�`� b!�R��A���A,��Bd��kA��P��_C4kP��!2�C��$Ɓ�]��ffA�À��+B�� �| ���/�/�T (��54a5 �}%/7/d?/M?_? q?�?�?�?�?�?O�? OO%O7OIO�OmOO �O�O�O�O�O�O�OJ_ !_3_�_�_3�_�_�_ �_�_o�_(ooLo^o Ё=?k_IoS_�o�o�o �o�o�o�o#5 G�k}���� ���H��1�~�U� g�y�ƏAo�Տ��� 2�D�/�h�S���go�� ��ԟ����ϟ��� R�)�;���_�q����� �����ݯ�<��%� 7�I�[�m�������� �}�&��J�5�n�Y� �ϤϏ��ϣ�ѿ�� ����F��/�Aߎ�e� w��ߛ߭��������� B��+�x�O�a��� ���������,���%� b�M���q��������� ������L#5 �Yk}���  ��61CU g������� �	//h/���/w/�/ �/�/�/�/
?�/.?@? I/[/1/_?q?�?�? �?�?�?�?�?OO%O rOIO[O�OO�O�O�O �O�O&_�O_\_3_E_ W_�_?�_�_�_�_�_ "ooFo1ojoE?s_�_ �om_�o�o�o�o�o0 f=Oa�� �������� b�9�K���o���Ώ�� [o��(��L�7�I����m������$DC�SS_SLAVE L���ё���_4�D  љ��C�FG Mѕ��������F�RA:\ĐL-�%04d.CSV���  }�� ���A� i�CHq�z��@����|�����"�������Ρޯ̩�Ґ-矩*����_CR�C_OUT N�������_FS�I ?њ ����k�}����� ��ſ׿ �����H� C�U�gϐϋϝϯ��� ������ ��-�?�h� c�u߇߽߰߫����� ����@�;�M�_�� ������������� �%�7�`�[�m���� ������������8 3EW�{��� ���/X Sew����� ��/0/+/=/O/x/ s/�/�/�/�/�/�/? ??'?P?K?]?o?�? �?�?�?�?�?�?�?(O #O5OGOpOkO}O�O�O �O�O�O _�O__H_ C_U_g_�_�_�_�_�_ �_�_�_ oo-o?oho couo�o�o�o�o�o�o �o@;M_� �������� �%�7�`�[�m���� ����Ǐ������8� 3�E�W���{�����ȟ ß՟����/�X� S�e�w���������� ����0�+�=�O�x� s���������Ϳ߿� ��'�P�K�]�oϘ� �ϥϷ���������(� #�5�G�p�k�}ߏ߸� ������ �����H� C�U�g������� ������ ��-�?�h� c�u������������� ��@;M_� ������� %7`[m� ������/8/ 3/E/W/�/{/�/�/�/ �/�/�/???/?X? S?e?w?�?�?�?�?�? �?�?O0O+O=OOOxO�sO�O�O�O�O�C�$�DCS_C_FS�O ?�����A P �O�O_?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo ~o�o�o�o�o�o�o�o 72DVz� ������
�� .�W�R�d�v������� ������/�*�<� N�w�r���������̟ ޟ���&�O�J�\� n���������߯گ� ��'�"�4�F�o�j�|� ������Ŀֿ�������G�B�T��OC_RPI�N_jϳ��� �ς��O����1�Z�U��NSL��@&�h߱� ��������"��/�A� j�e�w������� ������B�=�O�a� ���������������� '9b]o� ������� :5GY�}�� ����///1/ Z/U/g/y/�/�/�/�/ �/�/�/	?2?-???Q? z?u?��ߤ߆?�?�? �?OO@O;OMO_O�O �O�O�O�O�O�O�O_ _%_7_`_[_m__�_ �_�_�_�_�_�_o8o 3oEoWo�o{o�o�o�o �o�o�o/X Sew����� ���0�+�=�O�x� s���������͏ߏ� ��'�P�K�]�o������ �PRE_CH�K P۪�A ~��,8�2x��� 	 8�9�K���+�q���a� ������ݯ�ͯ�%� �I�[�9����o��� ǿ��׿���)�3�E� �i�{�YϟϱϏ��� ��������-�S�1� c߉�g�y߿��߯��� �!�+�=���a�s�Q� ����������� ���K�]�;�����q� ������������#5 �Ak{�� ����CU 3y�i���� ��/-/G/c/u/ S/�/�/�/�/�/�/? ?�/;?M?+?q?�?a? �?�?�?�?�?�?�?%O ?/Q/[OmOO�O�O�O �O�O�O�O_�O3_E_ #_U_{_Y_�_�_�_�_ �_�_�_o/ooSoeo GO�o�o=o�o�o�o�o �o=-s� c������� '��K�]�woi���5� ��ɏ��������5� G�%�k�}�[������� ן�ǟ����C�U� o�A�����{���ӯ�� ��	��-�?��c�u� S�������Ͽ῿�� ���'�M�+�=σϕ� w�����m������%� 7��[�m�K�}ߣ߁� ���߷����!���E� W�5�{��ϱ���e� ������	�/��?�e� C�U������������� ��=O-s� ���]���� '9]oM�� �����/�5/ G/%/k/}/[/�/�/� �/�/�/�/?1??U? g?E?�?�?{?�?�?�? �?	O�?O?OOOOuO SOeO�O�O�/�O�O�O _)__M___=_�_�_ s_�_�_�_�_o�_�_ 7oIo'omoo]o�o�o �O�o�o�o!�o1 W5g�k}�� ����/�A��e� w�U�������я��o ����	�O�a�?��� ��u���͟����� '�9��]�o�M����� ����ۯ��ǯ�#�ů G�Y�7�}���m���ſ �����ٿ�1��A� g�E�wϝ�{ύ����� ��	�߽�?�Q�/�u� ��e߽߫ߛ������� �)���_�q�O�� ������������ 7�I���Y��]����� ����������!3 WiG��}�� ��%�A�1 w�g����� �/+/	/O/a/?/�/ �/u/�/�/�/�/? �/9?K?�/o?�?_?�? �?�?�?�?�?O#OO GOYO7OiO�OmO�O�O �O�O�O_�O1_C_%? g_y__�_�_�_�_�_ �_�_o�_+oQo/oAo �o�owo�o�o�o�o �o);U__q� �������%� �I�[�9����o��� Ǐ�����ۏ!�3�M ?�i��Y�������՟ �ş����A�S�1� w���g�����������ӯ�+�=��$DC�S_SGN Q�K�c��7m� �16-MAY�-19 09:2�0   O�l�4-�JANt�8:38�}����� N.DѤ����������h�x,rWf*�σ�^M��  �O�VERSION� [�V3�.5.13�EF�LOGIC 1R�K��  	���P�?�P��N�!�PROG_E_NB  ��6����o�ULSE  �TŇ�!�_AC�CLIM�����Ö��WRSTgJNT��c��K�EMOx̘��� ���INIT S.��G�Z���OPT_S�L ?	,��
 	R575��VY�74^�6_�7_�+50��1��2_�@�����<�TO  �Hݷ���V�DE�X��dc����P�ATH A[�A�\�g�y��HC�P_CLNTID� ?��6� �@ȸ����IAG_�GRP 2XK�� , `���� �9�$�]�H������1234?567890����S�� |�������8!�� ��H؀��;�dC�S��� 6�����. �Rv�f�� H��//�</N/ �"/p/�/t/�/�/V/ h/�/?&??J?\?�/ l?B?�?�?�?�?�?v? O�?4OFO$OjO|OO E��Oy��O�O_�O 2_��_T_y_d_�_,
�B^ 4�_�_~_ `Oo�O&oLo^oI��T jo�o.o�o�o�o�o  �O'�_K6H�l �������#� �G�2�k�V���B]� ��Ǐُ�������(���L�B\Drx�@���PC�����4  79֐�$��>���:������ߟʟܟ���CT_�CONFIG �Y��Ӛ��egU���STBF/_TTS��
��b�����Û�u�O�MA�U��|��MSW_�CF6�Z��6��O�CVIEW��[ɭ������-�?� Q�c�u�G�	�����¿ Կ������.�@�R� d�v�ϚϬϾ����� ��ߕ�*�<�N�`�r� ��ߨߺ�������� ��&�8�J�\�n��� !�������������4�F�X�j�|����R%C£\�e��!*�B^ ������C2g�{�SBL_FAULT ]��ި�GPMSKk��*��TDIAG ^�:�աI��U�D1: 6789?012345�G�BSP�-?Qc u��������//)/;/M/� ��
@q��/$�TORECP��

� �/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOi/{/xO��/UMP_OPT�IONk���ATR�¢l��	�EPME�j��OY_TEMP�  È�3B��J�P�AP�DU�NI��m�Q��YN_BRK _ɩ��EMGDI_S�TA"U�aQK�XPN�C_S1`ɫ �PFO�_�_�^
�^dpO oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�E� ����y�Q���  �2�D�V�h�z����� ��ԏ���
��.� @�R�d��z������� ˟����%�7�I� [�m��������ǯٯ ����!�3�E�W�i� ��������ÿݟ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�{�iߗߩ� ��տ������'�9� K�]�o������� �������#�5�G�Y� s߅ߏ�����i����� ��1CUgy �������	 -?Qk�}��� ������//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?u?�?�?�?��? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_m?w_�_ �_�_�?�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 Ke_W����_�_ ����#�5�G�Y� k�}�������ŏ׏� ����1�C�]oy� �������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;���g�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�_�i� {ߍߟ߹��������� ��/�A�S�e�w�� ������������ +�=�W�E�s������� ��������'9 K]o����� ���#5O�a� k}�E����� �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-?GYc?u?�?�? ��?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_Q? [_m__�_�?�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /I_Sew� �_������� +�=�O�a�s������� ��͏ߏ���'�A 3�]�o�������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����9�K�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��������ߑ� C�M�_�q߃ߝ��߹� ��������%�7�I� [�m��������� �����!�;�E�W�i� {��ߟ����������� /ASew� ������ 3�!Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?+=G?Y? k?!?��?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ #?5??_Q_c_u_�?�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o-_7I [m�_����� ���!�3�E�W�i� {�������ÏՏ��� �%/�A�S�e�q� ������џ����� +�=�O�a�s������� ��ͯ߯����9� K�]�w���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�1�C�U�g߁� �ߝ߯���������	� �-�?�Q�c�u��� ���������m��)� ;�M�_�y߃������� ������%7I [m����� ���!3EWq� {������� ////A/S/e/w/�/ �/�/�/�/�/�/�/ +?=?O?i_?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O? �$EN�ETMODE 1�aj5� W 005�4_F[PRROR_PROG %#Z�%6�_�YdUTAB_LE  #[t?��_�_�_gdRSEV�_NUM 2R  �-Q)`dQ�_AUTO_EN�B  PU+SaT_;NO>a b#[EQ}(b  *��`���`��`��`4`+��`�o�o�oZdHIS�%c1+PSk_ALMw 1c#[ �4�l0+�o;M _q���o_b``  #[aFR�z�PTCP_VER� !#Z!�_�$�EXTLOG_R�EQ�f�Qi,�SsIZ5�'�STKR��oe�)�TOL�  1Dz�b��A '�_BWD�p��Hf��D�_DIn�� dj5Sd�DT1KRņSTEP�я�P��OP_D�Ot�QFACTO�RY_TUN�gd�<�DR_GRP s1e#YNad 	����FP��x�̹ ��� ��$�f?�� ���ǖ ��ٟ�ԟ���1�� U�@�y�d�v�����ӯ�����LW
 J�#Z&�,��tۯ��j�U���y�B�  �B୰���$  �A@��s�@UUU�Ӿ�������E��� E�`F@ Fǂ5U/�,��L����M��Jk��Lzp�JP���Fg�f�?�  s��9�Y�9}�9���8j
�6���6�;��A����O ���� � I ߵ�����[FE�ATURE f�j5��JQH�andlingT�ool � "�
PEngl�ish Dict�ionary�d�ef.4D �St�ard� � 
! hA�nalog I/�OI�  !
I�X�gle Shi�ftI�d�X�ut�o Softwa�re Updat?e  rt sѓ��matic Ba�ckup�3\s�t��ground Edit���fd
C_amera`�Fd��e��CnrRnd�Im���3�Co�mmon cal�ib UI�� E�the�n��"�M�onitor�L�OAD8�tr�R�eliaby�O�E�NS�Data A�cquis>��m�.fdp�iagn�os��]�i�Doc�ument Vi�eweJ��870�p�ual Ch�eck Safe�ty*� cy� �h�anced UsF��Fr����C ��xt. DIO 6:�fi�� m8���wend��ErrI��L��S������s _ t Pa�r[��� ���J944�FCTN M�enu��ve�M� �J9l�TP In�T�fac{�  7�44��G��p Mask Exc��g�� R85�T���Proxy S�v��  15 J��igh-Spe���Ski
� R7�38Г��mmuwnic��ons�oS R7��urr�T�d�022��aю��connect �2� J5��In{cr��stru,����2 RKA�REL Cmd.� L��ua��R8�60hRun-T�i��EnvL�oaz��KU�el +��s��S/Wѹ�7�License��޷�rodu� og�Book(Sys�tem)�AD �pMACRO�s,��/Offsl��2�NDs�MH��� ����MMRxC�?��ORDE� echStop��t? � 84fM�i$�|� 13dx���]е�׏���Mo}dz�witchIءVP��?��. �sv��2Optmp�8�2��fil���I ��2g 4 �!+ulti-T�����;�PC�M funY�P�o|���4$�b&Re�gi� r �Pr�i��FK+7���g Num SelW�  F�#�� A�dju���60.8��%|� fe���&Otatu�!$6����%��  9 J6�RDM Ro�bot)�scov�e2� 561��R�emU�n@� 8� (S�F3Serv�o�ҩ�)?SNPX b�I��\dcs�0}�Li�br1��H� İ5� f�0��58���So� tr�ss�ag4%G 91"�p ��&0���p{/I��  (ig ?TMILIB(MӞ��Firm����gqd7���s�Acc��2��0�XATX�H'eln��*LR"1Ҽ�Spac�Ar�quz�imula�H��� Q���TouF�Pa��I��T���c��&��ev. �f.svUS�B po��"�iP��a��  r"1Unexcept���`0i$/����H59� VC&�r��[�6���P{��RcJPR�IN�V�; d T�@�TSP CSUiI�� r�[XC�~�#Web Pl6��%d -c�1R��@4d�����I�R6�6?0FV�L�!FVGr�idK1play �C�lh@����5Ri�R�R.@���R-3�5iA���As�cii���"��� s51f�cUpl� N� (T����S���@rityAvo�idM �`��CE��rk�Col,%�@�GuF� 5P���j}P����
 B�L�t^� 120C C� Ao�І!J��P��y�ᤐ� o=q�b @D�CS b ./��c@��O��q��`�; �t��qckpaboE4��DH@�OTШ�m�ain N��1.�H��an.��A> aB!FRLM���!i� ���MI De�v�  (�1� h8j��spiJP��� �@��Ae1/�r���y!hP� M-2� �i��߂^0i�p6��PC��  iA�/'�Passwox�qT�ROS 4�d���qeda�SN��Cli����G6x9 Ar�� 47�!��:�5s�DER��T�sup>Rt�I�7� (M�a�T2DV��
�3D TriA-���&��_8;�:
�A�@Def?�����Ba: deRe p 4t0��e��+�V�st64M�B DRAM�hs86΢FRO֫�0�Arc� vis�I�ԙ�n��7| )�, �b�Heal�wJ�\h��Cel�l`��p� �sh�[��� Kqw�c� #- �v���p	VC�v�tyy�s�"Ѐ6�ut��v��m���xs ���TD`_0��J�m�` 2��ya[�>R tsi��MAILYk�/F�2�h��ࠛ 90 �H��F02]�q�P5'���T1C��5����FC��U�F9�G'igEH�S�t�0/�A� if�!2��b]oF�dri=c �/OLF�S����" H5k�OPT ��49f8����cro6��@���l�ApA�Syn.(RSS) 1L�d\1y�rH�L� (20x5�5�d�pCVx9��.��est�$SР���> \pϐSSF�en$�tex�D o�� �A�	� BP���a�(R00�Qirt��:���2)�D��1�e��VKb@l Bu�i, n��WAPLf��0��Va�kT�X#CGM��D��L����[CRG&a�YB	U��YKfL��pf�ܳk�\sm�ZTAPf�@�О�Bf2��@���V#�s���� r���CB���
f���WE��!��
��B�T�p��DT�&�4 Y�V�`��EH0����
�61Z��
b�R=2�
�E (Np��F�V�PK�B���#"��Gf1`?G���QH�р?I�e ��F��LD�L��N��7\s@���`���=M��dela<,��u2�M�� "L[P��`?��_�%�Ԍ���S��-F�TStO�W�J57���VGF�|�VP2֥ 5\b�`0&�c V:���T;T� �<�ce,?VPD^��$
T;F�־DI)�<I�a\�so<��a-�6Jc6s 6�4L�M�V9R�h���Tri�� ���5�` �f�@�������P
�� ����`��Img� PH�[l��IM/A  VP�S��U�Ow��!%S�Skastdpn)ǲt��� SWIMEST��BFe�00��-Q�� �_�PB�_�Rued�_�T�!�_�S �<�_bH573o2c12��-oNbJ5N�Io$jb)�Cdo�cxE��o �_�lp��o�TdP�o�c �B�or�2.rٱ(0Jsp�EfrSEo�f81�}�r3 RGoe'ELS��sL��� �s�����B	��S\ �$�F�ryz�ftl�o~�g�o������� ��?�����P  �n�&�"�l ��T�@<�@^��Y��e�u8Z���alib��Γ��`ɟ3���埿�\v �F�e\c�6�Z�f��T�v�R VW���8S��UJ91����i�Lů[c91+o�w8���847�:��A 4�j��Q��t6�m���vrc.����HR����ot�0ݿ���  ��8ޯ�4�60�>eS0L�9�7���U�ЄϦ�60 .� g�н�+��'�ܠd�Ϻ�8co��DM�B�U"�����ߕpi��f�T! ��na;�� ���u%��ⅰI��loR�d��1a�59gϱŭ���9I5�ϔ�R����1�� ?��o�#��1A�/��2�vt{�UWeǟ��L�ￇ73[���7��΁�C W��62$K�=fR���8���� ����d����2�ڔ@����@�@" "http���೿t7 �� v R7��78����4�8� ��TTPT�#8	��ePCV4/v�2��j�Q�Fa7��$1N�0�/2�rIO�)/8;/M/6.sv3�64�i�oS�l? tor�ah?*�|`�?��AM/�?
??.?0�k/��1 JO��� ,O�tro���[P��OB4�c.K?�g'�)�24g?�� (B�Od�3\iOA5sb�?U_�?vi�/i��/�/W!n��`�o%�Fo�4�l�$of��oXF I9)xo�cmp\7��3mp���duC��lh����o(A�_Bt� �o]6P��m�I?�w�@L���naO��4*O�0wi�%P�?"�bsg?�]7�YEM����8woVJ�/ե11�?o��DMs�BC���7J�\���(�52�XFa AP�ڟ<�qv�`/şaqs�����/Of��1$�9�VRK����ph�քH5+�=�I9N/¤SkiW�/�IF��_�%��#fs�I�O�l�����"<𜿚$�`����\�jԿz5bO�vrou�ς�3(�ΤH ( DϮ��?sG��|��F�O u�������D)O��*�3P$�FӅ�k���P����럴� �PL��<ʿ��pbox�ߦe3bo���Sh �>��R.�0wT{����fx6��P��D��3���#_I\m;YEe��OԆM�hxW�=Etse,���dct\���O$kR������Xm*���ro3��D�l�j9��V'�  FC���|@��ք f?6KARqE0�_�~ (Kh���.cf���Wp1oO�_K�up��a����H/j#- Eq�d/�84���$qu �o��/ o2o?Vo<�7C�)�s�NJԆ�<|?�3l\sy�?�40�?Τwio�u]?f�w58�?,F�$O�J�
?Ԇ"io�!�Vd��u&A��PR���5, s��v1\�  H55�2B�Q21p0�R78P510�.R0  nel J614Ҡ�/WATUqP��d8P545*��H8R6��9V�CAM�q97PCRqImP\1tPUIF�C�8Q28  ing`sQy0��4P P63P� @P PSCH��DOCVڀD �PGCSU���08Q0=P�qpVEIOC�r��� P54Pupd�PR69aP���PwSET�pt\hPQ�`Qt�8P7`Q�!�MASK��(POPRXY���R7B#�POCO  \pppb36���PR�Q���b1Pd60Q$cJ�539.eHsb��v�LCH-`(��OPLGq\b�PQ0]`��P(`HC�R��4`S�aun�d�PMCSIP`e0�aPle5=Ps�p(`DSW� �  qPb0`�aPa��(`PRQ`Tq�R�E`(Poa601P<cP�CM�PHcR0@q\j23b�V�`E`�S`UPvisP`E`p c�`UPcPRS	a��bJ69E`sFRyDmPsRMCN:e�H931PHcSNB�ARa�rHLB�USaM�qc�Pg52�f�HTCIP0cTMI�L�e"P�`eJ �PyA�PdSTPTX6p;967PTEL�p���P�`�`
Q8P8$Q4�8>a"PPX�8P95��P`[�95qqbU�EC-`F
PU�FRmPfahQCmP90ZQVCO�`@PwVIP%�537sQ7SUIzVSX�P�S�WEBIP�SHTTnIPthrQ62aPd�!tPG���cIG؁��`c�PGS�eIsRC%��cH76�P"�e Q�Q|�Ror��R51P s:P�P,t�53=P8u8=Py�C�Q6]`�b�PI��qs52]`sJ56E`0s���PDsCL�qPt�5�\rd�q75LUP cR8���u5P sR55]`,s� P 8s��P�`CP�PP�SwJ77P0\o��6��cRPP�cR6¼ap�`�QtaT�79�P`�64�Pd87]`�d90P0c��=P�,���5�9ta�T91P� ��1P(S���Q�pai�P06=P-+ C�PF�T	����!aLP PTS�pL�CKAB%�I БIQ`� ;�H�UPPaintPMS�Pa��D�IP�|�STY%�t\patPTO�b�P�PNLSR76�`�5�Q���WaNN�Paic�qNNE`�ORS��`�cR681Pin�t'�FCB�P(�6Hx�-W`M�r��!(`{OBQ`plug�`�L�aot �`OP�I-���PSPZ�PkPG�Q7�`73Β�PRQad�R]L��(Sp�PS���n�@�E`�� v�PTS-�� W��P�`apw�`��P�`cFVR�PlcV39D%�l�PBVI�SwAPL�Pcyc+P�APV1�pa_�C{CGIP - U���L�Prog+PCCQR�`�ԁB�P �PԁK=�"L�P��p��(h�<�P��h�̱��@g�Bـ
TX��%���CTC�pt�p��2��P927"�0ҝPs2�Qb��TC�-�rmt;�	`#1�ΒTC9`HcCTEֵPerj�EIPp.�p/�E�P�c��I�ukse��Fـvrv�F%���TG�P� CP\��%�d -h�H-�wTra�PCTI�p���TL� TRS����p�@נ��IP�PT�h�M%�lexsQT=MQ`ver, �p¸SC:���F��Pv\qe�PF�IPSV"+�H�$cj�ـtr�aC�TW-���CPVGF�-��SVP2mPv\fx���pc�b��e���bVP4�fx_m8��-��SVPD-��SwVPF�P_mo�`iV� cV��t\��=LmPove4��-�.sVPR�\|�tP]V�Qe5.W`V6� *u"��P}�o`���`��'CVK��N�IIP��sCV����IPN9�Gene���D��D��R�D����  ��f�谔�pos.��inal��n��De�R���`��d�P��o9mB���on,���Rh�D�R��\��TXf��D$b��omp�� #"N��P��m���s! ��=C-f����=FXU������g F��(��Dt CII��r�D��u��� "����Cx_u�i X������f20��h	Crl2��D�,r9ui�Ԣ� �it2c�0cov��e"����ا�(.)� ����� ��� I�QnQ �I[� ��_= wo���,bD� �w�|GG� ������4� �e� v�{�� ��&� �2��Z uz������� �ֻTW&q~q 5{�׷&�o? �;0��  �2�� �y� �{��W&��� �?�3� A�ޗe�/> �\��3&T��� 7�7߸ ����� ���� ֵ���&��8 �wl1��S�) ￸�d *J�� F's ~w��� 6:0� ���,��s�-� Q�v� ��{� �,�T ��ZBLx6���v6 ��6���'Par ��s>�E���j�6dsq��F�  �������ЁDh�el�����ti-S�� �Ob��D�bcf�O�����t OFT��P<A�_ �V�ZI��D��V\��qWS��= dtl�e�Ean�(bzd���titv�Z�zҀEz XWO Hq6�6���5 H�6/H691�E4܀To�fkstF� Y68�2�4�`�f804&�E91�g�`30oBkmon_�E��eݱ��� qlm��0 �J�fh��B�_  �ZDTfL0�f(;P7�EcklKV� �6|��D85��ّ�m\b����xo�k�7ktq��g2.g����yLbkLVts6��IF�bk���<���Id I/f��GR� �han��L��Vy��%��%er�e�����io�� �ac�- A�n��h���cuACl�_�^ir��)�g��	�.�@�& G��R630���p v�p�&0H�f��un��cR57v�OJavG��`Y��owc��-ASF��O��7�����SM�����
;af��rafLEa�vl�\F c�w� a���?VXpoV �3�0��NT "L�FFM��=����yh	a��G-�w�� �m2�.�,�t��̹�6�ԯ��sd_�MC'V����D���f�slm�isc.�  H5�522��21&dc.pR78�����0�708�J614Vip? ATUu�@��OL�545ҴIN�TL�6�t8 (�VCA���ss?eCRI��ȑ��UI���rt\r�L�28g��NRE6��.f,�63!��n,�SCH�d EkЏDOCV���p��C�,�<�L�0Q�isp���EIO��xE,�5�4����9��2\;sl,�SET����lр�lt2�J7��ՌMASK���̀PRXY�҇��7���OCO��J6l�3�l�� (SVl�A�H�LѸ@Օ��539Rs�v���#1��LCyH���OPLGf�outl�0��D��wHCR
svg��1S@�h��CSa�!�F{�50��D�l�5!�\lQ��DSW��S����̀��OP����7&��PR���L�ұ��(Sgd���PC�M���R0 \s"��5P՝���0���,n�q� AJ�1��N�:q�2��PRSa����69�� (Au�FRD�Խ��RgMCN���93A��ɐCSNBA:�F9� HLB��� AM��4���h�2A�;95z�HTCaԈ��TMIL6�j95�,��857.,P�A1�ito��TP�TXҴ JK�TEIL��piL�� XpL�80�I)��.�!���P;�J95��s �"N���H�UECޑ�7\cs�FR��<Q��C��57\�{VCOa�,���I�P1jH��SUI��	CSX1�A�WEBa��HTT\a�8�R62��m`���GP%�IG %t{utKIPGSj�v| RC1_me��H76��7P�w�s_+�?x�R51�\iw�N���H�S53!��wL�8!�h�R66��H����ࠡ��@;J56@��1���N0��9�j��L���R5`%�A|�%5q�r�`,�8 5��F{165!��@�"5��6H84!�29��0���PJ���n B�[�J77!Ԩ�R6 �5h3n���y36P��3R6��-`;о Ԩ�@��exeKJ8�7��#J90!�s�tu+�~@!䬵�vk90�kop�B����@!�p�@|BA��g*�n@!��Q��06�!�@[�F�FaP�6؁�́,�TS� N]C[�CAB$iͰl1I��R7��@q��y�CMS1�ro�g+QM�� �� TY�$x�CTOa�nvA\+��1�(�,�6��con�~0��15.��JNN�%e:��P��9ORS%x����8A�815[�FCBaUnZQ�P!��p{���CMOB��"G���OL��x�OPI.�$\lr[�SŠ�T�	D7�U��CPRQ&R9RL���S�V�p~`���K�ETS�$ 1��0���3�Ԩ��FVR1�LZQV31D$ ���BVa�SwAPL1�CLN[�sPV��	rCCGa�̙��CL�3CC�RA�n "W!B��H�CSKQn\`0�p��)�0CTP�n�ЌQe��p!$b�Ct�aT0U�pC�TC�yЋRC1�1� (�s��trl,��r��
TX��TC�aerrm�r�MCq"�s��#CTE���nrr�REa�XP8j�^��rmc�^�a"�P�QF!$���.$p "�rG1�tKTG$c8��QH�$�SCTI�! s���CTLqdACKЋRp)��rLa�R82��M��YPk�.����OF��.���e�{�C`N���^�1�"M� ^�a�С�Q`US��!$���M�QW�$m�V{GF�$R MH��;P2�� H5� ΐpq��ΐ�$(MH[�VP�uoY����$)���D��hg��VP=F��"MHG̑`et!�+�V/vpcm��N��ՙ�N��$�VP1Rqd)��CV�x�V� "�X�,�1�($T�Ia�t\mh��K��etpK�A%Y�1VP%ɠ�!PN����GeneB�rip�����8��exCtt���Y�m� "�(��HB��� )��x�������<Ȣ�res.�yA�ɠn����*����p�@M�_�NĀ6�L���Ș�y�AvL�Xr�Ȉ2��"9R;�Ƚ\ra��	Pދ� h86��Gu0+ʸ�Ͽ�SeLɨm�9�69�P�Ȩr��0�2�ɹ1��n2�h�a �0L�XR}�RI{�!e� L�x���c������N�vx�L��"��2\r�]�N�82�d���b�ɉa��y1���/�k�@���A��r�uk�ʘ L�sop��H�}�ts{������s��9��j96�5��Sc��h��5' J9�{�
�PL��J	een��t �I[
x�com��Fh�L�4 J�޻fo��DIF+�6x�Q����rati|�d�p��1�0�
R8l߂��M�����P��8� �j�mK�X�H�Z����N�odڠ��3�q��vi����80�~�l S0l�yQ��tpk�xb�j�.�@�R�d��@����,/n(�8�8�0���
:�O8�<�Q�}�CO���PT��O (��.�Xp|�~Hx���?�v �3wv��8�22�pm����722��j7`�^�@ƙ���cf��=Yvr���vcu ���O�O�O�O_#_�5_7�3Y_��wv4�{_�_w�ʈ�usst_�_�cus�_ �Z��oo,o>oPo�io��nge��(pLyw747�jWel��HM47ZKEq p{���[m�MFH�?�(wsK�8J�np���o��fhl;N��wmf���? :t�}(4	<g J{�N�II)̏މw�ڎX�774kﭏ/7n�tˏ݊e+���se�/�aw��8�ɐ��)EX \�!+: �p���~�00��nh�,:M�o+�xO��1 "K,�O��\a��#0�� .8���{h�L?�j+�'mon�:��t�/�st�?-�w�:��ڀ)�;��(=h�;
d� Pۻ�{:  ���� �J0��r�e����ST�D�!treL�ANG���81�\tqd�������rch.�����^�htwv�WWּ�� R79��"{Lo�51 (��I�W�h�Ո�4�aw)w� �vy �w623c�h a?�cti�֘!�X�Iiؠ�t ��n,� �։����j�Տ"AJP@�3p�v�r{�H�6��!��-7 SeT� E3�) �G�J934��LoW�4 (S�����8� <���91 ��8!4�j9�所+���y��
��	�btN�ite{�R ��I@Ո� ����P�������	 8����Z�vol��X ���9�<�I�p���ldt*���F�864{��?��K�	�k扐x�֘1�wmsk��AM�q�Xa�e�����p��0R�BT�1ks.OPTN�qf�U$ =RTCamT�� y��U��y��U��UlU6L�T�1Tx����SFq�Ue��6T��USP W��b DT�qT2 h�T�!/&+��TX�U\j6&�U 8U�UsfdO&��&ȁT���662_DPN�bi��%�Q�%62V��$����%�� �#(�(6To6e St�%��#�5y�$�)5(ToB�%tT0�%5�W6T��8�%�#�#orc��#�I���#���%cct��6ؑ?�4\W69�65"p6}"�#\j�536���4�"�?k#ruO O,Im?N�p�C �?t�0<O�;�e �%���?
;g=cJ7 "AV�?�;avsf�O__&_F8WtpD_V_0GT�FD|_:UcK6�_�_r�ON�3e\s�O2^y`O�:�migxGvgW! m�%��!�%T�$E A{6�po6��#337N�)5R5_2E���$0���$Ada�Vd���V�?;Tz7�_�e7DDTF9����#8�`�%��4y�ted Z@�A}�@�}�04N�}�}����}�dc& }����u 6�v��v1�u1\b�u$2}���}� R83�u�"}��"}�valg����Nrh�&�8�J�Y�ox�ue��� j70�v�=1��MIG�uer�fa��{q���E�N��ء��EYE�ce A���񁏯pV� e�A!���2Յ�Q�%��u1�e�i�@��H�e����J0� '��b���T��E In�B��  W�|��537�g����(MI�t��Ԇr��ݟ�am����nеv!g�U -�v J߆8⹖F���P�y�ac���2���R�ɏ jo��2�� �djd�8r}� o#g\k�0��g��wwmf�Fro/�� Eq'�4"}�3 sJ8��oni[���ᅩ}Ĵ�� o�� ��ʛ��m@�R�eD��{n�Д�V�o��x����  �����裆"POS�\����ͯ men�ϖ�⑥OMo�43���� �(Coc� �An[�t���"e�a�\�vp��.��cflx$�le��8�hr��tr�NT� C]F+�x E/�t	qi�M�ӓxc��p�f�clx����Z�cx���
0 h��h8��mo��=� H���)�{ (�vSER,�p��g�0߆0\r�v�X�= ��I � - ��ti��H��VC.�828�5��L"v�RC��n G/�d��w�P�y�\v�vm "o�lϚ�x`���=e�ߠ-�R-3�?������vM [�AX�/2�)�S�rxl2�v#�0��h8߷=�/ RAX�A���t��9�H�E/Rצt����h߶"RXk���F�˦85��2sL/�xB885_�:q�Ro�0iA��5\rO�9�K��v��Ĳ��8���.�n Y"�v��88��8s� i ?�9 ��/�8$�y O�MS"���<&�9R H74&�`�745�	p��p���ycr0C�c�hP0� j�-�a%?o��6D950R7trlܣ�ctlO�AP1C���j�ui"�L���  ����^���!�A��qH��&�-^7����; ��616C�q��794h���� M��ƔI��99���(��$FEA�T_ADD ?	����Q%P  	�H._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ��������TDEMO f~Y    WM_����� ���//%/R/I/ [/�//�/�/�/�/�/ �/�/?!?N?E?W?�? {?�?�?�?�?�?�?�? OOJOAOSO�OwO�O �O�O�O�O�O�O__ F_=_O_|_s_�_�_�_ �_�_�_�_ooBo9o Koxooo�o�o�o�o�o �o�o>5Gt k}������ ��:�1�C�p�g�y� ������܏ӏ���	� 6�-�?�l�c�u����� ��؟ϟ����2�)� ;�h�_�q�������ԯ ˯ݯ���.�%�7�d� [�m�������пǿٿ ���*�!�3�`�W�i� �ύϟ����������� &��/�\�S�eߒ߉� ���߿�������"�� +�X�O�a������ ����������'�T� K�]������������� ����#PGY �}������ LCU�y ������/	/ /H/?/Q/~/u/�/�/ �/�/�/�/???D? ;?M?z?q?�?�?�?�? �?�?
OOO@O7OIO vOmOO�O�O�O�O�O _�O_<_3_E_r_i_ {_�_�_�_�_�_o�_ o8o/oAonoeowo�o �o�o�o�o�o�o4 +=jas��� �����0�'�9� f�]�o���������ɏ �����,�#�5�b�Y� k���������ş�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c������� ������� ��)� V�M�_όσϕϯϹ� ��������%�R�I� [߈�ߑ߫ߵ����� ����!�N�E�W�� {����������� ��J�A�S���w��� ���������� F=O|s��� ���B9 Kxo����� �/�/>/5/G/t/ k/}/�/�/�/�/�/? �/?:?1?C?p?g?y? �?�?�?�?�? O�?	O 6O-O?OlOcOuO�O�O �O�O�O�O�O_2_)_ ;_h___q_�_�_�_�_ �_�_�_o.o%o7odo [omo�o�o�o�o�o�o �o�o*!3`Wi �������� &��/�\�S�e���� ����������"�� +�X�O�a�{������� ���ߟ���'�T� K�]�w���������� ۯ���#�P�G�Y� s�}��������׿� ���L�C�U�o�y� �ϝϯ��������	� �H�?�Q�k�uߢߙ� �����������D� ;�M�g�q������ ����
���@�7�I� c�m������������� ��<3E_i ������� 8/A[e�� ������/4/ +/=/W/a/�/�/�/�/ �/�/�/�/?0?'?9? S?]?�?�?�?�?�?�? �?�?�?,O#O5OOOYO �O}O�O�O�O�O�O�O �O(__1_K_U_�_y_ �_�_�_�_�_�_�_$o o-oGoQo~ouo�o�o �o�o�o�o�o ) CMzq���� �����%�?�I� v�m���������ُ����;�  2�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas��������'9  :>Ug y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{��������/=C 6Yk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ������/�A��$�FEAT_DEM�OIN  E���q��>�Y�INWDEXf�u��Y��ILECOMP �g������t�T���SET�UP2 h������  N �ܑ��_AP2BC�K 1i�� G �)B���%�C�>���1�n�E�� ��)���M�˯����� ��<�N�ݯr������ 7�̿[��ϑ�&ϵ� J�ٿWπ�Ϥ�3��� ��i��ύ�"�4���X� ��|ߎ�߲�A���e� ����0��T�f��� ������O���s�� ���>���b���o��� '���K��������� :L��p����5 �Y�}�$�H �l~�1�� g�� /2/�V/� z/	/�/�/?/�/c/�/ 
?�/.?�/R?d?�/�? ?�?�?M?�?q?O�?�O<O���P� }2�*.VRCO�O�0*�O�O�3�O�O�5w@PC�O_�0�FR6:�O=^�Oa_�KT���_�_&U��_�\h�R_�_�6*#.FzOo�1	(So�El�_io�[STM� �b�o�^+P�o�m��0iPenda�nt Panel�o�[H�o �g�o8Yor�ZGIF|���e�Oa��ZJPG �*��e���z�F�JJS�����0@����X�%
Java?Scriptُ��CSʏ1��f�ۏ �%Cascad�ing Styl�e Sheets�]��0
ARGNA�ME.DT���<�`\��^���Д៍�}АDISP*ן ���`$�d��V�e���CLLB.ZIX��=�/`:\��\������Colla�bo鯕�	PANgEL1[�C�%�` ,�l��o�o�2a�ǿ@V���r����$�3忀K�V�9���ϝ�$�4 i���V���zό�!ߘ��TPEINS.X3ML(�@�:\<�����Custom Toolbar}���PASSWOR�D���>FRS:�\��� %Pa�ssword Config��?J� ��C��"O��3����� i����"�4���X��� |�����A���e��� ��0��Tf��� ��O�s� �>�b�[�' �K���/�:/ L/�p/��/#/5/�/ Y/�/}/�/$?�/H?�/ l?~??�?1?�?�?g? �?�? O�?�?VO�?zO 	OsO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_;_M_�_q_o�_�_ <o�_`o�_�o�o%o�o Io�o�oo�o8�o �on�o�!��W �{�"��F��j� |����/�ďS�e��� ������T��x�� ����=�ҟa������ ,���P�ߟ񟆯��� 9����o����(�:� ɯ^�����#���G� ܿk�}�ϡ�6�ſ/� l�����ϴ���U��� y�� ߯�D���h��� 	ߞ�-���Q߻��߇���,��$FILE�_DGBCK 1�i������ ( ��)
SUMMAR�Y.DG,���M�D:`����D�iag Summ�ary���
CONSLOG��y�����$���Console log%����	TPACCN���%g�����T�P Accoun�tinF���FR�6:IPKDMPO.ZIP����
���)����Excep�tion-����MEMCHECK������8�Mem�ory Data|��LN�)�RIPE���0�%� Pa?cket LE����$Sn�STA�T*#� �%LStatuys�i	FTP��/�/�:�mment TBD=/�� >)ETHERNE�/o��/�/��Ethe�rnU<�figu�raL��'!DCSVRF1//)/B?��0 verif�y allE?�M�(5DIFF�:? ?2?�?F\8di�ff�?}7o0CH�GD1�?�?�?LOc �?sO~3&�
I�2BO)O;O�O 8bO�O�OGD3�O�O�OT_ �O{_
V�UPDATES�.�P�_��FRS�:\�_�]��Up�dates Li�st�_��PSRB?WLD.CMo����Ro�_9�PS_ROBOWEL^/�/:GIG��o>_��o�GigE ~��nosticW~�N�>�)�aHADOW�o�o�o�b�Shado�w Change���8+"rNOTI?=O���Notificx�"��O�A�PMIO�o��h�p�f/��o�^U�*��UI3�E�W��{�U	I������B���f� �_�������O���� �����>�P�ߟt�� ����9�ί]�򯁯� (���L�ۯp������ 5�ʿܿk� Ϗ�$�6� ſZ��~��wϴ�C� ��g���ߝ�2���V� h��ό�߰���Q��� u�
���@���d��� ���)��M������ ���<�N���r���� %�����[����& ��J��n��3 ��i��"� X�|��A� e�/�0/�T/f/ ��//�/=/�/�/�$�$FILE_�P{PR�P��� ����(�MDONLY 1�i5�  
 �z/Q?�/u?�/�?�? t/�?^?�?O�?)O�? MO_O�?�OO�O�OHO �OlO_�O_7_�O[_ �O_�_ _�_D_�_�_ z_o�_3oEo�_io�_ �oo�o�oRo�ovo �oA�oew� *��`�����&�O��*VISBC�K,81;3*.V�DV����FR:�\o�ION\DA�TA\��/���Vision V?D filȅ� �&�<�J�4�n���� ��3�ȟW������"� ��F�՟�|������ m�֯e������0��� T��x������=�ҿ a�s�ϗ�,�>���b� ��ϗϼ�K���o� �ߥ�:���^���������*MR2_GR�P 1j;��C4  B�}�	� 71������E��� E�  F?@ F�5U�������L���M���Jk�Lz�p�JP��Fg{�f�?�  S������9�Y9}��9��8j�
�6��6�{;��A�  �ﶵ�BH��B���B����$��������������@UUU #�����Y�D�}�h��� ������������
�C��_CFG =k;T M����]�NO ^:
F0� � �\�RM_CHKT_YP  0�}�h000��OM�_MIN	x����50X� SSuBdl5:0��bx�Y���%�TP_DEF_O�W0x�9�IR�COM��$G�ENOVRD_D�O*62�THR�* d%d�_E�NB� �RA�VC��mK�� ���՚�/3�/���/�/�� �M!O�UW s��}�x�ؾ��8�g��;?�/7?Y?[?  C��0����(7�?�<B�?B����2�ٸ*9�N SMTT#t�[)��X�4�$HO�STCd1ux����?�� MC�x��;zOx��  27.0�@1�O  e�O�O	_ _-_;Z�O^_p_�_�_��LN_HS	anonymous�_�_�_�oo1o yO��Fh Fk�O�_�o�O�o�o�o �oJ_'9K]�o �_�����4o �XojoG�~�o^��� ����ŏ����� 1�T���y������� ����,�>�@�-�t� Q�c�u���������ϯ ���(�^��M�_� q�����ܟ� �ݿ� �H�%�7�I�[Ϣ�� �ϣϵ����l�2�� !�3�E�Wߞ���¿Կ ����
�������/� v�S�e�w������ �������+�r߄� ��s�����߻����� �����'9K]�� �������4� F�X�j�l>��}� �����// 1/T��y/�/�/�/��/.D\AENT 1=v
; P!J/?  ��/3?"? W??{?>?�?b?�?�? �?�?�?O�?AOOeO (O�OLO^O�O�O�O�O _�O+_�O _a_$_�_ H_�_l_�_�_�_o�_ 'o�_Koooo2o{oVo �o�o�o�o�o�o5 �oY.�R�v���zQUICCA0���3��t14��"����t2��`�r��ӏ!ROUTE�Rԏ��#�!P�CJOG$���!�192.168�.0.10��sC�AMPRTt�P�!�d�1m�����RT�폟�����$NAM�E !�*!R�OBO���S_C�FG 1u�) ��Aut�o-starte�dFTP& ��=?/֯s���� 0�B��f�x������� ��S������,�� �������ϼ�ޯ���� �����ʿ'�9�K�]� oߒ�ߥ߷�������8��SM%y� {�U�ό������� ����
��.�@�c����v������������z �%�7�I�K�8�\ n���k���� �3�FXj|�����a��7 /M*/</N/`/ r/9�/�/�/�/��/ �/?&?8?J?\?�m? ���?�//�?�?O "O4O�/XOjO|O�O�O �?EO�O�O�O__0_ w?�?�?�?�O�_�?�_ �_�_�_o�O,o>oPo boto�_o�o�o�o�o �oK_]_o_L�o�_ �o�����o� � �$�6�Y�Y�~���𢏴�ƏZ�_ERR� w3�я�PDUSIZ  g��^�p���>�W�RD ?r�Cq��  guestb�Q�c�u��������`�SCDMN�GRP 2xr�;���H�g��\�b�K� 	P01.00 8`��   � ��   B  ���� ���_H���L��L�}�L�����O8�`����l�����a4�U  �Ȥ� �8����\���)�`�;��������d�.�@�R�ɛ_GWROUېy������	ӑ���QU�PD  ?u�����İTYg�����TTP_AUT�H 1z�� <�!iPenda�n��-�l���!�KAREL:*8-�6�H�KC]�m���U�VISION SET���ϴ�!�����R�0�� H�Bߏ�f�x��ߜ߮����CTRL {�����g�
��?FFF9E3��At�FRS:DEF�AULT;�F�ANUC Web Server;� )����9�K��ܭ����������߄WR_�CONFIG �|ߛ ;��I�DL_CPU_P5CZ�g�B�I�y�w BH_�MINj��)�}�GNR_IO���g���a�NPT?_SIM_D_������STAL_S�CRN�� ���T�PMODNTOL8������RTY��y����� �ENO���Ѳ�]�OLNK 1}��M���������eMAST�E��ɾeSLAV�E ~��c�O�_CFGٱBU�O�O@CYCL�En>T�_ASG� 1ߗ+�
  ����//+/=/ O/a/s/�/�/�/�/���NUM��
�@IPCH�^R?TRY_CNZ��@�@��������1 @kI�+E��z?E�a�P_MEMBERS 2�ߙ�� $���2����ݰ7�?�9a�SDT�_ISOLC  �����$J23�_DSM+�3J?OBPROCN���JOG��1�+��d8�?��+�O�/?
�LQ�O__/_�OS_e_w_�_`�O Hm@���E#?&BPOSRE�QO��KANJI_����a[�MONG ����b�yN_ goyo�o�o�o�Y�`3	�<� ��e�_ִ���_L���"?`EY�LOGGINL�E�������$L�ANGUAGE Y��<T� {q��LGa2�	�b����g�xP��  *��g�'��b����>�MC:�\RSCH\00�\<�XpN_DISP �+G�H��O��O߃LOCp�D�z���AsOGB?OOK ����`��󑧱����X� ����Ϗ����a�*��	p������!�m��!���=p_B�UFF 1�p��2F幟���՟�D� Collaborativǖ ���F�=�O�a�s��� ����֯ͯ߯����B�9�K���DCS ��z� =��� '�f��?ɿۿ���H@�{�IO 1��# ~?9Ø��9�I� [�mρϑϣϵ����� �����!�3�E�Y�i� {ߍߡ߱��������-E��TMNd�_B� T�f�x�������� ������,�>�P�b��t�������L��SE�VD0��TYPN1�$6���Q�RS"0&��<2FLg 1�"�J0��� �����G�TP:pOF�NGNAM1D�mr�t7UPS�GI"5�a�O5�_LOAD�N@G %�%�TI�pZUZAU�N#�(MAXUALRM�'���(��'_PR"4F0d��1��B_PNP� V� 2�C	M�DR0771ߕz�BL"8063%�@ �_#?�ߒ|/�C��z�6��/􈃟/Po@P 2���+ �ɖ	~T 	t  ��/ �%W?B?{?�k?�? g?�?�?�?O�?*OO NO`OCO�OoO�O�O�O �O�O_�O&_8__\_ G_�_�_u_�_�_�_�_ �_o�_4ooXojoMo �oyo�o�o�o�o�o �o0B%fQ�u �������� >�)�b�M�����{��� �����Տ��:�%��^�p�S�������D�_LDXDISA�pB�MEMO_{APjE ?C
 �,�(�:��L�^�p������� ;1�C ���� 4�������4��X����C_MSTR ����w�SCD 1���L�ƿH�� տ���2��/�h�S� ��wϰϛ��Ͽ���
� ��.��R�=�v�aߚ� �ߗ��߻������� <�'�L�r�]���� �����������8�#� \�G���k��������� ������"F1j Ug������ �B-fQ��u���h�MKCFG ����/�#�LTARM_��
7"0�0N/|V$� METPUᐶ�3����ND� A�DCOLp%A {.C7MNT�/ �%� ����.E#>!�/|4�%POSCF�'=�.PRPM�/9�ST� 1��� {4@��<#�
1 �5�?�7{?�?�?�? �?�?�?)OOO_OAO SO�OwO�O�O�O�O_��A�!SING_C�HK  �/$M/ODAQ,#�����.;UDEV 	���	MC:o\HOSIZEᝢ��;UTASK %���%$123456�789 �_�U9WT�RIG 1���l3%%��9o��"ocoFo�5#�VYP�QNe���:SEM_INF �1�3' �`)AT&F�V0E0po�m)��aE0V1&A3�&B1&D2&S0&C1S0=�m)ATZ�o;"t�H?g�a[o�xA���z����  �o>��o'��K �������я:� L�3�p�#�5���Y�k� }������$�[�H�� �~�9�����Ưد�� ������ӟ�V�	�z� ������c�Կ����
� �.���d��)�;� �Ͼ�q�������˿ <���`�G߄ߖ�IϺ� m�ϑϣ����8�J� ��n�!ߒ�M�����|��h_NITOR� �G ?�[   	EXEC1��/�25�35�45�5�5��P7�75�85�9�0�Қ�4��@� ��L��X��d��p��|�������2���2��2��2��2���2��2��2��2�23��3��3�@�;QR_GRP_�SV 1��k �(�A�z�4�~��K�������K:z�j]��Q_D��^�PL�_NAME !�3%,�!De�fault Pe�rsonalit�y (from �FD) �RR2�� 1�L6(�L?�,0	l d������ ��//(/:/L/^/ p/�/�/�/�/�/�/�/ZX2u?0?B?T?f?@x?�?�?�?�?\R<? �?�?O O2ODOVOhO�zO�O�O�OZZ`\R�?�N
�O_\TP�O:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHo_)_~o�o�o�o �o�o�o�o 2D Vhz�[omo�� ��
��.�@�R�d��v���������Џ�� Ef  Fb�� F7���  G ��!��d� �@�R�6�t����獀�l���ʝ����� ݘ����"�@� F�d���� "𩯹�ݐA�  ϩU[�$n�B�oE �� �� @D�  �?��� �?�@��A@��;f��FH� ;��	l,�	 �|��j�s�d�>���� ��� K(���Kd$2K ���J7w�K�YJ˷�Ϝ�J�	�ܿ�� @I����_f�@�z���f�γ��N������	X�l������W�S�ĽÔ��I �����5����  ����A?o�i#�;����� ���l� �Ϫ�-���ܛG�G�jѲ��@n�@�a   � � ��ܟ*�͵	�'� � H��I� �  y�Рn�:�Èl�?È=��̈́�в@�ߚЕ����D/�����̷NP�  ',���-��@
�@���?=�@A���B��  Cj�a�B�e�Ci��#�B�и�ee��^^ȹBР��P�����̠�����ADz ՟�n�3��C�i�@��R�R�Y����  �@� ��Ż����?�ff������n� ɠ#ѱy 9G
(���I�(�@u�P~����t�t���>�����;�Cd;���.<߈<��g�<F+<L �������,�d�,��̠?fff?��?�&&��@��@�x��@�N�@���@T�H �ِ�!-�ȹ�|� �
`������� //</'/`/r/]/�/��eF���/�/�/��/m?��/J?�(E��G�#�� FY�T?�?P?�?�?�? �?�?O�?/OO?OeO k���O�IQOG�?�O 1?�OmO_0_B_T_������A_�_	_��_�_�_ o��A��A0n0 bФ/o C�_Uo8�_�Op��؃o�o��o�o���W����v�oC�E� q�H�d��؜a@q���e�F�BµWB]��NB2�(A���@�u\?��D�������b��0�|�uR�����
x~�ؽ���Bu*C��$�)`�$� ���GC#����rAU�����1�e�G�D�I�mH��� I:�I��6[F���C��I��J��:\IT�H
?~QF�y��p��*J�/ I�8Y�I��KFjʻCe�o��s� ����Џ���ߏ�*� �N�9�r�]������� �����۟���8�#� \�G�����}�����گ ů���"���X�C� |�g�����Ŀ����� ��	�B�-�f�Qϊ� uχ��ϫ�������� ,��P�b�M߆�qߪ� ���߹�������(�� L�7�p�[����������s($���3�:����$���3Ï��d�,�4���@�R��񴲚�xl�~�wa���e��<��wa4 �{�������(L:ueP�P~�A�O�������	����G2W}h ������/�@��O�O7/m/[(d=� s/U/�/�/�/�/�/?��/1??U?C?y?�= � 2 Ef9gF[b��77�9fB)a,a)`C9A`�&`w`@-o�?w`e�O)O�?MO�Ow`�?�?�O�O��O�O9c?�0�A7hJt4w`w`!w`xn
 �O9_K_ ]_o_�_�_�_�_�_�_��_�_o#ozzQ ���h��G���$�MR_CABLE� 2�h ��a�T� @@��0�Ae��a�a�a���`��0�`C�`�aO�8�tB�n��d��`�aE�4��E�#�o�f#��0��0�DO���By`������bED4�E�c,��o�g8�  ���C�07n�d4
vے�0� �b��XE�Z&�l�`y`
q�C�p�bHE�
v{#g�5D�Ү�qz�lҠ`��0�q�p�b0�
v�%c����b=%	E;h��u/o�c-��4t H�\�?�9�K�]�o�ԏ Ϗ��
�ɏۏ@���?�:�eo �a����������b����� �����`�	 ����@������%� �*�0�6� ��ݐ�����`��	������@������*�,� ,�-�\cOM ��ii��3�� � $Q��%% 23456�78901i�{� �f�����������1�����
��`��not sen�t3�����;��TESTFEC�SALGR  eH�qiG�1d.�š
:�� �DCbS�Q��c�u��� 9UD�1:\maint�enances.Gxml��ֿq� �=��DEFAULT-��4\b�GRP 2�M� � =��a�{�p  �%Fo�rce�sor check  ��
�b�z��p����h5-[ �ϻ������ϖ��D�%!1st c�leaning �of cont.� v�ilatiCon��}�Rߗ+��@[�ߔߦ߸����mech�cal,`������0��h5k�@�R�d�v������(�rolle _Ƶ����/����(�:����Ba�sic quarterly��������,����������M�F�M��:C@"Gp P�a�b`�4��� ����#C���M"��{Pbt����Supp~q�grease���?/&/8/hJ/\/��C+ ge��_. batn�y`/��/h5	/�/�/�/`? ?_�ѷen'�!v��/�/��/��?`�?�?�?�?�G=?O�qp"CrB1O��0�/`OrO�O�O�O�Xt$��Lf��C-m��A�O:�OO$_6_H_�Z_l_�t*cabYl�Om���S<m��Q�_:�
_�_�_o o0oo)(Ӂ/�_�_���_�o�o�o�o�o�;O@hau1�l�2r xm�<qC:��op�������ReplaW�f Uȼ2�:�._4� F�X�j�|�m�$%��� o�������#���
�� .�@���d���ŏ׏�� ��П����U�*�y� ����r���������	� q��?�߯c�8�J�\� n���ϯ�����ڿ)� ���"�4�Fϕ�jϹ� ˿������������ [�0�ϑ�fߵϊߜ� ������!���E�W�,� {�P�b�t����߼� ����A��(�:�L� ^������������ �� $s�H���� ��q�����9 ]o�Vhz� ��U�#�G/ ./@/R/d/��/�/� �//�/�/??*?y/ N?�/�/�?�/�?�?�? �?�???Oc?u?JO�?�nO�O�O�O�O+J�r	 H�O�O__6M2_ @OBE:_p_>_P_�_�_ �_�_�_ o�_�_oHo o(oZo�o^opo�o�o��o�o�o �o :z� �bA?�  @�q _����Fw�� �H* �** @q>v�p 2T�f�x�:�������ҏ��eO^C7�Տ #�5�G�	�k�}���ُ ���c�����W�� C�U�g���ß)����� ӯ���	��-�w��� ��9�������m�Ͽ���=�O�E	A�$�MR_HIST �2�>uN�� 
� \$�Force se�nsor che�ck  1234?567890q�3�����ß�N�}SB� -3�19.8 hou�rs RUN 9�.�Y�!1st �cleaning� of cont�. ventilation0Äϖ�Ԩ�-�Y���me;ch��cali�%���4��o�DN��t��95��1�|���rolleh��+�=�O��Y�B�asic qua?rterlyߒ� �߶�
O4�F��(�� ����b�t������ �����M�_����:�����p���:�SKCFMAP  >u�Q��r5�������ONREoL  .��3���EXCFEN���:
��QFN�CXJJOGOVLIM8dNá ��WKEY8��_PAN7����ԧ�����SF?SPDTYPxC���SIG�:��TO1MOT�G���_CE_GRP [1�>u\�D �����/Ⱥ� �/�/U//y/0/ n/�/f/�/�/�/	?�/ ???�/c??\?�?P? �?�?�?�?�?O)OO�MO,���QZ_ED�IT5 )TCO�M_CFG 1����[�O�O�O 
>�ASI �y3�!
__+[_O_ċ�>O�_bHT_/ARC_Uք�T_MN_MOD�E5�	UAP�_CPL�_gNO�CHECK ?^�� �� o .o@oRodovo�o�o�o �o�o�o�o*!�NO_WAIT_�L4~GiNT�A���EUwT_ERMRs2���3��Ʊ J�����>_)�V�|MO�s��}x:O�v���8�?������ l��rPA�RAM�r�����j���5�5�G� =  r�b�t�s� X������������֟0�0����b�t������SUM_RSPACE�����Aѯ�ۤ�$ODRDS�P�S7cOFFS?ET_CARt@�_��DIS��PE?N_FILE:�7��AF�PTION�_IO��q�M_�PRG %��%�$*����M�WOR�K �yf '��춍�@��� � �������	 �������It��RG_DSBL  ���C�{u��RIE�NTTO7 ��Cٴ A �UT�_SIM_Dy����V�LCT ��}{B �٭�ď_PEX�P=��R[AT�W dc�>�UP ���`���e�w�]ߛߩ���$�2r�L�6(L?���	l d������ &�8�J�\�n���� �����������"�4�F�X���2�߈����� ��������*�<w�Tfx��������J`�ˣG���Tz�Pg���� ��/"/4/F/X/j/ |/�/�/�/���/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?�/�/ ,O>OPObOtO�O�O�O �O�O�O�O__(_:_��O��y_�]2����_�^�_�_�W^]@^]��/ooSog�� Hgrohozo�o�o�o�o��oF`�#|`�AG�  9y����OK��1�k�����<��EA�nq @D�  �q����nq?��C��s�q1�� ;�	l��	 '|�Q�s�r�q>��u
��qF`�H<zH~��H3k7GL�z�HpG�9�9l7�k_B�T�F`C4T��k�H���t��-��Ae���k������s���  ��ሏ����EeBVT����dZ��g���ڏ ����q-�Fk�y�{FbZU���n@6�_  ���z��Fo��Be	'� �� ��I� ��  �:p܋=����ڟ웆�@���B�,���B��g�AgN���� � '|���g��B�*��p�BӀC׏�����@  #�B�u�&�ee�^^މB:p2����>�m�6p�Z���Dz ?o}�܏������׿�������Ǒ��� f� � � �M���*�?�ff�_8�Jφܿ 3pϑ�ñ8@�Чϵʖq.·�(����P���'��s�tL��>��/�;�Cd;���.<߈<��g�<F+<AL ��^oiΚrd@�|�r6p?fff?��?&�п�@���@x��@�N��@���@T� ��Z���ћtމ�u�� �w	�x��ti�>�)�b� M��q��������� ����:�%�^��������W���S�E�  �G�aF�� Fk���������1 U@yd���� ��q��	��{�A ��h�����a��ird��A{/w�/J/5/n/vA��A0���":t�/ C^/�/xZ/ ލ?���/��/1??���W���t�g��pE� ~1��?04�0
1�1@�IӀ��BµW�B]�NB2�(�A��@�u\�?����������b�0�|�uR�����
�>��ؽ��Bu�*C��$�)`��? ���G�C#���r�AU����1��eG���I�m�H�� I:��I�6[F����C4OI���J�:\IT��H
~QF�y��Ol@�*J�/� I8Y�I��?KFjʻC��-? �O�O__>_)_b_M_ �_�_�_�_�_�_�_o �_(oo%o^oIo�omo �o�o�o�o�o �o$ H3lW�{� ������2�� V�h�S���w�����ԏ �������.��R�=� v�a�������П���� ߟ��<�'�`�K�]� ��������ޯɯ��&�8�#�\��3(J��g�3:a������J�3��c4�������������1��㚅ڿ��1����e���14 �{ 2�2�r�`ϖτϺϨ�J�%PR�P���!��h�!�K�6�o�Z�����u�|ߵߠ��� �������3��W�B� {�f�4���������d�A����!��1�3� E�{�i��������������  2 Efn�7Fb�7��6�B�!�!� C9� �� �0@�/`r������#x��+=�3?, V�8�v��0�0�:�0�.
 D� ����//%/7/�I/[/m//�/�:� ���ֻ�G����$PARAM_M�ENU ?2���  �DEFPUL�SE�+	WAI�TTMOUT�+�RCV? S�HELL_WRK�.$CUR_ST�YL� 4<OP9TJJ?PTB_?Y2�C/?R_DECSN 0�Ű<�?�?�?�? �?OO?O:OLO^O�O��O�O�O�O�!SSR�EL_ID  �.�����EUSE_PROG %�*q%�O0_�CCCR0��B���#CW_HOSoT !�*!HT�_=ZT��O_�Sh_zQ��S�_<[_TIM�E
2�FXU� GD�EBUG�@�+�CG�INP_FLMS�Ko5iTRDo5gP+GAb` %l�tk�CHCo4hTYPE
�,� �O�O�o# 0Bkfx�� �������C� >�P�b���������ӏ Ώ�����(�:�c��^�p�����7eWOR�D ?	�+
 �	RSc`��P�NS��C4�JO�v1��TE�P��COL�է�2��gLVP 3�����Oj�TRACECTL� 1�2��!{ Ѐ ��Қ�q�DT Q�2�Ǡ��D �� :��f��Ԡ�Ԡ���}�ׯ���;�4��4��4� ��;�u:�q:���;�U8�	8�
8�8�U8�8�8�8�T�@:�8�8����� ���ٱ޴���ؿ�$�6��� 
�l�~�@�R�dϞϰ� ��������
��V�h� zߌߞ߰��������� 
�,�>�P�*�<�v���*���; (�8� )��*��+ ����������1�C� U�g�y����������� ����	-,�>�P� b�t������������ С�*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6@ubt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀�V�߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h?�z?�?�?�?�?�1�$�PGTRACEL�EN  �1  ���0���6_UP �/���A@�1�@�1_CFG7 �E�3�1U
@�<D�0<D�ZO<C�0uO$BDEF�SPD �/L��1�0��0H_C�ONFIG �\E�3 �0�05d�D��2 �1�AaPpDsA�A�0��0�IN'@TRL ɽ/MOA8pEQPEv�E��G�A�<D�AILID(C��/M	bTGRP 1}ýI l�1�B  ������1A�33FC�� F8� E�� @eN	�A�AsA�Y��Y�A�@� 	 �vO�Fg�_ ´8cokB;`baBo,o�>oxobo�o�1>о�?B/�o�o~��o =%<��
C@yd ��"������  Dz@�I�@A 0�q� �������ˏ�� �ڏ���7�"�4�m��X���|���Ú)ґ�
V7.10be�ta1HF @�����Aq�ܢQ  �?�� �BܠP�p �C���&�B�EQ�A���Q�P�Q�� @ß[�m����<CA���0�b�@���f�������ҡ�R�ܣ�R����1�i������t<B!CeQ�KNOW_M  �lE7FbTSV ĽJ�BoC_�b� t�������������1��]aSM�SŽK ���	NB�0����ĿK���-�bb��A�R� �P����0�Ŗ��bQ+MR�S��T�iN�`��d���V]ST�Q�1 1�K
 4aMU�iǨj� K� ]�oߠߓߥ߷����� ��2��#�h�G�Y�� }�������
������,�27�I��1�#<t�H��P3^�p�����,�4���������,�5(:,�6 Wi{�,�7����,�8�!3n,�MAD�6 F�,�OVLD  �KD�xO.�PAR?NUM  �MC\/%�SCH� E�
9'!G)�3Y%UP�D/��E�/P�_C�MP_��0@�0'�7E�$ER_CH�K�%5H�&�/�+RqS���bQ_MO��+?=5_'?O�_RES_G6��:�I�o �?�?�?�?O�?O7O *O[ONOOrO�O�O�{4]��<�?�Oz5�� �O__|3 #_B_G_ |3V b_�_�_|3� �_ �_�_|3� �_�_o|3�Oo>oCo|2V 1��:�k1!�@c?��=2THR_IN�Rc0i!}�o5d�fM�ASS�o Z�gM�N�o�cMON_QUEUE �:ը"�j0��O�N� U�1Nv�+DpEND8Fqd?`yEXEo`uƅ BEnpPAsOP�TIOMwm;DpPR�OGRAM %�$z%Cp}o(/BrT�ASK_I��~O?CFG �$���K�DATA��&T���j12/ď ֏������+�=�O� a����������͟���INFO�͘�� 3t��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����
�Θ� '��FJ�a K_N��T��˶�ENBg ڽw1��2���GN�2�ڻ� P(O�=�{��]ϸ�@���v� �u�uɡd�Ʒ_EDIT ��T�����G�WER�FL�x�c)�RGA�DJ Ҷ�A�  $�?j00��a��Dqձӆ5'�?��ʨ�<u�)�%e������FӨ�2Y�R��	H;pl�G��b_�>�pAodɻt$�*�/� **:�j0�$�@�5Y�T���^��q�߈b~�L��\� n���������� �����4�F�t�j�|� ������������b LBT�x�� ��:��$, �Pb���/� ���/~/(/:/h/ ^/p/�/�/�/�/�/�/ V? ??@?6?H?�?l? ~?�?�?�?.O�?�?O O O�ODOVO�OzO�O _�O�O�O�O�Or__ ._\_R_d_�_�_�_�_�_�_�f	g�io�pWo �o{d�o�~o�ozo�B�PREF S�Rږp�p
�?IORITY�w[�}��MPDSP�q���pwUT6����OoDUCT3������OG��_T�G��8��ʯrTOE�NT 1׶� �(!AF_IN�E�p,�7�!t�cp7�_�!u�dN���!ic�mv��ޯrXYK��v����q)� ,�����p��&�	� �R�9�v�]�o����� П������*��N�`�*�sK��9}�ߢ�\��Ư ,�/6�H�������خ�At�?,  �Hp���P�b�t����u�w�HANCE �R��:�wd��连�2s��9Ks��POR_T_NUM�s�p����_CAR�TREP{p�Ω�SoKSTA�w dʷLGS)�ݶ���tӁpUnothing��������{��TEMP �޾y��'e��_a_seiban�o \��olߒ�}߶ߡ��� ������"���X�C� |�g���������� ���	�B�-�f�Q��� u������������� ,<bM�q� ������(|L�VERSIyp��w} di�sabledWS�AVE ߾z	�2600H76%8S?�!ؿ����/ 	5(�r)og+^/y�e{/�/�/��/�/�*�,/? ��p���_�p 1��Ћ� ������Wh?z?�W*pURGE��B�p}vgu6,�WF�0DO�vƲ©vW%��4(�C�WR�UP_DELAY� �\κ5R_HOT %Nf�q׿�GO�5R_NORM�AL&H�r6O�OZGS�EMIjO�O�O(qQ/SKIPF3��W3x=_98_J_\_] �_�_{_�_�_�_�_�_ �_	o/oAoSoowoeo �o�o�o�o�o�o�o +=aOq�� ������'���7�]�K�������)E�7$RA{���K/��zĀÁ_PARA�M�A3��K @�.�@`�61�2C�<��y��C��6$�BÀBTIF��4`�RCVTMO�Uu�c��ÀD�CRF3��I ��+UC�AqD���2=\�(�?��]�
�ޅ���4��+_����;�Cd;���.<߈<�g��<F+<L�A��Ѱ��d�u�L� ������ϯ�����)�;�M�_���RDI�O_TYPE  �M=U�k�EFPO�S1 1�\�
 	x4/�����+� $/<��$υ�pϩ�D� ��h��ό��'����� �o�
ߓ�.ߤ�Rߌ� ������5���Y��� i��*�<�v���r��� �������U�@�y�� ��8���\������������?��c����2 1�KԿX��T�x��3 1� ����nY�S4 1�'9K��/�'/�S5 1���/�/�/|�/:/S6 1�Q/�c/u/�/-??Q?�/S7 1��/�/
?D?��?�?�?d?S8 1�{?�?�?�?WOBO{O��?SMASK 1�L��O�D�GXN�O���F&�^��MOCTEZ�Ż��Q_ǁ��%]pA݂��PL_RANG!Q]�_QOWER �ŵ��P1VSM_DRYPRG %ź�%"O�_�UTART� �^�ZUME_PRO�_�_4o���_EXEC_EN�B  ��#�e�GS�PD`O`WhՅjbT3DBro�jRM�o�h�INGVERSI�ON Ź�#o�)I_AIRPURhP �O(�M�MT_�@T�P#_�ÀOBOT_ISOLC�NTV@A'q�huNAME�l���o�JOB_ORD_NUM ?�X�#qH76�8  j1Zc@n�r
�rV�sw��r�?�r�?�r�pÀPC�_TIMEu�a�x�ÀS232>R1��� LTE�ACH PENDcANw�:GX��!O Maint�enance C�onsj2����"���No UseB�׏������1�8C�y�V�NPO�P@��YQ�cS�C7H_L`�%^ ��	ő��!UD�1:럒�R�@VA#IL�q@�Ӏ�J�Q�SPACE1 2�ż ��YRs�i�@Ct�YRԀ'{��?8�?��˯ ����"���7�2�c� u�����G���߯ѿ� ���(��u�AC�c� u�����Ͻ�߿���� ���(��=�_�qσ� ��C߹������߱�� $��9�[�m�ߑߣ� Q������߭��� ��� 	�W�i�{���M��� ����5���.S� e�w�����I����� ��*?as ��E����� /&//;/]o�� ����/2/�/?"? �/7?Y/k/}/�/�/O? �/�/�?�?�?O0OO~KA��*SYPp�M*�8.302�61 yB5/21�/2018 A� �WPfG|�H�_�TX`� !$C�OMME��$USAp �$ENABLED�Ԁ$INN`QpI�OR�B�@RY�E_�SIGN_�`�AP��AIT�C�BWRKz�BD<�_TYP�CRINDXS�@W��@%VFRI{�_G�RPԀ$UFR�AM�rSRTOOL�\VMYHOL�A�$LENGTH_�VTEBTIRST��T  $SE�CLP�XUFINV�_POS�@$�MARGI�A$�WAIT�`�ZX2l�\�VG2�GG1�AAI�@�S�Q	g�`_WR��BNO_USE_�DI�BuQ_REQ��BC�C]S$CUR_TCQP�R"a^f� �GP_STA�TUS�A @ ��A3`�BLk�H$�zc1�h�P@���@_��FX �@E_MLT_CT�C�H_�J�`CO�@O�L�E�CGQQ$W��@w�b#tDEA�DLOCKuDELAY_CNT�a�3qGt�a$wf �2 R1[1T$X<�2[2�{3[3$Zwy�q%Y�y�q%V0�@�c�@�b$V�`�R�V�UV3oh>b�@� � �d�0arMSKJ�LgWaZ�C`�NRK�PS_RATE�0$���S
`�Qv�TAC��PRD��$�e�S*��a4�A�0:�DG�A 0�P�f�lp bquS2�ppI�#`
`�P 
��S\`  ؾA�R_ENBQ ��$RUNN�ER_AXI�<`A�LPL�Q�RU�THI�CQ$FLIP�7��DTFEREN|��R�IF_CHS�U�IW��%V)�G1�����$PřA�Q�Pnݖ_JF�PR_P��	�RV_DA�TA�A  =$�ETIM���_$VALU$�	��OP_   ��A  2 ��SC*�	�� �$ITP_0!�SQ]PNPOU}�o��TOTL�o�DSP>��JOGLIb��P'E_PKpc�Of�i���PX]PTAS��$KEPT_MI�R��¤"`M�b�A	Pq�aE�@�y�q��g@١c�q�PG�BCRK6�x���L�I��  ?�SJ�q�P��ADEz�ܠBSO�Cz�MOTNv�D�UMMY16Ӂ�$SV�`DE_O�P��SFSPD_�OVR
���@L�D����OR��TP8�LE��F������OV��SF��F����bF�d�ƣ&c)�fQ~c�LCHDLY��RECOV���`���W�PM��gŢ�ROȲ�����_F�?� �@v�S �NVER\�@�`OFS�PC,�CSWDٱc�ձ���B,����TRG�š�`�E_FDO��MB�_CM}���B��BALQ�¢	�Q�̄VzaF�BUP�g��G
��AM���@`KՊ�fe�_M!�d�AMf�<Q��T$CA����uDF���HBKd��v���IOU��I'R��PA�����������p��і�DVC_DB�S!�x�Q�!�s�Dd�9�1A��9�3A�^��ATIO�0���͠��US����WaAB��R+c�`tá`Dؼ�A��_AUXw�S�UBCPUP���S �`����3Եжc����3�FLA�B�HW�_Cwp"�Ns&�]sA�a��$UNIT�S�M�F�ATTR�Iz�Z�CYCL��CNECA���F�LTR_2_FI~��TARTUPJp0����A��LP����ޖ�_SCT*cF_�F�F_P���b�FS8��+�K�CHA/Q��p*�d�RSD��`Q����Q���_TH��PROr���հEM�PJ���G�T�c �Q�DI�@~y�RAILAC/��bMX�LOf�xS���ځ���拁���P�R#�S`app�C�� 	��FUsNC���RIN``QQP� ԱRA)]R ��AƠ��AgWAR֓��BLZa�WrAkg�ngD�AQ�B�rkLD@�र&q�M�K����TI���j���$�@RIA_SWV��AF��Pñ#���%%�p9r1��MO9IQ���DF_~P(��PD"LM-�FA��PHRDY�DORG�H; _QP�s%MULSE~Pz���**�� J��Jײ���FAN_ALMsLVG��!WRN�%�HARDP��UcO��� K2$SHADOW]�kp�a02��N� STOf�+�_^�w�AU{`R��eP_SBR�z5���:�F�� �3MPIN�F?�\�4��3R3EGV/1DG�+c1Vm �C�CFL(��?�DAiP���Z`Ɨ� �����Z�	 ��P(Q$�A$�Z�Q V�@�[�
7� ��EG��o����kAAR���㌵2p�axG��AXE��wROB��RED���W�QD�_�Mh�SY�A��AF��FS�GWRqI�P~F&�STR��(��E�˰EH�)��D�a\2kPB6P��=V���Dv�OTO�1)���ARYL�tR��v�3���FI&�ͣ$LINKb!\��Q%�_3S���E�N�QXYZ2�Z5�V'OFF���R�R�X%xPB��ds�G�cFI�03g�h������_J���'�ɲ�S&qR0LTV[6����aTBja�"�bCL���DU�F7�TUR� X��e�Qb�2XP�ЊgFL�@E���x@�`�U9Z8��^�� 1	)�K��	Mw��F9��劂����ORQj��G;W3���#�Ґd ���upz����1�tOVE�q_�M��ё?C�uEC�u KB�v'0�x-�wH��t ���& `��qڠ� B�ё�u�q�wh�ECh�L���ER��K	�!EP����AT�K�6e9e�W���AXs�'��v�/�R  ����!�� ��P ��`��`�3p�Yp�1�p�� �� � � (�� 8�� H�� X� � h�� x�� ������oDEBU�$`%3�I��·RAB�ȱ�ٱ�sV��� 
d�J、��@񘧕� ������Q���a���a ��3q��Yq+$�`%"<�.cLAB0b�u��'�GRO���b<��B_s��"Tҳ*`��0A�u��uq�p1}�ANDGp�������U��p1�� �ѷ0�Qθu�ݸ��PNT0����SERVE �Z@� $`EAV�!�PO����nP!��P@�$!Y@ w $>�TRQ�b�
=��BG�K�%"2�\��� _ � l��5�D6ERRVb(�I��V0`;���'TOQ:�7�L�@
�(R��e G�%�Q��q <�50F� ,��`�z�>�RA� �2 d!�����S�  M��px�U ����OCuG��  ��COU�NT6Q��FZN_wCFGF� 4#��6��TG4�_�=�����(���VC ���M �"��$6��q ��FA E� &��X�@�������A�����AP��P@H�EL�0��� 5b`B_BASN��RSR�6�C�SH����1�Ǌ�2���3��4��5��6ʭ�7��8��}�ROaO����P�PNLEAƭcAB)ë ��AC-Ku�INO�T��(B�$UR0� =�_P�U��!0��OU+�P�d�8j��� V��T�PFWD_KAR���� ��RE(ĉ P��P�>QUE�:RAO�p�`r0P1I� �x�j�P�f��6�QSCEM��0��� A��7STYL�SO j�DIX�&�����S!�_TMCMANR�Q��PENDIt�$KEYSWIT�CH���kHE��`BEATM83PE{@LE��>]���U��F��SpD_O_HOM# O�6@�EF�pPRaB(�A#PY�C� O�!���OV_M|b<0 �IOCM�dFQ���h�HKYA �D�Q�7��UF2��M����p�cFORC��3WAR�"�OM>|@  @S�#�o0U)SP�@1�2�&3&4E��p�S*T�O��L���8OUNLOv�D4K$�EDU1  �S�Y�HDDNF� �M�BLOB  �p�SNPX_;AS�� 0@�0|��81$SIZ�1�$VA{���MU/LTIP-��# �A� � A$��� /4`�BS���0�C���&FRIF�BO�S���3� N=F�ODBUP߰��%@3;9(��ҋ�Z@� x��SI��TE�s�r�cSGL�1T�Rp&�Н3B��@�0OSTMTq�3Pg@�VBW�p�4SHO�W�5@�SV��_�G�� 3p$PC�J�PИ���FB�PHSP AW�EP@�VD�0WC� ���A00��PB �XG XG XG$ XG5�VI6VI7VI8VI9
VIAVIBVI�XG�YF�0XGFVH��XbIU1oI1|I1�I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1Y1Y2UI2bIU2oI2|I2�I2�I@�`�X�I2p�X�I2�IU2�I2�I2�I2Y�2Y�p�hbI3oI3�|I3�I3�I3�I3��I3�I3�I3�I3��I3�I3�I3Y3�Y4�i4bI4oI4�|I4�I4�I4�I4��I4�I4�I4�I4��I4�I4�I4Y4�Y5�i5bI5oI5�|I5�I5�I5�I5��I5�I5�I5�I5��I5�I5�I5Y5�Y6�i6bI6oI6�|I6�I6�I6�I6��I6�I6�I6�I6��I6�I6�I6Y6�Y7�i7bI7oI7�|I7�I7�I7�I7��I7�I7�I7�I7��I7�I7�I7Y7ZT�VP� UD�#y"ՠ��
<A62���t�R��CSMD� ��M5�Rv�,]��Q_h�R���pe����<�YSL��>�  � �%\2 ��+4�'��W�BVALU��b��'�z��FH�ID_L����HI��I���LcE_��㴦�$0�C�SAC�! h� �VE_BL�CK��1%�D_CPU5ɧ 5ɛ ������C�� ��R " � PWj���#0��LA�1S�Bћì���RUN_FLG�Ś����ĳ  ����������H����Х�ցTBC2���# � @ B ��e �S�8=�F'TDC����V���3d�Q�THF�����R�L�ESERCVE9��F��3�2��E��Н�X -$��LEN9��F���f�RA��W"G�WI_5�b�1��д2�MO-�T%S60U�I�k�0�ܱF����[�DyEk�21LACEi�0�CCS#0�� _M�A� j��z��TCV����z�T�������.Bi�'A�z�'AJ$h�#EM5���J��@@Ri�V�z���2Q `�0&@o�h��JK��VK9��{���щ�J0����JJ��JJ��AAL���������4��5�ӕ NA1������.�LD��_�1* �CF�"% `�GRO�U���1�AN4�C��#m REQUIR��EBU�#��6�7$Tk�2$���pzя #�& \�/APPR� C� 0��
$OPEN�C'LOS�St��	ri�
��&' ��MfЩ���W"-_M	G�7CB@�A�ܸ�BBRK@NO�LD@�0RTMO!_5ӆp1J��P��������������6��1�@� | ��#�(�# �����'��+#PATH''@!6# @!�<#� � '��1�SCA���6I�N��UCJ�[1� C0@UM�(Y ��#�"������*���*��� P�AYLOA~J2=LؠR_AN^�3�L��91�)1AR?_F2LSHg2B4LO4�!F7�#T7�#ACRL_�%�0ȏ'�$��H��.�$yHA�2FLEX�u�J!�) P��2�D߽߫���0��* :����z�FG�]D����z���%�F1]A�E�G4�F�X�j�|���BE������ ������(��X�T*� A���@�XI�[�m�\At�T$g�QX<�=�� 2TX���emX������ ������������t+	�J>+ �-�`K]o|�٠AT�F�4�ELFPѪs��J� *� JEmC3TR�!�ATN�v�zHAND_VB�.��1��$, $�8`F2Av���S�Wu8-� $$M*0.�]�W�lg��PZ����A@��� 1����:AK��]AkAz��LTN�]DkDzPZ G��C�ST_K�lK�N}DY��� A ����0��<7]A<7W1@�'��d�@g`�P��������"0C$. M�2D%"�H����ASYM$j%0�� j&-��-W1�/_�{8� �$������/�/�/�/ 3J�<�:9�/�89�D_�VI�v����V_UNI�ӛ��cD1J����╴�W<��n5 Ŵ�w=4��9��?�?$<�uc�4�3��%�H���/�j��0��DIzuO���8�k�>0 �`��I��A��#���@ģ����@��IPl� �1 � /�MEB.Qp��9�ơT}�PT�;pG �+ GtA� ���'��T��0 $DUM�MY1��$PSm_�@RF�@  G �b�'FLA@ Y�P(c|��$GLB_TP�ŗ���p9 P�q��2 X� �z!ST9�� S�BRM M21_V��T$SV_ERb*0O�p����CL�����AGPO��f�GLv~�EW>�3 4H ��$YrZrW@�x�A1+�A���";��"�U&�4 8`N�Z�"�$GI�p}$&� -� �Y��>�5 LH {��}�$F�E��NEA�R(PN�CF��%PT�ANC�B;�JOG܌@� 6.@$JOINTwa?pd��MSET>�7  "x�E��HQtpS{r��|up>�8� �p�U.Q?�� LOC�K_FOV06���B�GLV�sGLt�T?EST_XM� 3�'EMP����Ҏ_�$U&@%�w`24� Y��5��2�d���3��CE- ����_ $KAR�QM��TPDRA)������VECn@��IUھ�6��HEf�TO�OL�C2V�DREN IS3ER6�N�@ACH� 7?1Ox �Q�29Z�H �I�  @$R�AIL_BOXEzwa�ROBO���?��HOWWA�R�1�_�zROLMj��:qw�jq� ��@ O_Fkp!� d�l>�9�� +�R O8B: �@��c�OU�;��Һ�3ơ�r�q_�/$PIP��N&`H��l�@��#@CORDEDd�p >f��fpO�� < D ��OB⁴sd����Kӕ���qS;YS�ADR�qf���TCHt� =� ,8`ENo��1A
k�_{�-$Cq,Be��VWVA��> Ǥ  &��PR�EV_RT�$�EDITr&VSHWRkq�֑ &R:�%v�D��JA�$�a?$HEAD�6�4� �z#KE:�E��CPSPD�&JM%P�L~��0R*P�ģ?��1%&I��S�rC�pNE; �q�wOTICK�C��M�1�<�3HN��@� @� 1Gu�!_GqPp6��0STY'"xLO��:�2l2?�_A t 
m G3%S%$R!{�=��S�`!$��w`���ճ�r��Pˠp6SQU��x�E��u�TERC��Q2�TSUtB ����hw&`gw�Q)b�pO����@IZ��4{��^�PR�kј�B1XPU���E_�DO��, XS�KN~�AXI�@���UR�pGS�r� ^0�d&��p_) �ET�BQPm��o��0Fo�2�0A|���Rԍ���a;�SR�Cl>@P��b_�yU r��Y��yU��yS��yS ���UЇ�U���U���U �]��Ul[��Y�bXk�]Cm�����YR�SC�� D h��DS~0��Q�SPL���eATހ���A�]0,2N�ADDRE�S<B} SHIF�{s��_2CH�pr�I��=q�TVsrI��E"���a�Ce�
��
;�VW�A��'F \��q��0l|\A@�rC�_B"R{z�p�ҩq�TXSCWREE�Gv��1TINA���t{�����A�b?�H T 1�ЂB�����I��Ap��BE�y RRO������� B��D��UE�4I �g�!p�S���RSM]0�GU�NEX(@~Ƴ�j�S_S�ӆ��Á։񇣣��ACY�0� 2-H�pUE;�J���\��@GMT��Lֱ��A��O	�BBL�_| W8���K �Լ0s�OM��LE�/r��� TO!�s�RwIGH��BRD
�%qCKGR8л�T�EX�@����WIDTH�� �B[�|�<���I_��Hi� OL 8K���_�!=r���R:�_��HYґ��O6q�Mg0I紐U��h�Rm��LUMh��FpE#RVw��P���`��N��&�GEU�R��FP)�)� LIP��(RE%@�a)ק@�a�!��f �5�6�7�8Ǣ#B�à�@���tP�fW�Sv@M�USR&�OO <����U�Qs�FOC)��P�RI;Qm� :���T�RIP�m�U)N����Pv��0���f%��'���@�0 qQ����AG �0aT� �a>q�OSт%�RPo���8�R�/�A�H�L4����U¡�SU�g��¢5N��OFF���T��}�O�� 1R������S�GUN���6�B_SUqB?���,�SRTN��`TUg2��mCOR�| D�RAUrPE�T<Z�#'�VCC��	3�V AC36MgFB1f$c�PG ��W (#��AST�EM�����0P�E��T3G�X �<\ ��MOVEz�<���AN�� ���M�>��LIM_X��2� ��2��7�,�����ı�
��VF�`E�� �}��04Y��IB(�7���5S��_Rp� x2��� WİGp+@��}СP��3�Zx ���3A���A�ݠCZ��DRID����V�y08�90� De�MY_UBYd���6�ш@��!��X��P�_S��3��L�KB�M,�$+0DEY�(#EX`�����UM_MU� X����ȀCUS�� ���G0`PACI���а@�Հ:��:,�:����R!E/�3qL�+��:z[��TARG�БP�r��R<�\C d`��A��$�	���AR��SW2 ��-I��@Oz�%qA7p�yREU�U�01�,��HK�2]g0��qP� N� �EAM0GWOR����MRCV3�^ ����O�0M�C�s	p���|�REF_� ��x(�+T� ����������3_RCH4(a�P�І��hrj�NA�5��0�_ ���2����L@��n�@@OU~7w6����Z��a2[��RE�p�@;0\�c�a'2]K�@SUL��]���C��0�^��� NT��L�3��(6I�(6q�(3� L��Q5��Q5(I�]7q�}�Tg`4D�`�0.`0�AP_�HUC�5SA��CMPz�F�6�5�5�0_�aR��a�1I\!�X�9|"GFS��a/d ��M��0p�UF_x��B� ���,RO��Q��'����UR�3GR�`.�3AIDp���)�D��;��A��~�IN��H{D���V@AJ���S͓UWmi=������TYLO*�5�����bt +��cPA� �cCACH�vR�UvQ��P�Y��p�#CF�I0s�FR�XT���Vn+$HO����P!A3� ��XBf�(1 ���$�`�VPy� ^b_SZ�313he6K3he12�J�eh chG�chWA��UMP�j��IMG�9uPAD�iiI�MRE�$�b_SI�Z�$P����0 ��A�SYNBUF��V�RTD)u5tqΓOLE_2DJ�Qu5RJ��C��U��vPQ�uECCUlVE�MV �U�r�WVIR9C�aIuVTPG����rv1s��5qMPLAHqa��v�V0�cm}� CKLAS�q	�Q�"��d  ��H�%ӑӠ@}¾�$�Q���Ue |�0!�rSr�T�#0! �r��iI��m�vK�BGf��VE�Z�PK= p�v�Q�&�_HO�0>��f � >֦3x�@Sp�SLOW>��RO��ACCE0���!� 9�VR�#���p:���AD�����PAV�j�� D�����M_B"���^�J�MPG ��g:�#E$SSC��x&�vP$q��hݲvQS�`qV�N��LEXc�i# T`�sӂ��Q��FLD �DEsFI�3�02���:���VP2�Vj� ��A��V�4[`MV_PIs��t����A�@��FI��|�Z ��Ȥ�����A���A���~�GAߥ1 LOO��1 JCB���Xcx��^`�#PLANE��R��1F�c�����pr�M� [`�噴��S����f����Af��R��Aw�״tU��pR�KE��d�VANCp�A���� k��q�ϲ�BR_AA� l��2� ��p�#Hć�m h���O !K�$������kЍ0SOU&A�"A�
pցpSK�TM@FVI=EM 2l ��P=���n <<��d^K�UMMYK1P�j�`D�ȟ��CU��#AU��o� $��TIT��$PR����OP����VSHIF<�r�p`J�Q�sԙ�fOxE$� _R�`U�#����s�� q������G�"G�޵r'�T�$�SCO{D7�CNTQ i�l�> a�-�a�;�a�H�a�V�P��1�+�2u1���D����  D��MO�Uq��a�YJQ�����a_�R�[�r�n�*@LIxQ�AA/`�XVR���s�n�TL���ZABC�t�t�c��
L�ZIP��u,���LVbcLn"�{ ��MPCFx�Mv:�$�� ���?DMY_LN����8���@y�w Ђ(a\�u� MCM�@Cbc�CART_�DP~N� $J71D��=NGg0S�g0�BUXW� ��U�XEUL|B yX���	������x 	���m��YH�Db  y� 80���0EIGH�3n�?(� H��9��$z ���|�,����$B� Kd'���_��L3�RVS�F8`���OVC�2@'�$|�>P&��
q�4��5D�TR�@ �9Vc��SPHX��!�{ ,� *<��$R�B2 2 ����C!�  ��� V+L�b*c%g!`+g"��`V*�,8�?�V+�/V.�/�/ ?�/�/V(7%3@/R/ d/v/�/6?�/�/�?�?@�?O4OOION;4]? o?�?�?�?SO�?�?�O�_�O0_Q_8_f_N;5 zO�O�O�O�Op_�O_ o8o�_MonoUo�oN;6�_�_�_�_�_�oo %o4Uj�r�N;7�o�o�o�o�o�  BQ�r�5���������N;8����� Ǐ=�_�n���R���şx��ڟN;G � џ�
�� ����W�i�{����� ��ï�.�������A��dW�<�N�|� ������Ŀֿ�ޯ� ��0�B�_�R�d�� �϶������������ �*�L�^��rτ�
� �����������&�p8�J�l�~� `ҟ @����������-����&�,� ��9�{�����a��� ������������A 'Y����� ����a#�1�
��N;_MO�DE  ��S ��[�Y�AB���
/\/*	|/��/R4CWORK_{AD�	��DT1/R  ���� ��/� _INTVA�L�+$��R_O�PTION6 ��q@V_DAT�A_GRP 2,7���D��P�/~? �/�?�9��?�?�?�? OO;O)OKOMO_O�O �O�O�O�O�O_�O_ 7_%_[_I__m_�_�_ �_�_�_�_�_!ooEo 3oioWoyo�o�o�o�o �o�o�o/e S�w����� ��+��O�=�s�a� ������͏���ߏ� �9�'�I�o�]������$SAF_DO_PULS� �~�������CAN_T�IM����ΑR� ��Ƙ/��5�;#�U!P"�1!���  �?E�W�i�{�����.��ïկ�����'(~�T"2F���dR�I�Y��2�o+@a얿����)�u���� k0ϴ��_ ��  T� � ��2�D�)�T D��Q�zόϞϰ����� ����
��.�@�R�d��v߈ߚ�/V凷�����߽��R�_;�o �W��p��
�t���Diz$� �0 � �T"1!��� ������������ ��*�<�N�`�r��� ������������ &8J\n��� �����"4FX ��࿁�� �����/`4� =/O/a/s/�/�/�/�/ �/�/�!!/ �0޲k� ݵu�0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ ok$o6oHoZo lo~o�o�o�o�o1/�o �o 2DVhz �/5?������ ��&�8�J�\�n��� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-��?�Q�c�u��� �� ��`Ò�ϯ���� )�;�M�_�q������� ��˿ݿ� ����\3� ���&2,���	12345�678v�h!B_!��2�Ch���0�ϵ����� �����!�3�9ѻ�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� h�K߰���������
� �.�@�R�d�v����� ���������* <N`r���� ���&��J \n������ ��/"/4/F/X/j/ |/;�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�/�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_�? L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o=_�o�o�o�o�o �o 2DVhz@�����h��� ���u�o.�@�R���Cz  B��_   ���2&�_ � _�
����  	�_�2��Տ����_�p������ďi�{� ������ß՟���� �/�A�S�e�w����� ����N������+� =�O�a�s��������� Ϳ߿���'�9�K�"_������<v�_���$SCR_GR�P 1
� ��� t ���� ��	 �����������������_������)�a�����&�DE� D�W8���l�&�G��CR-35iA �90123456�7890��M-�20��8��CRg35 ��:�
��D�������������:֦�Ӧ�G���&������	��]�o������:���H���>��������@���&���ݯ:���j����g������B��t����������A����  @�`��s@� ( ?�=���Ht�P
��F@ F�`z�y� ����� �$ H��Gs^p��B��7�� /�0//-/f/Q/�/ u/�/�/�/8���P�� 7%?����"?W?-2<?<���]? �H�1�?t�ȭ7@�������?-4A, ��&E@�<�@G�B-1 3OZOlO-:HA��H�O�O|O P��B(�B�O�O_��E�L_DEFAUL�T  �����`SHO�TSTR#]JA7RM�IPOWERFL�  i�/UYTW7FDO$V /UR�RVENT 1�����NU L�!DUM_EI�P_-8�j!AF_INE#P�_-4O!FT�_->�_r;o!��`o �*o��o!RPC_M'AIN�ojh�vo�oN�cVIS�oii��o�!TPpPU��Ydk!
P�MON_PROX	Yl�VeZ�2r���]f��!RD�M_SRV��Yg�O�!R��k��XYh>���!
�`M���\i���!RL�SYNC�-98|֏3�!ROS�_�-<�4"��!
C}E4pMTCOM����Vkn�˟!	��C'ONS̟�Wl����!��WASRCd��Vm�c�!��'USBd��XnR��� Noӯ�������!���E��i�0���WRV�ICE_KL ?�%�[ (%S?VCPRG1��-:"Ƶ2ܿ�˰3�	�"˰4,�1�˰5T�Y�"˰6|ρ�˰7�ϩϐ˰�����9���� ȴf�!�˱οI�˱�� q�˱ϙ�˱F���˱ n���˱���˱��9� ˱��a�˱߉��7� ���_������� ��)����Q����y� �'���O����w� �������� ˰��İd�c��� ���=(a s^������ /�/9/$/]/H/�/ l/�/�/�/�/�/�/�/ #??G?2?k?V?}?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O��O�O�O	_�O-_��_�DEV �Y��MC:5Xd��GTGRP 2�SVK ��bx 	�� 
 ,�PK 5_�_�T�_�_�_ o�_'o9o o]oDo�o hozo�o�o�o�o�o �o5{�_g�� �������� ?�&�c�u�\������� Ϗ���J\)���M� 4�q���j�����˟ݟ ğ��%���[�B� �f������ٯ���� ���3��W�i�P��� t���ÿ���ο�� �A�(�e�L�ί��R� ���ϸ������ �� O�6�s�Zߗߩߐ��� �������'�~ϐ�]� ��h�������� �����5��Y�@�R� ��v���������@�	 ��?&cu\� ������� ;M4qX���� ���/�%//I/ [/B//f/�/�/�/�/ �/�/�/�/3??W?� L?�?D?�?�?�?�?�? O�?/OAO(OeOLO�O �O�O�O�O�O�O�O_�iV �NLy�6� * 		S=>��+c"_VU@T�n_Y_B���B��2�J�j~Q��~_g_�_�Q%J?OGGING�_�^�7T(?VjZ�R{f��Y���/e�_%o7e�Tt�]/o�o {m�_�o�m?Qi�o�o�;)Kq%� �o�}os���� ��9�{`��)��� %���ɏ���ۏ�S� 8�w��k�Y���}��� ş���+��O�ٟC� 1�g�U���y������ �'����	�?�-�c� Q���ɯ����w���s� ���;�)�_ϡ��� ſOϹϧ�������� �7�y�^ߝ�'ߑ�� �ߣ��������Q�6� u���i�W��{��� ���=��M���A�/� e�S���w�������� ����=+aO ������u�� �9']��� M������/ 5/w\/�%/�/}/�/ �/�/�/�/=/"?4?�/ ?�/U?�?y?�?�?�? ?�?9?�?-OO=O?O QO�OuO�O�?�OO�O _�O)__9_;_M_�_ �O�_�Os_�_�_o�_ %oo5o�_�_�o�_[o �o�o�o�o�o�o!co H�o{��� ���; �_�S� A�w�e�������я� ��7���+��O�=�s� a������П���� �'��K�9�o����� ��_���[�ɯ���#� �G���n���7����� ����ſ����a�F� ���y�gϝϋϭϯ� ����9��]���Q�?� u�cߙ߇ߩ���%��� 5���)��M�;�q�_� ���߼��߅������ %��I�7�m������ ]�����������! E��l��5��� ����_D� we����� %
//���=/s/ a/�/�/�/��/!/�/ ??%?'?9?o?]?�? �/�?�/�?�?�?O�? !O#O5OkO�?�O�?[O �O�O�O�O_�O_sO �Oj_�OC_�_�_�_�_ �_�_	oK_0oo_�_co �_so�o�o�o�o�o#o Go�o;)_Mo ����o��� �7�%�[�I�k���� ������ُ���3� !�W���~���G�i�C� ���՟���/�q�V� �����w�������� ѯ�I�.�m���a�O� ��s�������߿!�� E�Ͽ9�'�]�Kρ�o� ������Ϸ���� 5�#�Y�G�}߿Ϥ��� m���i������1�� U��|��E����� ����	���-�o�T��� ���u����������� G�,k���_M� q����� ��%[Im� ��	���// !/W/E/{/��/�k/ �/�/�/�/	???S? �/z?�/C?�?�?�?�? �?�?O[?�?RO�?+O �OsO�O�O�O�O�O3O _WO�OK_�O[_�_o_ �_�_�__�_/_�_#o oGo5oWo}oko�o�_ �oo�o�o�oC 1Sy�o��oi� ����	�?��f� x�/�Q�+���Ϗ��� ��Y�>�}��q�_� ������˟���1�� U�ߟI�7�m�[�}�� ��ǯ	��-���!�� E�3�i�W�y�ϯ��ƿ ��������A�/� eϧ���˿UϿ�Q��� ������=��dߣ� -ߗ߅߻ߩ������� �W�<�{��o�]�� ��������/��S� ��G�5�k�Y���}��� ������������C 1gU������{ ����	?-c ���S���� ��/;/}b/�+/ �/�/�/�/�/�/�/C/ i/:?y/?m?[?�?? �?�?�?? O??�?3O �?COiOWO�O{O�O�? �OO�O_�O/__?_ e_S_�_�O�_�Oy_�_ �_o�_+oo;oao�_ �o�_Qo�o�o�o�o �o'ioN`9 ������A&� e�Y�G�i�k�}��� ��׏���=�Ǐ1�� U�C�e�g�y����֟ ���	���-��Q�?� a���ݟ��퟇��ϯ ��)��M���t��� =���9���ݿ˿�� %�g�Lϋ���mϣ� �ϳ�������?�$�c� ��W�E�{�iߟߍ߯� �����;���/��S� A�w�e��������� �����+��O�=�s� �����c��������� ��'K��r��; �������# eJ�}k�� ���+Q"/a� U/C/y/g/�/�/�// �/'/�/?�/+?Q??? u?c?�?�/�?�/�?�? �?OO'OMO;OqO�? �O�?aO�O�O�O�O_ _#_I_�Op_�O9_�_ �_�_�_�_�_oQ_6o Ho�_!o�_io�o�o�o �o�o)oMo�oA/ QSe�����%{,p�$SER�V_MAIL  �+u!��+q�O�UTPUT��$�@�RV 2��v  $� (�q�}��SAVE�7�(�TOP10 �2W� d O6 *_�π(_� �����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u�����`����Ͽݷ��YP���'�FZN_CFGw �u$��~����GRP �2�D� ,B�   A[�+qD;� B\��  �B4~�RB2�1��HELL�!�u��j�k�2���>��%RSR���� ���
�C�.�g�Rߋ� v߈��߬�����	����-�?�Q��  �_�%Q���_�슨�,p����)ޖ�g�2,pd��ﾆ�HK 1�� ��E�@�R�d��� �������������� *<e`r���?OMM ������FTOV_EN�B�_���HOW_?REG_UI�(��IMIOFWDL� �^�)WAIT���$V1��^�NTIM���VA�_)_UNIT�����LCTRY�B�
�MB_HDD�N 2W�  2�:%0 �pQ/�qL/ ^/�/�/�/�/�/�/�/��"!ON_ALI_AS ?e�	f�he�A?S?e?w?�: /?�?�?�?�?�?OO &O8OJO�?nO�O�O�O �OaO�O�O�O_"_�O F_X_j_|_'_�_�_�_ �_�_�_oo0oBoTo �_xo�o�o�o�oko�o �o,�oPbt �1������ �(�:�L�^�	����� ����ʏu�� ��$� Ϗ5�Z�l�~���;��� Ɵ؟����� �2�D� V�h��������¯ԯ ���
��.�ٯR�d� v�����E���п��� ϱ�*�<�N�`�r�� �ϨϺ���w����� &�8���\�n߀ߒߤ� O�����������4� F�X�j�|�'����� �������0�B��� f�x�������Y����� ����>Pbt ������ (:L�p�� ��c�� //$/ �H/Z/l/~/)/�/�/ �/�/�/�/? ?2?D?�V?]3�$SMON�_DEFPRO ����1� *S�YSTEM*0�m6RECALL �?}9 ( ��}0copy m�db:*.* v�irt:\tmp�back\=>1�47.87.14�9.40:102�96 �6�9517q2]?O+M}4x�2fr:\�?I@�?�1p�?O�O�O }5?EaGOYO�6uO�O_*_�}9@Ds:ord�erfil.dat�?�O�O�_�_.M�? Y_�?t_�_o)o<O�O �_rOo�o�o�OKo]o��O�o%8c
xy�zrate 61 �o�o�o ��6ey?w_192 � q��&�9~���� �����6e��U9308 ^�p�����%�8c8�R�Sout�put\tcpserv3.pc�P�: over =>370278�P357235 �� ����.�@_R_ʏ܀y�
��/l/�_ڟ҉������7d3?oR΍ s����(�;i�oدՆ �������<�N�`�r� ���'Ϻ�̟U�p�� �ϥ�8�J�e�n���� #߶�I�[���Ϗߡ� 4�F�W�j�|���2� D���h��ߋ����� ]���x�	��.�@��� d������,���O�a� t���)<�N����� ����U��p� %8�����n� � ���GY��~/!/ 4�F����/�/�<ď�Q7516ގo/��/?$?7dtpdisc 0�/�!�/��/?�?�?7Ttp?conn 0I�X? j?|?OO2_D��. �?�O�O�_�\O�(pO �O_%_8oK/]/�#�O _�_�_�oM___� u_؇_o*o}<��te�st_Աerټ1�62791424�:263469  �_�o�o2ODO�O�?zo �O�O�o�O�o����|�$SNPX�_ASG 2�����q�� P 0 '�%R[1]@g1.1��y?��s%�!��E�(�:�{� ^�������Տ��ʏ� ��A�$�e�H�Z��� ~���џ����؟�+� �5�a�D���h�z��� ��ů�ԯ���
�K� .�U���d�������ۿ ������5��*�k� N�uϡτ��ϨϺ��� ���1��U�8�Jߋ� nߕ��ߤ�������� ��%�Q�4�u�X�j�� ������������;� �E�q�T���x����� ������%[ >e�t���� ��!E(:{ ^������/ �/A/$/e/H/Z/�/ ~/�/�/�/�/�/�/+? ?5?a?D?�?h?z?�? �?�?�?�?O�?
OKO .OUO�OdO�O�O�O�O �O�O_�O5__*_k_ N_u_�_�_�_�_�_�_ �_o1ooUo8oJo�o�no�o�o�d�tPAR�AM �u��q �	��jP��d9p�ht���pOFT_KB_?CFG  �c�u��sOPIN_SI/M  �{vn���p�pRVQS�TP_DSBW~�r"t�HtSR �Zy � & �ROB195_?SERV M����vTOP_O�N_ERR  �uCy8�PTN �Zuk�A�4�RING_PR��D��`VCNT?_GP 2Zuq�!px 	r��ɍ`���׏��wVD���RP 1�i p �y��K�]�o����� ����ɟ۟����#� 5�G�Y���}������� ůׯ�����F�C� U�g�y���������ӿ ��	��-�?�Q�c� uχϙϫ��������� ��)�;�M�_�qߘ� �ߧ߹��������� %�7�^�[�m���� ����������$�!�3� E�W�i�{��������� ������/AS ew������ �+=Ovs �������/ /</9/K/]/o/�/�/ �/�/�/�/?�/?#? 5?G?Y?k?}?�?�?�?��?�?�?�?OO)�P�RG_COUNT�8v�k�GuKBEN�B��FEMpC:t}O_�UPD 1�{T  
4Or�O�O �O__!_3_\_W_i_ {_�_�_�_�_�_�_�_ o4o/oAoSo|owo�o �o�o�o�o�o +TOas��� �����,�'�9� K�t�o���������ɏ ۏ����#�L�G�Y� k���������ܟן� ��$��1�C�l�g�y� ��������ӯ����	� �D�?�Q�c������� ��ԿϿ����)��;�d�_�q�=L_IN�FO 1�E[�@ �2@����������� �ٽ`�y*�d�h�'��¬��=�`y;MYSDEBSUGU@�@���d�I�f�SP_PASS�UEB?x�LOGW  ���C��9*ؑ�  ��A��UD1:\��<�Υ�_MPC�ݵEH&�8�A��V� �A~�SAV !�ݰ�����X���S�VZ�TEM_TI_ME 1"���@ 0  JX����������$T1SVGUNS�@�VE'�E��AS�K_OPTION�U@�E�A�A+�_D�I��qOG�BC2_?GRP 2#�I�������@�  C����<Ko�CFG %z��� �����`��	�.> dO�s���� ���*N9r ]��������/�8/#/\/n/v$ Y,�/Z/�/�/H/�/? �/'??K?]�k?=�@0 s?�?�?�?�?�?�?O �?OO)O_OMO�OqO �O�O�O�O�O_�O%_ _I_7_m_[_}__�_ �_�X� �_�_oo/o �_SoAoco�owo�o�o �o�o�o�o=+ MOa����� ����9�'�]�K� ��o���������ɏ�� �#��_;�M�k�}��� �����ß�ן�� 1���U�C�y�g����� ����������	�?� -�c�Q�s��������� �Ͽ����)�_� Mσ�9��ϭ������� m���#�I�7�m�� ��_ߵߣ��������� ��!�W�E�{�i�� ������������� A�/�e�S�u�w����� ��������+=O ��sa����� ��9']K mo������ �#//3/Y/G/}/k/ �/�/�/�/�/�/�/? ?C?��[?m?�?�?�? -?�?�?�?	O�?-O?O QOOuOcO�O�O�O�O �O�O�O__;_)___ M_�_q_�_�_�_�_�_ o�_%oo5o7oIoo mo�oY?�o�o�o�o �o3!CiW�� ������� -�/�A�w�e������� ���я���=�+� a�O���s�������ߟ ͟��o�-�K�]�o� ퟓ�����ɯ���צ���$TBCSG_GRP 2&ץ��  ��� 
 ?�  6�H�2�l�V��� z���ƿ��������(�d�E�+�?�	 HC�=���>���G���~�C�  A�.��e�q�C��>ǳ3�3��S�/]϶�Y���=Ȑ� C\  B�ȹ��B���>�c���P���B�Y��z��L�H�0�$�����J�\�n�����@ �Ҿ���������=��Z�%�7����?3������	V3�.00.�	cr;35��	*�����
�������� �3��4�   �{�CT�v�}��J�2�)������C�FG +ץ�'� *������rI���� .<
�<bM�q �������( L7p[�� ����/�6/!/ Z/E/W/�/{/�/�/�/ �/.�H��/??�/L? 7?\?�?m?�?�?�?�? �? OO$O�?HO3OlO WO|O�O����Oӯ�O �O�O!__E_3_i_W_ �_{_�_�_�_�_�_o �_/oo?oAoSo�owo �o�o�o�o�o�o+ O=s�E��� Y�����9�'� ]�K�m�������u�Ǐ ɏۏ���5�G�Y�k� %���}�����ßşן ���1��U�C�y�g� ������ӯ������ 	�+�-�?�u�c����� �����Ͽ���/� A�S�����qϓϕϧ� �������%�7�I�[� ��mߣߑ߳����� �߷��3�!�W�E�{� i����������� ��A�/�e�S�u��� ������������ +aO�s�� e�����'K 9o]���� ���#//G/5/k/ }/�/�/[/�/�/�/�/ �/??C?1?g?U?�? y?�?�?�?�?�?	O�? -OOQO?OaO�OuO�O �O�O�O�O�O___ M_�e_w_�_3_�_�_ �_�_�_oo7o%o[o moo�oOo�o�o�o�o �o!3�o�oiW �{������ �/��S�A�w�e��� ����я������� =�+�M�s�a������� ��ߟ�_	���_ן ]�K���o�������ۯ ɯ���#���Y�G� }�k�����ſ׿���� ����U�C�y�g� �ϋ��ϯ�������� 	�?�-�c�Q�s�u߇� �߫��������)�� 9�_�M����/���� i������%��I�7� m�[������������� ������EWi{ 5������� �A/eS�w �����/�+/ /O/=/_/a/s/�/�/ �/�/�/�/?'?��?? Q?c??�?�?�?�?�? �?�?O�?5OGOYOkO�)O�O}O�O�O�O�N s �@S V�_R�$TBJO�P_GRP 2,��E� / ?�V	-R4S�.;\��@|�u0{SPU >���UT @��@LR	 �C�� �Vf  C����ULQLQ>�33��U�R����U�Y?~�@=�ZC��P׌�ͥR��P � B��W$o/gC���@g�dDb�^���eeao�P�&ff�e=�7L3C/kaB o�o�P��P�efb-C�p��^g`�d�o��PL�Pt<�eVoC\  �Q@�'p}�`�  A�o�L`�_wC�BrD�S�^�]�_�S~�`<PB��P0�anaa`C�;�`L�w�aQoxp��x�p:��XB$4'tMP@�PCHS��n���=�P����trd<M�gE�2pb ����X�	��1�� )�W���c�������� ����󟭟7�Q�;�PI�w���;d�Vɡ��U	V3.00�RScr35QT�*�QT�A�� �E�'E�i��FV#F"w�qF>��FZ�� Fv�RF�~�MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
�D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt���ٵ=�_t��V �R�p�V9� ]ESTP�ARtp�HFP*SH�R\�ABLE 1%/;[%�SG��Q �W�G�G�GȨ WQG�	G�
G��GȖ�QG�G�8G�ܱv�RDI~�EQ�ϧϹ�������W�O_�q�{ߍߟ߱���w�S]�CS !ڄ�� �����������&� 8�J�\�n��������� ���� ]\�`��	� �(�:�����
��.��@�w�NUM  ��EEQ�P�	P ۰ܰw�_CFG 0��)r-P�IMEBF_TT�b��CSo�,VER�ڳ-B,R 1=1;[ 8��R��@� �@&   �������/ /)/;/M/_/q/�/�/ �/�/�/?�/?J?%? 7?M?[?m?>�@�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_l_�Y�@cY�MI_CWHAN8 c c�DBGLV��:�cX�	`ETHER_AD ?f�\`��?�_uo�oQ��	`ROUTV!�	
!�d�o�lSN�MASKQhcba255.uߣ'�9ߣY�OOLOF/S_DIb��U;i�ORQCTRL �2		�Ϸ~T �����#�5�G� Y�k�}�������ŏ׏ �����.��R�V��PE_DETAI�/h|zPGL_CONFIG 8�	����/cel�l/$CID$/grp1V�̟ޟ����Ӏ�o?�Q�c� u�����(���ϯ�� ����;�M�_�q��� ��$�6�˿ݿ��� %ϴ�I�[�m�ϑϣ� 2����������!߰� ��W�i�{ߍߟ߱�%}F�������/�A��C�i�H�Eߞ�� ��������?��.�@� R�d�v���������� ������*<N` r������ �&8J\n� �!�����/ �4/F/X/j/|/�// �/�/�/�/�/??�/ B?T?f?x?�?�?+?�? �?�?�?OO�?>OPO�bOtO�O�O�O����User Vi�ew ��}}12�34567890 �O�O�O_#_5_=T�P,��]_���I2�I:O �_�_�_�_�_�_X_j_�B3�_GoYoko}o�o�o o�op^46o�o�1CU�ovp^5 �o�����	�h*�p^6�c�u����� �����ޏp^7R�� )�;�M�_�q�Џ��p^8�˟ݟ���%����F�L� lCamera�J ��������ӯ���E~��!�3��OM�_�`q��������y  e� �Yz���	��-�?�Q� ��uχϙ�俽���������>��e�5i�� c�u߇ߙ߽߫�d��� ���P�)�;�M�_�q� ��*�<��i������� ��)���M�_�q��� ��������������<� û��=Oas�� >����*' 9K]f�Q��� ����/�%/7/ I/�m//�/�/�/�/ n<��^/?%?7?I? [?m?/�?�?�? ?�? �?�?O!O3O�/<׹� �?O�O�O�O�O�O�? �O_!_lOE_W_i_{_�_�_FOXG9+_�_�_ oo(o:o�OKopo�o )_�o�o�o�o�o 
��	g�0�oM_q ���No����o �%�7�I�[�m�& l�n��Ə؏����  ��D�V�h������� ��ԟ柍�g�ڻ}� 2�D�V�h�z���3��� ¯ԯ���
��.�@� R���3uF�鯞���¿ Կ������.�@ϋ� d�vψϚϬϾ�e�w� ��U�
��.�@�R�d� ψߚ߬��������� ��*���w���v� �������w���� �c�<�N�`�r����� =�w��-����� *<��`r�����������  ��1CUgy��������   -/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E_W_i_�  
���(  �%( 	 y_�_�_�_ �_�_�_o	o+o-o?o@uoco�o�o�o�Z* �Q&� J\n������o ���9�(�:�L� ^�p���������܏ � ��$�6�}�Z�l� ~�ŏ����Ɵ؟��� C�U�2�D�V���z��� ����¯ԯ���
�� c�@�R�d�v������ ��п�)���*�<� N�`ϧ����ϨϺ�� ������&�8��\� n߀��Ϥ߶������� ��E�"�4�F��j�|� ����������� �e�B�T�f�x����� ��������+�, >Pb������� ���(o� ^p������ � /G$/6/H/�l/ ~/�/�/�/�//�/�/ ?U/2?D?V?h?z?�?�/�`@ �2�?�?��?�3�7�P��!�frh:\tpg�l\robots�\m20ia\c�r35ia.xml�?;OMO_OqO�O�O�O�O�O�O�O �� �O_(_:_L_^_p_�_ �_�_�_�_�_�O�_o $o6oHoZolo~o�o�o �o�o�o�_�o 2 DVhz���� ��o�
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟�ݟ� �&�8�J�\�n����� ����ȯߟٯ���"� 4�F�X�j�|��������Ŀ־�8.1 ��?@88�?�ֻ�ֿ�3�5�G� iϓ�}ϟ��ϳ����� ���5��A�k�U�w���߿��$TPGL�_OUTPUT �;�!�! ��������,� >�P�b�t����� ��������(�:�L�@^�p�������������2345678901�������� �"��BTfx� �4�����
}$L^p�� ,>��� //$/ �2/Z/l/~/�/�/:/ �/�/�/�/? ?�/�/ V?h?z?�?�?�?H?�? �?�?
OO.O�?<OdO vO�O�O�ODOVO�O�O __*_<_�OJ_r_�_ �_�_�_R_�_�_oo &o8o�_�_no�o�o�o �o�o`o�o�o"4 F�oT|����\��}�����0�B�T�e�@������� ( 	 �� Џ������<�*� L�N�`���������ޟ ̟���8�&�\�J� ��n���������ȯ���"�������*�X� j�F�����|�¿Կ�� C���ϱ�3�E�#�i� {�忇ϱ�S������� ���/ߙ�S�e�߉� ��y߿���;����� ��=�O�-�s���ߩ� ��]��������'��� �]�o���������� ��E�����5G% W}������g� ��1�Ug	 w�{��=O	/ /�?/Q///u/�/� �/�/_/�/�/�/�/)? ;?�/_?q??�?�?�? �?�?G?�?O�?OIO [O9OO�O�?�O�OiO �O�O�O!_3_�O_i_ {__�_�_�_�_�_�R��$TPOFF_�LIM >�op:���mqbN_�SV`  l��jP_MON M<6�dopop�2l�aSTRTC�HK =6�f�� bVTCOMP�AT-h�afVWV_AR >Mm�h.1d �o �oop�`ba_DEFPROG %|j�%ROB195�_SERV	�j_DISPLAY`�|n"rINST_M�SK  t| �^zINUGp�odtL�CK�|}{QUIC�KMEN�dtSC�RE�p6��btpscdt�q�h�b*�_.�ST�j�iRACE_CF�G ?Mi�d�`	�d
?�u�H_NL 2@|i����k r͏ߏ����'�9�K�]�w�IT�EM 2A�� ��%$12345�67890���� � =<��П�� G !���p�� =��c��^������� ���.���R��v�"� H�ί��Я������ *�ֿ���r�2ϖ��� ��4�޿�ϰ���&��� J�\�n���@ߤ�d�v� �ς������4���X� �*��@������ ��������T���x� ������l������ ��,�>�P�������F X��d������ :�p"��o �����F6H Zt~��N/t/�/ ��// /2/�/V/? (?:?�/F?�/�/�/j? �??�?�?R?�?v?�? QO�?lO�?�O�OO�O *O|O_`O _�O0_V_ h_�Ot_�O__�_8_ �_
oo�_@o�_�_�_ Lodo�_�o�o4o�oXo jo3�oN�or��o���s�S�B|���z�  h���z ��C�:y
 �P�v�]����UoD1:\�����q�R_GRP 1C���� 	 @Cp���$��H�6�l�Z��|�����f�৏˟���ڕ?�  
���<�*�`�N� ��r�������ޯ̯���&��J�8�Z���	��u�����sSCBw 2D� �� ���(�:�L�^�p�����|V_CONFIG E���@�����ϖ�OUTPU�T F�������6�H�Z�l�~� �ߢߴ���������� ��#�6�H�Z�l�~�� ������������� 2�D�V�h�z������� ��������
�.@ Rdv����� ��)<N` r������� //%8/J/\/n/�/ �/�/�/�/�/�/�/? !/4?F?X?j?|?�?�? �?�?�?�?�?OO/? BOTOfOxO�O�O�O�O �O�O�O__+O>_P_ b_t_�_�_�_�_�_�_ �_oo'_:oLo^opo �o�o�o�o�o�o�o  $����!�bt� �������� (�:�-o^�p������� ��ʏ܏� ��$�6� G�Z�l�~�������Ɵ ؟���� �2�D�U� h�z�������¯ԯ� ��
��.�@�Q�d�v� ��������п���� �*�<�M�`�rτϖ� �Ϻ���������&� 8�J�[�n߀ߒߤ߶� ���������"�4�F� W�j�|�������� ������0�B�S�f� x��������������� ,>Pa�t� �������(:L/x���k}gV�K� ��//&/8/J/\/ n/�/�/�/W�/�/�/ �/?"?4?F?X?j?|? �?�?�?�/�?�?�?O O0OBOTOfOxO�O�O �O�?�O�O�O__,_ >_P_b_t_�_�_�_�O �_�_�_oo(o:oLo ^opo�o�o�o�o�_�o �o $6HZl ~����o��� � �2�D�V�h�z��� �����ԏ���
�� .�@�R�d�v������� ��Ϗ�����*�<� N�`�r���������˟ ޯ���&�8�J�\��n���������Ż�$�TX_SCREE�N 1G�g�}ip�nl/��gen.htmſ�*�<�N��`ϽPanel setupd�}�dϥϷ����������ω�6�H�Z�l� ~ߐ�ߴ�+������� � �2�߻�h�z�� �����9�g�]�
�� .�@�R�d������� ��������}���< N`r��;1 ��&8�\ �������Q�ȾUALRM_M_SG ?��� �Ȫ-/?/p/c/ �/�/�/�/�/�/�/?�?6?)?Z?%SEV7  -�6"ECFG I嵻�  ȥ@�  A�1   ;B�Ȥ
 [?ϣ ��?OO%O7OIO[O�mOO�O�O�G�1GR�P 2J�; 0�Ȧ	 �?�O I�_BBL_NOT�E K�:T��lϢ�ѡ��0RDEFPR�O %+ (% N?u_Ѡc_�_�_�_�_ �_�_o�_o>o)obo�Mo�o\INUSE�R  R]�O�oI�_MENHIST� 1L�9  �(_P ��)/�SOFTPART�/GENLINK�?current�=menupag�e,1133,1`�oDVhz~�(
50�����ޛzedit(rONE�I�[�m���	#�OPEN8�Ώ����� �'���~7�1��P�b�t����0����ROB195t0RV?�ݟ����� z37̟X�j�|�0���/�)r95G�ݯ ���6Q�`q|oB� T�f�x�������1�ƿ ؿ���� ϯ�D�V� h�zόϞ�-������� ��
�߫Ͻ�R�d�v� �ߚ߬�;�������� �*��N�`�r��� ��7�I�������&� 8�#�\�n��������� ��������"4F ��j|����S ��0BT� x�����a� //,/>/P/�t/�/ �/�/�/�/�/o/?? (?:?L?^?I��?�?�? �?�?�?�?�/O$O6O HOZOlO�?�O�O�O�O �O�OyO_ _2_D_V_ h_z_	_�_�_�_�_�_ �_�_o.o@oRodovo o�o�o�o�o�o�o �o*<N`r�o? ������ 8�J�\�n�����!��� ȏڏ��������F� X�j�|�����/�ğ֟ �������B�T�f� x�����+�=�ү��� ��,���P�b�t���������z�$UI_�PANEDATA 1N���ڱ�  	��}/frh/�cgtp/wid�edev.stm����%�7�I�Y�)Gpriρ�@�}����ϻ�������� ) �)��M�4�q߃�j� �ߎ����������%��7��[�7����     H�d�Ϙ��� ������E����:�L� ^�p������������ ����$H/l ~e������o� ݰܳ7�<N `r����-�� �//&/8/�\/n/ U/�/y/�/�/�/�/�/ ?�/4?F?-?j?Q?�? �?%�?�?�?OO 0O�?TO�xO�O�O�O �O�O�OKO_�O,__ P_b_I_�_m_�_�_�_ �_�_oo�_:o�?�? po�o�o�o�o�oo�o  sO$6HZl~ �o�������  �2��V�=�z���s� ����ԏGoYo�.� @�R�d�v�ɏ���� П������<�N� 5�r�Y�������̯�� �ׯ�&��J�1�n� ������ȿڿ��� �c�4ϧ�X�j�|ώ� �ϲ���+�������� 0�B�)�f�Mߊߜ߃� �ߧ��������� P�b�t�������� ��S���(�:�L�^� ���i�����������  ��6ZlS`�w�'�9�}��@�"4FX)� }��l����� /j'//K/2/D/�/ h/�/�/�/�/�/�/�/�#?5??Y?��C�=���$UI_POST�YPE  C��� 	 �e?�?�2QUICK�MEN  �;��?�?�0RESTO�RE 1OC��  ��L?��6OCC1O��m aO�O�O�O�O�OuO�O __,_>_�Ob_t_�_ �_�_UO�_�_�_M_o (o:oLo^oo�o�o�o �o�o�oo $6 H�_Ugy�o�� ���� �2�D�V� h��������ԏ ����w�)�R�d�v� ����=���П���� ��*�<�N�`�r��� �����ޯ���&� ɯJ�\�n�������G��ȿڿ�����7SC�RE�0?�=�u1sc+@uU2K�3K�4K�5Kĕ6K�7K�8K��2U�SER-�2�D�ksTMì�3��4��5�ĕ6��7��8���0N�DO_CFG �P�;� ��0PDA�TE ����None�2��_INFO 1QC�@��10%�[��� Iߊ�m߮��ߣ����� �����>�P�3�t���i���<-�OFFS_ET T�=�� ��$@������1�^� U�g������������ ����$-ZQcu���?�
�����UFRAME  �����*�RTO?L_ABRT	(��!ENB*GR�P 1UI�1Cz  A��~��@~���������0UJ�9MSK  M@�;-N%8�%��/��2VCCM��V��ͣ#RG�#Y�9����/����D�BeH�p71C����3711?�C0�$MRf2_�*S��괰	���~XC56 *�?�6�Y��1$�5����A@3C��. 	��8�?��OO KOx1FOsO�5�51ⴰ_O�O�� B����A2�DWO �O7O_�O8_#_\_G_ �_k_}_�__�_�_�_��_"o�OFoXo�%TCC�#`mI1�i���u��� GFS�»2aZ; �| 2�345678901�o�b�����o@��!5a�4BwB�`�56 311:�o=L�Br5v1�1~1�2 ��}/��o�a��# �GYk}�p�� �����ُ�1�C� U�6�H���5�~���ߏ����	���4�dSEGLEC)M!v1b3��VIRTSYN�C�� ���%�SIONTMOU�������F��#b�ֳ�ֵ(�u FR:\�H�\�A\�� ��� MC��L�OG��   U�D1��EX����'� B@ �����̡m��̡  �OBCL�1�H�� �  =	 �1- n6 � -������[�,xS�A�`=��͗���ˢ��TRA�IN⯞b�a1l�
�0d�$j�T2cZ; (aE2ϖ�i�� ;�)�_�M�g�qσϕ� ���������	��F�STAT dmB~2@�zߌ�*j$i�\���_GE�#eZ;7�`0�
� 0}2��HOMIN� �f־�ֿ� ~�����БC�g��X���JMPERR� 2gZ;
   ��*jl�V�7������ ��������
��2�@��q�d�v�B�_ߠREr� hWޠ$LEX�ԹiZ;�a1-e��V�MPHASE  �5��c&��!OF�F/�F�P2n�jJ�0�㜳E1�@��0ϒE1!1?s#33�����ak/�@kxk䜣!W�m[�䦲�[����o3;� [ i{���� /�O�?/M/_/q/ ��/��//�/'/9/ �/=?7?I?s?�/�?�/ �/�?�??Om?O%O 3OEO�?�?�O�?�O�O �?�O�O�O__gO\_ �OE_�O�_�O�O/_�_ �_�_oQ_Fou_�_|o �o�_�oo�o�o�o�o ;oMo?qof-�oI �����7� [P��������� ˏ��!�3�(�:�i��[�ŏg�}������TD_FILTEW��n�� �ֲ:���@���+�=�O�a� s���������֯� ����0�B�T�f�x����SHIFTME�NU 1o[�<��%��ֿ����ڿ� ���I� �2��V�h� ���Ϟϰ�������3��
�	LIVE/�SNAP'�vs�fliv��E�����ION * U<b�h�menu~߃������ߣ���p����	����E�.ォ50�s�P�@� �Z�AɠB8z�z�!�}��x�~�P��� ���MERb���<�0���kMO��q���z��WAITDINE�ND������O9K1�OUT���SD��TIM����o�G���#����C���b������RELEASE������TM�������_�ACT[�����_DATA r�%L����xRD�ISb�E�$X�VR�s���$Z�ABC_GRP �1t�Q�,#�r0�2���ZIP�u'�&����[�MPCF_G 1	v�Q�0�/� �w�ɤ� 	|�Z/  85�`�/�/H/�/l$?��+ �/�/�/?�/�/???|r?�?  �D0 �?�?�?�?�?�;����x�]hYLI�ND֑y� ���� ,(  * VOgM.�SO�OwO�O�M i?�O�O^PO1_ �OU_<_N_�_�O�_�_ �__�_�_x_-ooQo�8o�_�o�oY&#2z� ���oC� e?a?>N|�oq��햋qA�$DSPH�ERE 2{6M� �_�;o���!�io |W�i��_��,��Ï ���Ώ@��/�v��� e�؏��p�����������ZZ�� � N