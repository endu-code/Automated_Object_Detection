��   ��A��*SYST�EM*��V8.3�0261 5/�21/2018 A 	  ����DRYRUN�_T   � �$'ENB �4 NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��SAW_� G �%$INIT�	RESUME_/TYPEN &J�_  4 �$($FST_IcDX�P_ICI�0 �MIX_BG�-A
_NAM�c MODc_U�Sd�IFY_T�I� sxMK�R-  $�LINc   �_SIZcv� �k. , $?USE_FL4 ���&i*SIM�A�Q#QB6'S�CAN�AXS+I�NS*I��_COU�NrRO��_!_?TMR_VA�g�h>�i)  �'` ��R��!�+�WAR�$}H��!{#NPCH���$$CLASS  ���01���5��5%0VER�S�.7 � �@2IRTU�� .?@0'/ l5W5��������Y0�6m071�5��%@71�?���?
O��}5I2�;�GOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_���%FW?N8�0 ����_�_�_��s@�o { 2�;� 4%L_AOND_Bt_���Q?I��%L Jo���:dLmu�%[o�o7g�1zo�o 
�X�o�o�o�o���p
Oa @�dvu�S���=��9Y0ma`�s�1�t�al1Y0�>�&�8� J�\�n���������ȏ ڏ����6�1��1 � 2�D�V�h�z������� ԟ���
�44�6�S�!2�9 �[�m�������� ǯٯ����!�3� � M�f�x���������ҿ �����,�>�I�b� tφϘϪϼ������� ��(�:�L�W�p߂� �ߦ߸������� �� $�6�H�S�e�~��� ����������� �2� D�V�a�z��������� ������
.@R do������� �*<N`k }������/ /&/8/J/\/n/F