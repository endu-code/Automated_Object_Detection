��   $��A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN �/ MON_DAT�A6 p	$�ENABLF$�BASF   ��_NORMG ?$LIMIT��>�ERROR��ơIOCO/ CN�TR_CTM6� �$PF_�ENBG 	VL��PDD_POSRGN%��� LF� CTP�U-a>TDsIS� � FCG΍FRQ>/ EL�CPN F6 P�$�DTMA�NU �SE�RNO�OPFL��MODE�SFoTVER� q�C_GRP6�� 2$FS_FGORC� ��P�S_MEA2'%� 	1GF#2G0 �GTSK_CHKY%�O RIc"]!A�PP�$PS_oAAML��$�"v�	$/!_MI2�$AS�!!�#'#��#�!�3  2 �ROM_RU2�$J� EST2!y$� �N_NU��$u �  
$�SB*BSCNC�TOINS29FS� _NG$G�AGEx� � C�UTFREQY#L=R*REAL%� ��2MOMEN�TV�VC�F�C�f�2NC�K1DT�>�1DEVIDS�7� 	�3PATuH�0A�3FNA� 6!	AEX� �5O n�8BUF�7TDP8�Y�FLGEJ5���  � N I2U
@!(UF*����4OS0�	 DMM�A@ ? @ $�AbE?REG_OF�B�BME�HAS�C1�A� �DRE-  ? � �0�BB{F S{T� M�D|TRS$STD6XlQCWFA� 7X�QCW��"YV�"eS/ �A7 �  $�@TI�Nd@�0SULگ �R_@ g $}@ SW�@�RO�RR%	� �P�T� �@J�U� �SqFS4DN6
 �2P�0_@�cFOL[d!$�FIL� jjE�P��C�S�aDIG4R_C_SCA��c�INTTHRS�_BIdA�dSMA9L�bCOL�b9G�`� �� ��_IVTIM��$!0B"$S�?0xCCBDDN���-qI2wT2wDE�BUdA\!SCHN�"TOfa0�! �  Q0mr<0V� �;!�r~AUTTUN�� TRQa�uE�40N �qFS3A	XG  � 1eb}tj�rI�v	"G_gr>7 l �!�3>@WEIGH�q�2� uS_5QF(�T�2�WA� 	pEsNTERVA�; -  Q�� S!�t�AS0S��$J-_STAF�p JQg���1(�U��2��3��W����� hqx��"COG+_X�Y�Z�ҁCM�p?�p�܂RSLT�4��D��D��	"_�p_�q7  �~�b#0�VROUNDCMV�PERIODA�1�PUU3F2D�'TaM1� �Ƒ_D��GAMMc1��TRXI�K�K��K��CLbP�&On00ADJ�GAu��UPDB	"I%�0 ,$M"Pp30f��� d��:pG p"��HCDv�GV�#GVY��Z�JDO5�,q���S��$R��E_�8@{٣�pAP�HBC��$VF6�P��2L��蘨@IL[����;����;�d@���RG���NGEW_���r�Q}�8��ڡ�5OBOA@fQY�sW2/�G<�	����ȴ\�2�E�KP��NUCNPRGOVp����@`d_TW�cj,�G�E^!NV2#�C�c0@�WTS�T�RL_SKI2!�$SJ�Q��NQpG�W��u���7 \� ;0FR]b� � CMDC���T���b���TO?��� �5گ���_�Ah 0 |'��ALARM��_�*�TOT6�FRZn l�,!Y 3��X! ��mӥ�X �Œ`X ��(��U#��2��2
�X#�Z���FIX�8��Fȯ"��IT�`IB2�PN_d��CH�%�Υ�_DFL _�BF2N�ڶ�3������ ��3�"������P��� ����3��3
�8�X��DIA����/#� ���%�����[1��g1�[��� Z��#��!���%���$0�@
p��7F��YD�� HA�pU�5x����v�FSIW6� �2PN@�`R�>!�PHMP�`HCK%���>0G�'*#�e A����pNTడ^H	��HUFR zs3��A��UgvCa��$v0Q �����@p@p ̷  SI0�� P�5�IR�TU_��� %SV� 2���   A�6>0]@]�	Q�EF@ �oP�   �p � �//�'/9/K/U%@pd@p
m hK�/w/�/�/�( ��$��/� �/�/? .8e"�/?J?\?r?8? �?|?�?�?�?�?�?�? >O4ObOO�OTO�O�O jO|O�O�O�O_�O(_ _\_f_�_B_�_�_�_ �_ o�_$o�_Ho>oo ^b�/�ot��%�/�o�o��k	MC: �5678  A�fsdt1 78?901234q�#5w  	q �6xz.Ops�'��j l�o�o����������,�5�DMM 1�)5�A ���x�������=���ORw 2	Q� ���m��_� tu�B?)DN~�S4D 
Q�#!tY�d�!Ls|��q`rƈ̀?�l�B�𴐠�$ ONF�IG ��(� -� �����i!s�� 2��,
Hand� guide��?��3���  ��X��с��ь��g#�=���A ��ύ�������p� ݯ�(��L�7�p�[�<���m*���� ��ʿܿ� ��$�6� H�Z�lɌ��ό��ϰπ�������
�C�E�I� 2Q�(�0�� -�zՀ�Fտ&��_`πB���Ԟd�C�  ��uq=�#�
_aNnk(���K����̥@���e��=D�����_a;����8�I��_aIt$� �$F�>����k"���Q�Fۀ3]儢ѯǯ�����!�/�``+��̞��.�����_a$�敕��(4$�x����>�E���B<~w%�_a8E{�y5�;�jA���Ҝ�Q�>�	�]�_a?��m��箑�����~u1�?�33x����0�:�o�� ��0�����LSB��~uq�ӻ��m��S]���8��� ���t�	eF|���(]��߯����<n��;�.����=3�'	�����B���4* �2/V��%D�DH#  *%v�+��^-��
�/��/u/~u#�J/l/�)AI��/p�/�?/ A��n5��p��4vO?;)@�7�?�?�o�?�8Jhq�?�?zyjG�_FSIW Q��9�� O�O�Ou�