��   ʇ�A��*SYST�EM*��V8.3�0261 5/�21/2018 A   ����DCSS_C�PC_T� �$COMMENT� $ENA�BLE 6 MO�DJGRP_NU�MKL\  ?$UFRM\] ?_VTX 6 � �  $Y�Z�1K $Z2�STOP_TYPK�DSBIO�ID�XKENBL_C�ALMD�USE_PREDIC? � &S. �c 8J\TC�~u
SPD_LI_0���SOL�&|Y0  � 1CHG_SIZO$APGESDIS��G�!C����Jp 	�J�� &�"��))$'2_SE��� XPANIN�  �STAT�/ D $F�P_BASE �$_ K�$!� �&_V�.H�#:g%J- ��ZAXS\UPR�JLW7Se���&� | 
 �/�/�/D&?8?zh$�ELEM/ Tc ��2�"NOG<�0�3UTOOi�2�HAD�� $D7ATA"g%e�0  @@p:�0 _2 
&Pp%' � p!U*n   �FS�Cz�B�� �B(�F�D(�R|UC�DROBOT�H��CqBo�E�F$�CUR_2Rh$SwETU�	 l� ��P_MGN�I?NP_ASS�0 "@�� �3�8B7gP@U��^V�Sp!�h$T1�
`B|8�8�TM 0 �6P�+ Ke�1VRCFY�8
dD5F1� ��W��1$R��8SPH/ (�{ �CA�CA�CA3�BOX/ 8 �0������b'o�EjTUIR�0 � ,{ FR`ER��02 $�` ��a_S�b��gZN/ 0 �{9F0� -a0rZ	_0�_0�u0  @Q�Yv	�o:o� �$$CLLP ? ����q���Q��Q�pVERSwION�xZ0��5�qIRTU�AL��q' 2 ��xQ   ��Double �Parts Si�de�� �0�p����#PD  �DM-�N�� � �@k����� ����M@2���q��/�A�S�f D���
�y�DJ@ QD�p+������� ����r��a�W�u�� ��ٟ�Z��~���Ɵ ��F�{������� �2� h�����/���S�¯ ԯ毛�
���ѿ@��� d�v���=Ϭ�a�s�� �ς��*���N��� ��%�Kߺ��ρ��ϥ� ��N�8���\�n�#�� G�Y�k��ߏ������ 4������|�1���� 9���w��������B� T���x�
?Q��u ����,����b ���_��� �(:L/p%/ 7/�[/F/���// �/�/H/�/?~/�/E? �/i?{??�/�? ?2? �?V?OO/O�?SO�? �?�O�?�O�O�O@O�O dOvO�O�O;_a_s_�O �___N_<_�_oo �_9o�_�_�_�opo�o �o&o�oJo\ono#�o GY�o}�o�o� 4��j�
��� g���������ӏB� T�	�x�-�?�֏��u� ������ϟ��b� �����M���q����� ���(�:���^���%� 7���[�ʯܯ� ��� ǿٿH���l�~���E��4�i�{���$DC�SS_CSC 2�!���Q  D����� ��*ƶ������A�� S�4߉�X߭�|��ߠ� ���������<�a�0� B��f������� ��'���K��o�>�P� ��t����������� 5Y(}L^����'ɘ�GRP ;2�� ��,�	Z�?*cN�r ������/)/ /M/8/q/\/�/�/�/ �/�/�/?�/�/7?"? [?F??j?�?�?�?�? �?�?�?!OOEO0OiO TO�O�O�O|O�O�O�O �O�O/__S_>_w_�_ �_f_�_�_�_�_�_o o=o(oaoso�oPo�o �o�o�o�o�o�o' K]o:�~��������5��_�GSTAT 2���1�,8���}OH�Ơ-��ۣ�����?{#�>!6��=�2�>+�&��{O�B7�b�ı��B����$�8t�<�m���`/�4�z�2
�A?� � �����4��Z�@v����T�/������痿-���?;�l���v�?;ڌ?-�ـ̉A���+��D�Z���J��%��?�C?��<�n�{�탳��T��?B��?%���A�	��C��iD-��䅽��Y�%y?A��<�@��~���=9�ս����B�sĳ��HC	/j䅼�� �|�/�[?u��9���=���2���+�;?{O� ��v�����ȑ���� �� �F�X�6�|����� ȁ'ɰ�%�����ԯ � �
��>�@�R�t� ������Կ⇔��`� ��D�V�4�zόϦ�� �ϼ���������"�� .�X�B�dߎ�xߊ��� ��l�����<�N�,��r��b�ȁ�C�C���y]�C�ｿɀ6_Ɔ��p�_}d��D|����2DQ���͸�R�-�IB�ԁ���ԁC?  ��!'���7��'4��Ȃɀ8�T�!���t��D�E��8i��4w�q1ȁ8�ǂﴨ��$��F�P��C����}�Dk�P��6��AN �Wp�����R��ঽOt�Dj����~���b(�"ȁ�u�u�8�yr6u[M ȁ�������h�:L *p�`������ ����$N8 J�n����� /�2/D/�h/z/X/ �/�/�/�//�/? �/?.?0?B?d?�?x? �?�?�?�?�? /*O<O �/`OrOPO�O�O�O�� 
���������"�4� F�X�j�|��������� ���_�O�O�Ojo�O Zo�o�o�o�o�o�/O �?H2T~h ������� � 
��ob�t�R������� Ώ���o4�
���@� *�L�v�`�r������� ʟ̟ޟ �*���Z�l� ��������Ưد�O(o :o�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo��No�Ϛϴ� ���Ϯ�������8� B��N�x�b߄߮ߘ� ����������&�P� :�ߒ��ς������ ���*�d�:�@�F�p� Z�|������������� ��H2��� z�����X� j�(�:�L�^�p����� ����ʿܿ� ��$� 6� 2D~ϸ/�/� �/ ?�/$?6?�F`? j\?~?�?�?�?�?�? �?O�? OJO4OVO�O r�O�O?�O�O�O_ ._H?Z?�Oj_pOv_�_ �_�_�_�_�_o�_o Bo,oNoxobo@_�o_ �o�o�o&8v/�/ �/Xj|���� ���//h/B/T/ f/Pbt���؏ �0��T�f�L_�o�� �o��Ɵ������� ��.�P�z�d����� �o��D��(��L� ^�x�����Ư������ ��ܿ���<�&�H� r�\�~Ϩ�ί����<� �� ���0�V�4ߦ��� ʏ������� ��*�<�N���r��� ��ߒ�̏F��*�� N�`�>�����|����� ��������,8 bL^����� v�" FX6| ��������� �$// /B/D/V/x/ �/�/�/�/�??l >?P?.?t?�?p����� �߸������� ��$� 6�H�Z�l�~���� �O�?�?��?H_�?X_ ~_\_n_�_�_��/�_ �/�_&oo2o\oFoho �o|o�o�o�o�o�o�o �_@R0v�f� ��_��o��� *�T�>�`���t����� ����ޏ���8�J�(��n���^������u�$�DCSS_JPC� 2�uQ ( D���#�� �%��G� �(�}�L�^�p�ů�� ӯ���ܯ1� �U�$� 6�x���l�~�ӿ���� ƿ��?��c�2χ� Vϫ�zό��ϰ����� )���7��q�@ߕ�d� �߈ߚ��������7� ��*��N��r��� ����������E�� &�8���\��������� ��������@e4 F�j|��� �+�OsBT �x������ 9//]/,/�/P/b/�/ �/�/�/�/�/�/�/G? ?k?:?�?^?�?�?�? �?�?O�?�? OUO$O�cO"�ԕSݐ�@ NO�OrODO�O�O_�O ?__$_u_H_Z_l_�_ �_�_�_�_�_�_;oo  o^o�oVoho�o�o�o �o�o�o7
E. Rd����� ��3���*�{�N� `���Ï������̏� ��A��&�w�J���n� ��������ȟڟ�=� �"�s�F�X�j����� ��ޯ�֯�9��]� 0���T�f�����ſ�� ��ҿ�5���,�}� P�bϳφϘϪ����� ���C��(�y�Lߝ� p��ߔߦ�������߀?��$�u�H�Z�HMODEL 2�K�xp�e�
 <���c��  g���l����� R�)�;�M�_�q����� ��������% 7�[m���� ���a�J��! �	w����/ ��B//+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?t?K?]?�?E W�?�?O?�?�?LO #O5O�OYOkO�O�O�O �O _�O�O6___l_ C_U_g_�_�_�_�_�_ �_ o�?�?�?oo�_ couo�o�o�o�o�o�o �o)vM_� ������*�� �`�7�I�[�1o��Uo ����k�ُ�8��!� n�E�W�i�{������ ß՟"�����/�A� S���w���֯����ѯ ��0�ˏ���x�O�a� ������俻�Ϳ߿,� ��b�9�KϘ�oρ� ���Ϸ��������L� #�5�G����A�o߁� ������$�����1� C�U��y������� ������	�V�-�?��� c�u����������� ������d;M�q ������ N%7I[m� ��/���/!/ 3/	�/-[/m/�/�/ �/?�/�/?X?/?A? �?e?w?�?�?�?�?O �?�?BOO+OxOOOaO sO�O�O�O/�/�/�O �OP_�O9_K_]_o_�_ �_�_�_o�_�_�_o #o5o�oYoko�o�o�o �o�o�o�o6l __GY�A�� ���D��-�z�Q� c�u���������Ϗ� .���)�;�M�_��� �����}���ϟ<� ��%�7���[�m����� ���ǯٯ�8��!� n�E�W���{������ ÿտ"����X��� �E�W�-ϛϭ����� ��0���+�=�O�a� �߅ߗ��߻������� ��b�9�K��o�� ��i���ϻ����� #�p�G�Y���}����� ������$��Z1 CUgy���� ��	��h�1 C������/ �//d/;/M/�/q/ �/�/�/�/�/?�/? N?%?7?�?[?m??U �?y�?�?&O�?O\O 3OEOWOiO{O�O�O�O �O_�O�O__/_A_ �_e_w_�_�_�_�_�_��_�_�:�$DCS�S_PSTAT ����_a�Q    �po~j no (��o�o�o�o�o | �```q�`7o0B�9*c_elpa�~�PdSETUP �	_iB�"d�3��1�tKiT1SC �2
�zp�1Cz��3��+��uCP [R�|��0D�? v����?����Џ��� ���<�N�`�/��� ��e���̟ޟ���� &���J�\�n�=����� ����گ��>d�!�3� ��W�i�{�J�����ÿ ������ڿ/�A�� "�wω�XϭϿ��Ϡ� ������=�O�a�0� �ߗ��������f�� �'���K�]�o�>�� �����������#� 5��Y�k�}�L����� ����������1C �߼�y���� ��	�?Qc 2��hz��� //)/�M/_/q/@/ �/�/�/�/�/�/Vh %?7?�/[?m??N?�? �?�?�?�?�?O�?3O EOO&O{O�O\O�O�O �O�O�O__�OA_S_ e_4_�_�_??�_�_ j_oo+o�_Ooaoso Bo�o�o�o�o�o�o�o �o'9]o�P �������� 5�G��_�_}������ ŏ׏�������C� U�g�6�����l�~�ӟ 埴�	��-���Q�c� u�D����������� Z�l�)�;�¯_�q��� R�����˿����� �7�I��*�ϑ�`� �����Ϩ����!��πE�W�i�8ߍߟ߯���$DCSS_TC�PMAP  ������Q_ @ z�zХz�z���z��z�z�z�	� � z�z�z��z�z�z�z��z�z�z�z�Jz�z�z�z�z�Uz�z�z�z�Uz� z�!z�"z�U#z�$z�%z�&z�U'z�(z�)z�*z�U+z�,z�-z�.z�U/z�0z�1z�2z�U3z�4z�5z�6z�U7z�8z�9z�:z�U;z�<z�=z�>z��?z�@��UIROw 2����� ���0�B�T�f� x���������������@,>Py�� y������� 	-?Qcu� ����Z�~� )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?�?
/�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O�r?_��UIZN �2��	 ��� ��L_^_p_u�G_�_�_ �_�_�_�_o�_,o>o Pooto�o�ogo�o�o �o�o�o(�oL^ p�E�����  ���6�H�Z�)�~� ����e�Ə؏ꏹ��  �2���V�h�z�I��� ��ԟ����
�ٟ.��@�R�_��UFRM� R����8 }ߪ���{���ͯ� (��L�^�9�����o� ��ʿ��� �ۿ$�6� �G�l�~ϕ��ϴ�S� ������� ���D�V� 1�zߌ�g߰��ߝ��� ��
���.�@��d�v� �Ϛ��K������� ���<�N�)�_����� q�����������& 8\n���C ����"�F X3|�i��� ���/0//T/f/ }t/�/�/�/�/�/�/ ??�/>?P?+?t?�? a?�?�?�?�?�?�?O (OOLO^Ou/�/�O�O EO�O�O�O __�O6_ H_#_l_~_Y_�_�_�_ �_�_�_�_ o2ooVo hoO�o�o=o�o�o�o �o
�o.@dv Q������� �*��N�`�wo���� 5���̏�����ݏ� 8�J�%�n���[����� ��ڟ�ǟ�"���F� X�2�